magic
tech sky130A
magscale 1 2
timestamp 1654519532
<< viali >>
rect 3065 47141 3099 47175
rect 29929 47141 29963 47175
rect 31033 47141 31067 47175
rect 47961 47141 47995 47175
rect 2053 47073 2087 47107
rect 12357 47073 12391 47107
rect 12633 47073 12667 47107
rect 16957 47073 16991 47107
rect 43177 47073 43211 47107
rect 47041 47073 47075 47107
rect 1777 47005 1811 47039
rect 3801 47005 3835 47039
rect 4813 47005 4847 47039
rect 6377 47005 6411 47039
rect 7297 47005 7331 47039
rect 9413 47005 9447 47039
rect 14105 47005 14139 47039
rect 14933 47005 14967 47039
rect 16681 47005 16715 47039
rect 19257 47005 19291 47039
rect 20913 47005 20947 47039
rect 22017 47005 22051 47039
rect 24869 47005 24903 47039
rect 28549 47005 28583 47039
rect 29745 47005 29779 47039
rect 31217 47005 31251 47039
rect 38393 47005 38427 47039
rect 40509 47005 40543 47039
rect 41889 47005 41923 47039
rect 42625 47005 42659 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 2789 46937 2823 46971
rect 4077 46937 4111 46971
rect 6653 46937 6687 46971
rect 9597 46937 9631 46971
rect 15117 46937 15151 46971
rect 19533 46937 19567 46971
rect 28733 46937 28767 46971
rect 40325 46937 40359 46971
rect 42809 46937 42843 46971
rect 45385 46937 45419 46971
rect 4905 46869 4939 46903
rect 7481 46869 7515 46903
rect 14289 46869 14323 46903
rect 21833 46869 21867 46903
rect 5825 46597 5859 46631
rect 13369 46597 13403 46631
rect 1409 46529 1443 46563
rect 24593 46529 24627 46563
rect 38117 46529 38151 46563
rect 47961 46529 47995 46563
rect 3985 46461 4019 46495
rect 4169 46461 4203 46495
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 13829 46461 13863 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 31585 46461 31619 46495
rect 32137 46461 32171 46495
rect 32321 46461 32355 46495
rect 32597 46461 32631 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 22017 46393 22051 46427
rect 1593 46325 1627 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 4629 46121 4663 46155
rect 5365 46121 5399 46155
rect 13093 46121 13127 46155
rect 14197 46121 14231 46155
rect 20177 46121 20211 46155
rect 24777 46121 24811 46155
rect 31861 46121 31895 46155
rect 38301 46121 38335 46155
rect 11713 45985 11747 46019
rect 20729 45985 20763 46019
rect 21281 45985 21315 46019
rect 25329 45985 25363 46019
rect 26709 45985 26743 46019
rect 41337 45985 41371 46019
rect 41889 45985 41923 46019
rect 46305 45985 46339 46019
rect 47041 45985 47075 46019
rect 2053 45917 2087 45951
rect 5273 45917 5307 45951
rect 11989 45917 12023 45951
rect 13001 45917 13035 45951
rect 14105 45917 14139 45951
rect 20085 45917 20119 45951
rect 24685 45917 24719 45951
rect 31769 45917 31803 45951
rect 38209 45917 38243 45951
rect 43913 45917 43947 45951
rect 45661 45917 45695 45951
rect 20913 45849 20947 45883
rect 25513 45849 25547 45883
rect 41521 45849 41555 45883
rect 45845 45849 45879 45883
rect 46489 45849 46523 45883
rect 44097 45781 44131 45815
rect 20821 45577 20855 45611
rect 25513 45577 25547 45611
rect 41429 45577 41463 45611
rect 42533 45577 42567 45611
rect 43177 45509 43211 45543
rect 43821 45509 43855 45543
rect 47685 45509 47719 45543
rect 1777 45441 1811 45475
rect 13921 45441 13955 45475
rect 20729 45441 20763 45475
rect 25421 45441 25455 45475
rect 41337 45441 41371 45475
rect 42441 45441 42475 45475
rect 43085 45441 43119 45475
rect 46765 45441 46799 45475
rect 47593 45441 47627 45475
rect 1961 45373 1995 45407
rect 2789 45373 2823 45407
rect 26249 45373 26283 45407
rect 44465 45373 44499 45407
rect 44649 45373 44683 45407
rect 45845 45373 45879 45407
rect 43913 45237 43947 45271
rect 46949 45237 46983 45271
rect 2237 45033 2271 45067
rect 43821 45033 43855 45067
rect 45109 45033 45143 45067
rect 45753 45033 45787 45067
rect 44465 44897 44499 44931
rect 48145 44897 48179 44931
rect 2145 44829 2179 44863
rect 45017 44829 45051 44863
rect 45661 44829 45695 44863
rect 46305 44829 46339 44863
rect 46489 44761 46523 44795
rect 46305 44489 46339 44523
rect 47685 44489 47719 44523
rect 45753 44353 45787 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 38577 44285 38611 44319
rect 38761 44285 38795 44319
rect 40049 44285 40083 44319
rect 45109 44149 45143 44183
rect 46949 44149 46983 44183
rect 28181 43945 28215 43979
rect 38761 43945 38795 43979
rect 45845 43945 45879 43979
rect 46305 43809 46339 43843
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 28089 43741 28123 43775
rect 38669 43741 38703 43775
rect 1409 43265 1443 43299
rect 46857 43265 46891 43299
rect 1685 43197 1719 43231
rect 47777 43061 47811 43095
rect 46305 42721 46339 42755
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 48145 41497 48179 41531
rect 2145 41225 2179 41259
rect 46949 41225 46983 41259
rect 2053 41089 2087 41123
rect 46857 41089 46891 41123
rect 47961 41089 47995 41123
rect 48145 40953 48179 40987
rect 47685 40681 47719 40715
rect 1869 40409 1903 40443
rect 1961 40341 1995 40375
rect 47777 39797 47811 39831
rect 24961 39457 24995 39491
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 23397 39389 23431 39423
rect 24777 39389 24811 39423
rect 46489 39321 46523 39355
rect 23213 39253 23247 39287
rect 24409 39253 24443 39287
rect 24869 39253 24903 39287
rect 46857 39049 46891 39083
rect 20269 38981 20303 39015
rect 22753 38981 22787 39015
rect 20453 38913 20487 38947
rect 44281 38913 44315 38947
rect 46765 38913 46799 38947
rect 47869 38913 47903 38947
rect 22477 38845 22511 38879
rect 45017 38845 45051 38879
rect 48053 38777 48087 38811
rect 20637 38709 20671 38743
rect 24225 38709 24259 38743
rect 22753 38505 22787 38539
rect 20545 38437 20579 38471
rect 23857 38437 23891 38471
rect 23397 38369 23431 38403
rect 42993 38369 43027 38403
rect 44373 38369 44407 38403
rect 45477 38369 45511 38403
rect 17141 38301 17175 38335
rect 17325 38301 17359 38335
rect 20361 38301 20395 38335
rect 22661 38301 22695 38335
rect 23489 38301 23523 38335
rect 42625 38301 42659 38335
rect 43821 38301 43855 38335
rect 45109 38301 45143 38335
rect 46305 38301 46339 38335
rect 46489 38233 46523 38267
rect 48145 38233 48179 38267
rect 17233 38165 17267 38199
rect 26433 37961 26467 37995
rect 46857 37961 46891 37995
rect 21925 37893 21959 37927
rect 23305 37893 23339 37927
rect 21833 37825 21867 37859
rect 23581 37825 23615 37859
rect 27813 37825 27847 37859
rect 44281 37825 44315 37859
rect 46765 37825 46799 37859
rect 47777 37825 47811 37859
rect 19533 37757 19567 37791
rect 19809 37757 19843 37791
rect 23489 37757 23523 37791
rect 24685 37757 24719 37791
rect 24961 37757 24995 37791
rect 45109 37757 45143 37791
rect 21281 37689 21315 37723
rect 23305 37621 23339 37655
rect 23765 37621 23799 37655
rect 27905 37621 27939 37655
rect 20453 37417 20487 37451
rect 21097 37417 21131 37451
rect 25145 37417 25179 37451
rect 44281 37417 44315 37451
rect 20269 37281 20303 37315
rect 2053 37213 2087 37247
rect 20085 37213 20119 37247
rect 20453 37213 20487 37247
rect 20913 37213 20947 37247
rect 21925 37213 21959 37247
rect 24409 37213 24443 37247
rect 25329 37213 25363 37247
rect 25881 37213 25915 37247
rect 25973 37213 26007 37247
rect 26709 37213 26743 37247
rect 44189 37213 44223 37247
rect 22201 37145 22235 37179
rect 24501 37145 24535 37179
rect 26985 37145 27019 37179
rect 20177 37077 20211 37111
rect 23673 37077 23707 37111
rect 28457 37077 28491 37111
rect 22109 36873 22143 36907
rect 23489 36873 23523 36907
rect 25789 36873 25823 36907
rect 26985 36873 27019 36907
rect 28365 36805 28399 36839
rect 1777 36737 1811 36771
rect 15761 36737 15795 36771
rect 17325 36737 17359 36771
rect 21833 36737 21867 36771
rect 23305 36737 23339 36771
rect 23673 36737 23707 36771
rect 23857 36737 23891 36771
rect 25605 36737 25639 36771
rect 27169 36737 27203 36771
rect 27261 36737 27295 36771
rect 27537 36737 27571 36771
rect 28181 36737 28215 36771
rect 29009 36737 29043 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 17601 36669 17635 36703
rect 22109 36669 22143 36703
rect 27445 36669 27479 36703
rect 27997 36669 28031 36703
rect 21925 36601 21959 36635
rect 15853 36533 15887 36567
rect 19073 36533 19107 36567
rect 23765 36533 23799 36567
rect 29101 36533 29135 36567
rect 2237 36329 2271 36363
rect 18245 36261 18279 36295
rect 22661 36261 22695 36295
rect 24961 36261 24995 36295
rect 25145 36261 25179 36295
rect 14749 36193 14783 36227
rect 19533 36193 19567 36227
rect 2145 36125 2179 36159
rect 18429 36125 18463 36159
rect 18613 36125 18647 36159
rect 18705 36125 18739 36159
rect 19441 36125 19475 36159
rect 22845 36125 22879 36159
rect 23121 36125 23155 36159
rect 23581 36125 23615 36159
rect 27629 36125 27663 36159
rect 15025 36057 15059 36091
rect 24685 36057 24719 36091
rect 27445 36057 27479 36091
rect 16497 35989 16531 36023
rect 19809 35989 19843 36023
rect 23029 35989 23063 36023
rect 23673 35989 23707 36023
rect 27813 35989 27847 36023
rect 18337 35785 18371 35819
rect 19533 35785 19567 35819
rect 23213 35785 23247 35819
rect 23673 35785 23707 35819
rect 24317 35785 24351 35819
rect 24977 35785 25011 35819
rect 25145 35785 25179 35819
rect 27261 35785 27295 35819
rect 27445 35785 27479 35819
rect 19253 35717 19287 35751
rect 22753 35717 22787 35751
rect 24777 35717 24811 35751
rect 1593 35649 1627 35683
rect 15577 35649 15611 35683
rect 16865 35649 16899 35683
rect 16957 35649 16991 35683
rect 17233 35649 17267 35683
rect 18245 35649 18279 35683
rect 18981 35649 19015 35683
rect 19165 35649 19199 35683
rect 19349 35649 19383 35683
rect 23029 35649 23063 35683
rect 26249 35649 26283 35683
rect 26433 35649 26467 35683
rect 27386 35649 27420 35683
rect 27905 35649 27939 35683
rect 28641 35649 28675 35683
rect 48145 35649 48179 35683
rect 15669 35581 15703 35615
rect 17141 35581 17175 35615
rect 22937 35581 22971 35615
rect 24041 35581 24075 35615
rect 24133 35581 24167 35615
rect 28917 35581 28951 35615
rect 1409 35445 1443 35479
rect 15853 35445 15887 35479
rect 16681 35445 16715 35479
rect 23029 35445 23063 35479
rect 24961 35445 24995 35479
rect 26249 35445 26283 35479
rect 27813 35445 27847 35479
rect 30389 35445 30423 35479
rect 47961 35445 47995 35479
rect 15577 35241 15611 35275
rect 15945 35241 15979 35275
rect 20729 35241 20763 35275
rect 22845 35241 22879 35275
rect 24593 35241 24627 35275
rect 25237 35241 25271 35275
rect 27261 35241 27295 35275
rect 24501 35173 24535 35207
rect 27445 35173 27479 35207
rect 24685 35105 24719 35139
rect 25697 35105 25731 35139
rect 15761 35037 15795 35071
rect 16037 35037 16071 35071
rect 18337 35037 18371 35071
rect 20545 35037 20579 35071
rect 21741 35037 21775 35071
rect 21925 35037 21959 35071
rect 22017 35037 22051 35071
rect 23029 35037 23063 35071
rect 23213 35037 23247 35071
rect 23489 35037 23523 35071
rect 24410 35047 24444 35081
rect 25421 35037 25455 35071
rect 25513 35037 25547 35071
rect 25789 35037 25823 35071
rect 26341 35037 26375 35071
rect 27169 35037 27203 35071
rect 27261 35037 27295 35071
rect 28089 35037 28123 35071
rect 28181 35037 28215 35071
rect 28365 35037 28399 35071
rect 28457 35037 28491 35071
rect 30021 35037 30055 35071
rect 30389 35037 30423 35071
rect 48145 35037 48179 35071
rect 23121 34969 23155 35003
rect 23331 34969 23365 35003
rect 26985 34969 27019 35003
rect 30205 34969 30239 35003
rect 30297 34969 30331 35003
rect 18429 34901 18463 34935
rect 21557 34901 21591 34935
rect 26433 34901 26467 34935
rect 27905 34901 27939 34935
rect 30573 34901 30607 34935
rect 47961 34901 47995 34935
rect 23489 34697 23523 34731
rect 27353 34697 27387 34731
rect 29377 34697 29411 34731
rect 21833 34629 21867 34663
rect 23121 34629 23155 34663
rect 24041 34629 24075 34663
rect 25237 34629 25271 34663
rect 30941 34629 30975 34663
rect 15301 34561 15335 34595
rect 17417 34561 17451 34595
rect 20361 34561 20395 34595
rect 20545 34561 20579 34595
rect 20913 34561 20947 34595
rect 22109 34561 22143 34595
rect 23305 34561 23339 34595
rect 26157 34561 26191 34595
rect 26985 34561 27019 34595
rect 27169 34561 27203 34595
rect 28641 34561 28675 34595
rect 28825 34561 28859 34595
rect 28917 34561 28951 34595
rect 29193 34561 29227 34595
rect 30757 34561 30791 34595
rect 31033 34561 31067 34595
rect 47777 34561 47811 34595
rect 17693 34493 17727 34527
rect 20637 34493 20671 34527
rect 20729 34493 20763 34527
rect 22017 34493 22051 34527
rect 25421 34493 25455 34527
rect 26433 34493 26467 34527
rect 29009 34493 29043 34527
rect 24225 34425 24259 34459
rect 15393 34357 15427 34391
rect 19165 34357 19199 34391
rect 21097 34357 21131 34391
rect 21833 34357 21867 34391
rect 22293 34357 22327 34391
rect 26249 34357 26283 34391
rect 26341 34357 26375 34391
rect 27077 34357 27111 34391
rect 30573 34357 30607 34391
rect 47593 34357 47627 34391
rect 18521 34153 18555 34187
rect 21741 34153 21775 34187
rect 22293 34153 22327 34187
rect 23581 34153 23615 34187
rect 24593 34153 24627 34187
rect 31106 34153 31140 34187
rect 22753 34085 22787 34119
rect 14197 34017 14231 34051
rect 16865 34017 16899 34051
rect 18153 34017 18187 34051
rect 19993 34017 20027 34051
rect 20269 34017 20303 34051
rect 26433 34017 26467 34051
rect 29929 34017 29963 34051
rect 30849 34017 30883 34051
rect 47133 34017 47167 34051
rect 47409 34017 47443 34051
rect 1593 33949 1627 33983
rect 16589 33949 16623 33983
rect 16681 33949 16715 33983
rect 16957 33949 16991 33983
rect 17785 33949 17819 33983
rect 17969 33949 18003 33983
rect 18061 33949 18095 33983
rect 18337 33949 18371 33983
rect 22201 33949 22235 33983
rect 22477 33949 22511 33983
rect 24409 33949 24443 33983
rect 26157 33949 26191 33983
rect 26249 33949 26283 33983
rect 26525 33949 26559 33983
rect 26985 33949 27019 33983
rect 27169 33949 27203 33983
rect 30021 33949 30055 33983
rect 14473 33881 14507 33915
rect 23213 33881 23247 33915
rect 23397 33881 23431 33915
rect 47225 33881 47259 33915
rect 1409 33813 1443 33847
rect 15945 33813 15979 33847
rect 16405 33813 16439 33847
rect 25973 33813 26007 33847
rect 27077 33813 27111 33847
rect 30389 33813 30423 33847
rect 32597 33813 32631 33847
rect 15117 33609 15151 33643
rect 18429 33609 18463 33643
rect 20729 33609 20763 33643
rect 27445 33609 27479 33643
rect 30021 33609 30055 33643
rect 32873 33609 32907 33643
rect 48053 33609 48087 33643
rect 29377 33541 29411 33575
rect 14473 33473 14507 33507
rect 14657 33473 14691 33507
rect 15301 33473 15335 33507
rect 17877 33473 17911 33507
rect 18245 33473 18279 33507
rect 18889 33473 18923 33507
rect 19073 33473 19107 33507
rect 19349 33473 19383 33507
rect 20637 33473 20671 33507
rect 21833 33473 21867 33507
rect 22109 33473 22143 33507
rect 24225 33473 24259 33507
rect 25973 33473 26007 33507
rect 26157 33473 26191 33507
rect 27353 33473 27387 33507
rect 27997 33473 28031 33507
rect 29716 33473 29750 33507
rect 32137 33473 32171 33507
rect 32781 33473 32815 33507
rect 46857 33473 46891 33507
rect 47593 33473 47627 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 15577 33405 15611 33439
rect 26249 33405 26283 33439
rect 14565 33337 14599 33371
rect 15485 33337 15519 33371
rect 24409 33337 24443 33371
rect 28181 33337 28215 33371
rect 18245 33269 18279 33303
rect 19257 33269 19291 33303
rect 25789 33269 25823 33303
rect 29542 33269 29576 33303
rect 29653 33269 29687 33303
rect 32229 33269 32263 33303
rect 46949 33269 46983 33303
rect 47869 33269 47903 33303
rect 1961 33065 1995 33099
rect 14841 33065 14875 33099
rect 15393 33065 15427 33099
rect 17141 33065 17175 33099
rect 18061 33065 18095 33099
rect 21097 33065 21131 33099
rect 21925 33065 21959 33099
rect 15761 32997 15795 33031
rect 19625 32997 19659 33031
rect 24869 32997 24903 33031
rect 27169 32997 27203 33031
rect 30021 32997 30055 33031
rect 31217 32997 31251 33031
rect 32413 32997 32447 33031
rect 2329 32929 2363 32963
rect 14933 32929 14967 32963
rect 15485 32929 15519 32963
rect 17233 32929 17267 32963
rect 18245 32929 18279 32963
rect 25421 32929 25455 32963
rect 30389 32929 30423 32963
rect 1869 32861 1903 32895
rect 2973 32861 3007 32895
rect 14657 32861 14691 32895
rect 14749 32861 14783 32895
rect 15393 32861 15427 32895
rect 17141 32861 17175 32895
rect 17417 32861 17451 32895
rect 18337 32861 18371 32895
rect 19257 32861 19291 32895
rect 21005 32861 21039 32895
rect 23121 32861 23155 32895
rect 24777 32861 24811 32895
rect 28181 32861 28215 32895
rect 29929 32861 29963 32895
rect 30205 32861 30239 32895
rect 31125 32861 31159 32895
rect 31401 32861 31435 32895
rect 31493 32861 31527 32895
rect 32045 32861 32079 32895
rect 45845 32861 45879 32895
rect 46305 32861 46339 32895
rect 16221 32793 16255 32827
rect 16405 32793 16439 32827
rect 18061 32793 18095 32827
rect 19441 32793 19475 32827
rect 21833 32793 21867 32827
rect 25697 32793 25731 32827
rect 32229 32793 32263 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 2789 32725 2823 32759
rect 16589 32725 16623 32759
rect 17601 32725 17635 32759
rect 18521 32725 18555 32759
rect 22937 32725 22971 32759
rect 28273 32725 28307 32759
rect 31585 32725 31619 32759
rect 23857 32521 23891 32555
rect 25605 32521 25639 32555
rect 28365 32521 28399 32555
rect 29653 32521 29687 32555
rect 46949 32521 46983 32555
rect 48053 32521 48087 32555
rect 2421 32453 2455 32487
rect 15669 32453 15703 32487
rect 22385 32453 22419 32487
rect 28273 32453 28307 32487
rect 2237 32385 2271 32419
rect 15853 32385 15887 32419
rect 15945 32385 15979 32419
rect 17233 32385 17267 32419
rect 20821 32385 20855 32419
rect 22109 32385 22143 32419
rect 24317 32385 24351 32419
rect 27353 32385 27387 32419
rect 27445 32385 27479 32419
rect 27721 32385 27755 32419
rect 29285 32385 29319 32419
rect 29469 32385 29503 32419
rect 30389 32385 30423 32419
rect 32137 32385 32171 32419
rect 46857 32385 46891 32419
rect 47961 32385 47995 32419
rect 4077 32317 4111 32351
rect 17509 32317 17543 32351
rect 30113 32317 30147 32351
rect 32413 32317 32447 32351
rect 33885 32317 33919 32351
rect 16129 32249 16163 32283
rect 1777 32181 1811 32215
rect 15669 32181 15703 32215
rect 17509 32181 17543 32215
rect 17785 32181 17819 32215
rect 21005 32181 21039 32215
rect 27169 32181 27203 32215
rect 27629 32181 27663 32215
rect 16221 31977 16255 32011
rect 16589 31977 16623 32011
rect 22661 31977 22695 32011
rect 24409 31977 24443 32011
rect 25605 31977 25639 32011
rect 29929 31977 29963 32011
rect 30757 31977 30791 32011
rect 32505 31977 32539 32011
rect 33057 31977 33091 32011
rect 28733 31909 28767 31943
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 3985 31841 4019 31875
rect 4629 31841 4663 31875
rect 16681 31841 16715 31875
rect 17877 31841 17911 31875
rect 20085 31841 20119 31875
rect 20361 31841 20395 31875
rect 23489 31841 23523 31875
rect 23765 31841 23799 31875
rect 24869 31841 24903 31875
rect 25053 31841 25087 31875
rect 26985 31841 27019 31875
rect 27261 31841 27295 31875
rect 32045 31841 32079 31875
rect 46581 31841 46615 31875
rect 47409 31841 47443 31875
rect 3801 31773 3835 31807
rect 16405 31773 16439 31807
rect 17601 31773 17635 31807
rect 17785 31773 17819 31807
rect 17969 31773 18003 31807
rect 18153 31773 18187 31807
rect 22569 31773 22603 31807
rect 23397 31773 23431 31807
rect 24777 31773 24811 31807
rect 25513 31773 25547 31807
rect 25789 31773 25823 31807
rect 26065 31773 26099 31807
rect 29929 31773 29963 31807
rect 30113 31773 30147 31807
rect 30757 31773 30791 31807
rect 30941 31773 30975 31807
rect 31769 31773 31803 31807
rect 31953 31773 31987 31807
rect 32137 31773 32171 31807
rect 32321 31773 32355 31807
rect 32965 31773 32999 31807
rect 1593 31705 1627 31739
rect 46673 31705 46707 31739
rect 18337 31637 18371 31671
rect 21833 31637 21867 31671
rect 25973 31637 26007 31671
rect 30297 31637 30331 31671
rect 2237 31433 2271 31467
rect 19533 31433 19567 31467
rect 21281 31433 21315 31467
rect 22661 31433 22695 31467
rect 23597 31433 23631 31467
rect 23765 31433 23799 31467
rect 24593 31433 24627 31467
rect 25237 31433 25271 31467
rect 27905 31433 27939 31467
rect 29285 31433 29319 31467
rect 18061 31365 18095 31399
rect 21925 31365 21959 31399
rect 23397 31365 23431 31399
rect 24225 31365 24259 31399
rect 24425 31365 24459 31399
rect 27077 31365 27111 31399
rect 27261 31365 27295 31399
rect 2145 31297 2179 31331
rect 14473 31297 14507 31331
rect 15301 31297 15335 31331
rect 15485 31297 15519 31331
rect 17141 31297 17175 31331
rect 20545 31297 20579 31331
rect 20729 31297 20763 31331
rect 21097 31297 21131 31331
rect 22569 31297 22603 31331
rect 25145 31297 25179 31331
rect 25789 31297 25823 31331
rect 28089 31297 28123 31331
rect 28181 31297 28215 31331
rect 28457 31297 28491 31331
rect 28917 31297 28951 31331
rect 29101 31297 29135 31331
rect 29929 31297 29963 31331
rect 32137 31297 32171 31331
rect 32321 31297 32355 31331
rect 32689 31297 32723 31331
rect 14565 31229 14599 31263
rect 14841 31229 14875 31263
rect 17785 31229 17819 31263
rect 20821 31229 20855 31263
rect 20913 31229 20947 31263
rect 25881 31229 25915 31263
rect 28365 31229 28399 31263
rect 30205 31229 30239 31263
rect 32413 31229 32447 31263
rect 32505 31229 32539 31263
rect 17325 31161 17359 31195
rect 22109 31161 22143 31195
rect 15301 31093 15335 31127
rect 23581 31093 23615 31127
rect 24409 31093 24443 31127
rect 30021 31093 30055 31127
rect 30113 31093 30147 31127
rect 32873 31093 32907 31127
rect 16037 30889 16071 30923
rect 17877 30889 17911 30923
rect 19349 30889 19383 30923
rect 21005 30889 21039 30923
rect 27445 30889 27479 30923
rect 29745 30889 29779 30923
rect 30757 30889 30791 30923
rect 31125 30889 31159 30923
rect 28733 30821 28767 30855
rect 14289 30753 14323 30787
rect 20821 30753 20855 30787
rect 23305 30753 23339 30787
rect 25973 30753 26007 30787
rect 26249 30753 26283 30787
rect 30849 30753 30883 30787
rect 32229 30753 32263 30787
rect 17049 30685 17083 30719
rect 17233 30685 17267 30719
rect 17877 30685 17911 30719
rect 18061 30685 18095 30719
rect 19257 30685 19291 30719
rect 20729 30685 20763 30719
rect 23029 30685 23063 30719
rect 25881 30685 25915 30719
rect 26709 30685 26743 30719
rect 26893 30685 26927 30719
rect 27353 30685 27387 30719
rect 29009 30685 29043 30719
rect 29561 30685 29595 30719
rect 30573 30685 30607 30719
rect 31953 30685 31987 30719
rect 14565 30617 14599 30651
rect 28733 30617 28767 30651
rect 17417 30549 17451 30583
rect 26801 30549 26835 30583
rect 28917 30549 28951 30583
rect 33701 30549 33735 30583
rect 15485 30345 15519 30379
rect 25145 30345 25179 30379
rect 25881 30345 25915 30379
rect 31125 30345 31159 30379
rect 16037 30277 16071 30311
rect 27077 30277 27111 30311
rect 28457 30277 28491 30311
rect 29653 30277 29687 30311
rect 32965 30277 32999 30311
rect 14841 30209 14875 30243
rect 14934 30209 14968 30243
rect 15117 30209 15151 30243
rect 15209 30209 15243 30243
rect 15347 30209 15381 30243
rect 15945 30209 15979 30243
rect 17325 30209 17359 30243
rect 17509 30209 17543 30243
rect 17601 30209 17635 30243
rect 18797 30209 18831 30243
rect 20729 30209 20763 30243
rect 20913 30209 20947 30243
rect 23949 30209 23983 30243
rect 24317 30209 24351 30243
rect 24961 30209 24995 30243
rect 25697 30209 25731 30243
rect 27721 30209 27755 30243
rect 28641 30209 28675 30243
rect 32873 30209 32907 30243
rect 28825 30141 28859 30175
rect 28917 30141 28951 30175
rect 29377 30141 29411 30175
rect 34345 30141 34379 30175
rect 34529 30141 34563 30175
rect 34897 30141 34931 30175
rect 18981 30073 19015 30107
rect 27261 30073 27295 30107
rect 17141 30005 17175 30039
rect 20821 30005 20855 30039
rect 24317 30005 24351 30039
rect 24501 30005 24535 30039
rect 27905 30005 27939 30039
rect 17877 29801 17911 29835
rect 20913 29801 20947 29835
rect 21925 29801 21959 29835
rect 29561 29801 29595 29835
rect 30665 29801 30699 29835
rect 34805 29801 34839 29835
rect 25053 29733 25087 29767
rect 16129 29665 16163 29699
rect 25789 29665 25823 29699
rect 47593 29665 47627 29699
rect 18337 29597 18371 29631
rect 20177 29597 20211 29631
rect 20821 29597 20855 29631
rect 21005 29597 21039 29631
rect 21741 29597 21775 29631
rect 22017 29597 22051 29631
rect 22937 29597 22971 29631
rect 23673 29597 23707 29631
rect 24869 29597 24903 29631
rect 29745 29597 29779 29631
rect 29837 29597 29871 29631
rect 30021 29597 30055 29631
rect 30113 29597 30147 29631
rect 30573 29597 30607 29631
rect 34713 29597 34747 29631
rect 47317 29597 47351 29631
rect 16405 29529 16439 29563
rect 18429 29529 18463 29563
rect 26065 29529 26099 29563
rect 20269 29461 20303 29495
rect 21557 29461 21591 29495
rect 23029 29461 23063 29495
rect 23765 29461 23799 29495
rect 27537 29461 27571 29495
rect 17325 29257 17359 29291
rect 21281 29257 21315 29291
rect 22201 29257 22235 29291
rect 25237 29257 25271 29291
rect 26433 29257 26467 29291
rect 27077 29257 27111 29291
rect 22017 29189 22051 29223
rect 26157 29189 26191 29223
rect 16681 29121 16715 29155
rect 16774 29121 16808 29155
rect 16957 29121 16991 29155
rect 17049 29121 17083 29155
rect 17187 29121 17221 29155
rect 21833 29121 21867 29155
rect 22661 29121 22695 29155
rect 25053 29121 25087 29155
rect 25789 29121 25823 29155
rect 25882 29121 25916 29155
rect 26065 29121 26099 29155
rect 26295 29121 26329 29155
rect 26985 29121 27019 29155
rect 28825 29121 28859 29155
rect 19533 29053 19567 29087
rect 19809 29053 19843 29087
rect 22937 29053 22971 29087
rect 24409 29053 24443 29087
rect 32689 29053 32723 29087
rect 32873 29053 32907 29087
rect 33149 29053 33183 29087
rect 28917 28917 28951 28951
rect 21005 28713 21039 28747
rect 21741 28713 21775 28747
rect 22201 28713 22235 28747
rect 23397 28713 23431 28747
rect 30021 28713 30055 28747
rect 30205 28713 30239 28747
rect 30665 28713 30699 28747
rect 32873 28713 32907 28747
rect 36461 28713 36495 28747
rect 17509 28577 17543 28611
rect 22937 28577 22971 28611
rect 29837 28577 29871 28611
rect 31033 28577 31067 28611
rect 16497 28509 16531 28543
rect 16589 28509 16623 28543
rect 17417 28509 17451 28543
rect 20361 28509 20395 28543
rect 20509 28509 20543 28543
rect 20826 28509 20860 28543
rect 21649 28509 21683 28543
rect 21925 28509 21959 28543
rect 22661 28509 22695 28543
rect 22845 28509 22879 28543
rect 23029 28509 23063 28543
rect 23213 28509 23247 28543
rect 30021 28509 30055 28543
rect 30849 28509 30883 28543
rect 31125 28509 31159 28543
rect 32781 28509 32815 28543
rect 34713 28509 34747 28543
rect 47685 28509 47719 28543
rect 20637 28441 20671 28475
rect 20729 28441 20763 28475
rect 29745 28441 29779 28475
rect 34989 28441 35023 28475
rect 16773 28373 16807 28407
rect 17785 28373 17819 28407
rect 20453 28169 20487 28203
rect 24501 28169 24535 28203
rect 26341 28169 26375 28203
rect 26985 28169 27019 28203
rect 28365 28169 28399 28203
rect 33701 28169 33735 28203
rect 35357 28169 35391 28203
rect 24409 28101 24443 28135
rect 29469 28101 29503 28135
rect 29561 28101 29595 28135
rect 17601 28033 17635 28067
rect 17749 28033 17783 28067
rect 17877 28033 17911 28067
rect 17969 28033 18003 28067
rect 18107 28033 18141 28067
rect 20085 28033 20119 28067
rect 20269 28033 20303 28067
rect 21833 28033 21867 28067
rect 21925 28033 21959 28067
rect 23581 28033 23615 28067
rect 26157 28033 26191 28067
rect 26433 28033 26467 28067
rect 27353 28033 27387 28067
rect 28181 28033 28215 28067
rect 29285 28033 29319 28067
rect 29653 28033 29687 28067
rect 30481 28033 30515 28067
rect 33609 28033 33643 28067
rect 34437 28033 34471 28067
rect 35265 28033 35299 28067
rect 47593 28033 47627 28067
rect 27445 27965 27479 27999
rect 27537 27965 27571 27999
rect 30389 27965 30423 27999
rect 34529 27965 34563 27999
rect 34805 27965 34839 27999
rect 23765 27897 23799 27931
rect 18245 27829 18279 27863
rect 21833 27829 21867 27863
rect 22201 27829 22235 27863
rect 25973 27829 26007 27863
rect 29837 27829 29871 27863
rect 30757 27829 30791 27863
rect 47685 27829 47719 27863
rect 31677 27625 31711 27659
rect 26617 27557 26651 27591
rect 15577 27489 15611 27523
rect 20177 27489 20211 27523
rect 29929 27489 29963 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 15117 27421 15151 27455
rect 19901 27421 19935 27455
rect 20085 27421 20119 27455
rect 20269 27421 20303 27455
rect 20453 27421 20487 27455
rect 21097 27421 21131 27455
rect 21281 27421 21315 27455
rect 24501 27421 24535 27455
rect 24593 27421 24627 27455
rect 27445 27421 27479 27455
rect 28089 27421 28123 27455
rect 28273 27421 28307 27455
rect 29009 27421 29043 27455
rect 32505 27421 32539 27455
rect 33333 27421 33367 27455
rect 15301 27353 15335 27387
rect 26433 27353 26467 27387
rect 28181 27353 28215 27387
rect 28733 27353 28767 27387
rect 30205 27353 30239 27387
rect 20637 27285 20671 27319
rect 21189 27285 21223 27319
rect 24777 27285 24811 27319
rect 27537 27285 27571 27319
rect 28831 27285 28865 27319
rect 28917 27285 28951 27319
rect 32505 27285 32539 27319
rect 33425 27285 33459 27319
rect 15393 27081 15427 27115
rect 28733 27081 28767 27115
rect 30205 27081 30239 27115
rect 31217 27081 31251 27115
rect 34069 27081 34103 27115
rect 21833 27013 21867 27047
rect 22845 27013 22879 27047
rect 29285 27013 29319 27047
rect 30573 27013 30607 27047
rect 34529 27013 34563 27047
rect 34729 27013 34763 27047
rect 15301 26945 15335 26979
rect 15945 26945 15979 26979
rect 19901 26945 19935 26979
rect 20637 26945 20671 26979
rect 20821 26945 20855 26979
rect 22017 26945 22051 26979
rect 22661 26945 22695 26979
rect 23673 26945 23707 26979
rect 23857 26945 23891 26979
rect 24501 26945 24535 26979
rect 24593 26945 24627 26979
rect 26985 26945 27019 26979
rect 29469 26945 29503 26979
rect 30389 26945 30423 26979
rect 30665 26945 30699 26979
rect 31125 26945 31159 26979
rect 32321 26945 32355 26979
rect 35357 26945 35391 26979
rect 35541 26945 35575 26979
rect 17233 26877 17267 26911
rect 17509 26877 17543 26911
rect 19717 26877 19751 26911
rect 20177 26877 20211 26911
rect 21005 26877 21039 26911
rect 23029 26877 23063 26911
rect 27261 26877 27295 26911
rect 29653 26877 29687 26911
rect 32597 26877 32631 26911
rect 24041 26809 24075 26843
rect 34897 26809 34931 26843
rect 16037 26741 16071 26775
rect 18981 26741 19015 26775
rect 20085 26741 20119 26775
rect 22109 26741 22143 26775
rect 24685 26741 24719 26775
rect 24869 26741 24903 26775
rect 34713 26741 34747 26775
rect 35357 26741 35391 26775
rect 18613 26537 18647 26571
rect 19520 26537 19554 26571
rect 21005 26537 21039 26571
rect 21833 26537 21867 26571
rect 33149 26537 33183 26571
rect 33885 26537 33919 26571
rect 22017 26469 22051 26503
rect 26617 26469 26651 26503
rect 30113 26469 30147 26503
rect 15025 26401 15059 26435
rect 16497 26401 16531 26435
rect 19257 26401 19291 26435
rect 21649 26401 21683 26435
rect 24409 26401 24443 26435
rect 24685 26401 24719 26435
rect 24894 26401 24928 26435
rect 26709 26401 26743 26435
rect 27537 26401 27571 26435
rect 32873 26401 32907 26435
rect 34989 26401 35023 26435
rect 36461 26401 36495 26435
rect 39313 26401 39347 26435
rect 14841 26333 14875 26367
rect 18521 26333 18555 26367
rect 21833 26333 21867 26367
rect 23489 26333 23523 26367
rect 23581 26333 23615 26367
rect 23673 26333 23707 26367
rect 23857 26333 23891 26367
rect 26157 26333 26191 26367
rect 26341 26333 26375 26367
rect 28181 26333 28215 26367
rect 29009 26333 29043 26367
rect 29561 26333 29595 26367
rect 29745 26333 29779 26367
rect 29929 26333 29963 26367
rect 32781 26333 32815 26367
rect 33885 26333 33919 26367
rect 34161 26333 34195 26367
rect 34713 26333 34747 26367
rect 37473 26333 37507 26367
rect 21557 26265 21591 26299
rect 23213 26265 23247 26299
rect 24777 26265 24811 26299
rect 27353 26265 27387 26299
rect 28641 26265 28675 26299
rect 28825 26265 28859 26299
rect 29837 26265 29871 26299
rect 34069 26265 34103 26299
rect 37657 26265 37691 26299
rect 25053 26197 25087 26231
rect 27997 26197 28031 26231
rect 19349 25993 19383 26027
rect 20269 25993 20303 26027
rect 24317 25993 24351 26027
rect 30113 25993 30147 26027
rect 33793 25993 33827 26027
rect 34897 25993 34931 26027
rect 35725 25993 35759 26027
rect 24961 25925 24995 25959
rect 25053 25925 25087 25959
rect 28641 25925 28675 25959
rect 34345 25925 34379 25959
rect 34529 25925 34563 25959
rect 12265 25857 12299 25891
rect 19257 25857 19291 25891
rect 19901 25857 19935 25891
rect 20085 25857 20119 25891
rect 22569 25857 22603 25891
rect 24777 25857 24811 25891
rect 25145 25857 25179 25891
rect 28365 25857 28399 25891
rect 33609 25857 33643 25891
rect 34621 25857 34655 25891
rect 34713 25857 34747 25891
rect 35633 25857 35667 25891
rect 44925 25857 44959 25891
rect 12357 25789 12391 25823
rect 16681 25789 16715 25823
rect 16865 25789 16899 25823
rect 17141 25789 17175 25823
rect 22845 25789 22879 25823
rect 12633 25721 12667 25755
rect 20085 25653 20119 25687
rect 25329 25653 25363 25687
rect 45017 25653 45051 25687
rect 47777 25653 47811 25687
rect 12725 25449 12759 25483
rect 19441 25449 19475 25483
rect 21465 25449 21499 25483
rect 21649 25449 21683 25483
rect 23305 25449 23339 25483
rect 26525 25449 26559 25483
rect 29653 25449 29687 25483
rect 32781 25449 32815 25483
rect 37933 25449 37967 25483
rect 20177 25381 20211 25415
rect 16681 25313 16715 25347
rect 21557 25313 21591 25347
rect 24777 25313 24811 25347
rect 39957 25313 39991 25347
rect 41797 25313 41831 25347
rect 45477 25313 45511 25347
rect 46857 25313 46891 25347
rect 11989 25245 12023 25279
rect 12633 25245 12667 25279
rect 12817 25245 12851 25279
rect 14105 25245 14139 25279
rect 16221 25245 16255 25279
rect 19257 25245 19291 25279
rect 19993 25245 20027 25279
rect 21373 25245 21407 25279
rect 21741 25245 21775 25279
rect 23489 25245 23523 25279
rect 23581 25245 23615 25279
rect 23765 25245 23799 25279
rect 23857 25245 23891 25279
rect 29561 25245 29595 25279
rect 32597 25245 32631 25279
rect 37197 25245 37231 25279
rect 37841 25245 37875 25279
rect 45293 25245 45327 25279
rect 47777 25245 47811 25279
rect 1869 25177 1903 25211
rect 16405 25177 16439 25211
rect 25053 25177 25087 25211
rect 40141 25177 40175 25211
rect 2145 25109 2179 25143
rect 12081 25109 12115 25143
rect 14197 25109 14231 25143
rect 21097 25109 21131 25143
rect 37289 25109 37323 25143
rect 28457 24905 28491 24939
rect 40141 24905 40175 24939
rect 12817 24837 12851 24871
rect 47041 24837 47075 24871
rect 11989 24769 12023 24803
rect 12541 24769 12575 24803
rect 15025 24769 15059 24803
rect 15761 24769 15795 24803
rect 16681 24769 16715 24803
rect 17325 24769 17359 24803
rect 17417 24769 17451 24803
rect 18153 24769 18187 24803
rect 19349 24769 19383 24803
rect 23489 24769 23523 24803
rect 23581 24769 23615 24803
rect 25513 24769 25547 24803
rect 25605 24769 25639 24803
rect 27445 24769 27479 24803
rect 28273 24769 28307 24803
rect 31217 24769 31251 24803
rect 31401 24769 31435 24803
rect 32873 24769 32907 24803
rect 33057 24769 33091 24803
rect 33517 24769 33551 24803
rect 33701 24769 33735 24803
rect 34713 24769 34747 24803
rect 40049 24769 40083 24803
rect 45201 24769 45235 24803
rect 47593 24769 47627 24803
rect 14289 24701 14323 24735
rect 14841 24701 14875 24735
rect 15209 24701 15243 24735
rect 15301 24701 15335 24735
rect 19533 24701 19567 24735
rect 27537 24701 27571 24735
rect 32689 24701 32723 24735
rect 34621 24701 34655 24735
rect 37289 24701 37323 24735
rect 37473 24701 37507 24735
rect 38485 24701 38519 24735
rect 45385 24701 45419 24735
rect 11805 24565 11839 24599
rect 15853 24565 15887 24599
rect 16773 24565 16807 24599
rect 18337 24565 18371 24599
rect 27813 24565 27847 24599
rect 31217 24565 31251 24599
rect 33517 24565 33551 24599
rect 35081 24565 35115 24599
rect 47685 24565 47719 24599
rect 16773 24361 16807 24395
rect 19993 24293 20027 24327
rect 20729 24293 20763 24327
rect 33241 24293 33275 24327
rect 36921 24293 36955 24327
rect 11805 24225 11839 24259
rect 15025 24225 15059 24259
rect 28825 24225 28859 24259
rect 30757 24225 30791 24259
rect 35449 24225 35483 24259
rect 37473 24225 37507 24259
rect 40325 24225 40359 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 14381 24157 14415 24191
rect 14565 24157 14599 24191
rect 17325 24157 17359 24191
rect 19717 24157 19751 24191
rect 19809 24157 19843 24191
rect 20729 24157 20763 24191
rect 21005 24157 21039 24191
rect 21465 24157 21499 24191
rect 25329 24157 25363 24191
rect 26341 24157 26375 24191
rect 26985 24157 27019 24191
rect 29561 24157 29595 24191
rect 30481 24157 30515 24191
rect 32873 24157 32907 24191
rect 33977 24157 34011 24191
rect 35173 24157 35207 24191
rect 39865 24157 39899 24191
rect 12081 24089 12115 24123
rect 15301 24089 15335 24123
rect 26433 24089 26467 24123
rect 27169 24089 27203 24123
rect 32689 24089 32723 24123
rect 33057 24089 33091 24123
rect 37657 24089 37691 24123
rect 39313 24089 39347 24123
rect 40049 24089 40083 24123
rect 13553 24021 13587 24055
rect 14565 24021 14599 24055
rect 17509 24021 17543 24055
rect 20913 24021 20947 24055
rect 21649 24021 21683 24055
rect 25421 24021 25455 24055
rect 29653 24021 29687 24055
rect 32229 24021 32263 24055
rect 32965 24021 32999 24055
rect 34069 24021 34103 24055
rect 1961 23817 1995 23851
rect 12081 23817 12115 23851
rect 13461 23817 13495 23851
rect 14013 23817 14047 23851
rect 14749 23817 14783 23851
rect 15117 23817 15151 23851
rect 20821 23817 20855 23851
rect 21005 23817 21039 23851
rect 23581 23817 23615 23851
rect 29745 23817 29779 23851
rect 30481 23817 30515 23851
rect 33063 23817 33097 23851
rect 35449 23817 35483 23851
rect 36001 23817 36035 23851
rect 37565 23817 37599 23851
rect 39313 23817 39347 23851
rect 47685 23817 47719 23851
rect 14565 23749 14599 23783
rect 20453 23749 20487 23783
rect 28273 23749 28307 23783
rect 31309 23749 31343 23783
rect 32137 23749 32171 23783
rect 32337 23749 32371 23783
rect 32965 23749 32999 23783
rect 33977 23749 34011 23783
rect 1869 23681 1903 23715
rect 11989 23681 12023 23715
rect 12357 23681 12391 23715
rect 12909 23681 12943 23715
rect 13093 23681 13127 23715
rect 13185 23681 13219 23715
rect 13277 23681 13311 23715
rect 13921 23681 13955 23715
rect 14841 23681 14875 23715
rect 14933 23681 14967 23715
rect 15761 23681 15795 23715
rect 17141 23681 17175 23715
rect 19717 23681 19751 23715
rect 19901 23681 19935 23715
rect 19993 23681 20027 23715
rect 20637 23681 20671 23715
rect 20729 23681 20763 23715
rect 21833 23681 21867 23715
rect 25789 23681 25823 23715
rect 27445 23681 27479 23715
rect 30389 23681 30423 23715
rect 31493 23681 31527 23715
rect 31585 23681 31619 23715
rect 33149 23681 33183 23715
rect 33241 23681 33275 23715
rect 35909 23681 35943 23715
rect 37473 23681 37507 23715
rect 39221 23681 39255 23715
rect 42809 23681 42843 23715
rect 42993 23681 43027 23715
rect 45937 23681 45971 23715
rect 47041 23681 47075 23715
rect 47593 23681 47627 23715
rect 12173 23613 12207 23647
rect 15669 23613 15703 23647
rect 22109 23613 22143 23647
rect 27537 23613 27571 23647
rect 27997 23613 28031 23647
rect 33701 23613 33735 23647
rect 16129 23545 16163 23579
rect 31309 23545 31343 23579
rect 32505 23545 32539 23579
rect 12357 23477 12391 23511
rect 17233 23477 17267 23511
rect 19533 23477 19567 23511
rect 25973 23477 26007 23511
rect 32321 23477 32355 23511
rect 42809 23477 42843 23511
rect 45753 23477 45787 23511
rect 46857 23477 46891 23511
rect 12357 23273 12391 23307
rect 17877 23273 17911 23307
rect 22201 23273 22235 23307
rect 23213 23273 23247 23307
rect 29745 23273 29779 23307
rect 31677 23273 31711 23307
rect 33701 23273 33735 23307
rect 34805 23273 34839 23307
rect 42901 23273 42935 23307
rect 48145 23205 48179 23239
rect 16405 23137 16439 23171
rect 20545 23137 20579 23171
rect 24501 23137 24535 23171
rect 27997 23137 28031 23171
rect 38853 23137 38887 23171
rect 39957 23137 39991 23171
rect 45477 23137 45511 23171
rect 46397 23137 46431 23171
rect 12357 23069 12391 23103
rect 12541 23069 12575 23103
rect 15577 23069 15611 23103
rect 15669 23069 15703 23103
rect 16129 23069 16163 23103
rect 18337 23069 18371 23103
rect 19717 23069 19751 23103
rect 20085 23069 20119 23103
rect 20913 23069 20947 23103
rect 21005 23069 21039 23103
rect 21465 23069 21499 23103
rect 22201 23069 22235 23103
rect 22385 23069 22419 23103
rect 23121 23069 23155 23103
rect 26801 23069 26835 23103
rect 29561 23069 29595 23103
rect 30849 23069 30883 23103
rect 31585 23069 31619 23103
rect 33701 23069 33735 23103
rect 34713 23069 34747 23103
rect 37013 23069 37047 23103
rect 38945 23069 38979 23103
rect 42625 23069 42659 23103
rect 42717 23069 42751 23103
rect 43361 23069 43395 23103
rect 43545 23069 43579 23103
rect 45293 23069 45327 23103
rect 19533 23001 19567 23035
rect 24777 23001 24811 23035
rect 26985 23001 27019 23035
rect 40141 23001 40175 23035
rect 41797 23001 41831 23035
rect 47961 23001 47995 23035
rect 18429 22933 18463 22967
rect 19809 22933 19843 22967
rect 19901 22933 19935 22967
rect 20821 22933 20855 22967
rect 21649 22933 21683 22967
rect 26249 22933 26283 22967
rect 31033 22933 31067 22967
rect 37197 22933 37231 22967
rect 39313 22933 39347 22967
rect 43453 22933 43487 22967
rect 16037 22729 16071 22763
rect 16773 22729 16807 22763
rect 19073 22729 19107 22763
rect 19901 22729 19935 22763
rect 20913 22729 20947 22763
rect 23581 22729 23615 22763
rect 24777 22729 24811 22763
rect 25973 22729 26007 22763
rect 27261 22729 27295 22763
rect 40049 22729 40083 22763
rect 48053 22729 48087 22763
rect 19533 22661 19567 22695
rect 19809 22661 19843 22695
rect 22109 22661 22143 22695
rect 24133 22661 24167 22695
rect 38117 22661 38151 22695
rect 11713 22593 11747 22627
rect 13461 22593 13495 22627
rect 15117 22593 15151 22627
rect 15853 22593 15887 22627
rect 16681 22593 16715 22627
rect 19717 22593 19751 22627
rect 20637 22593 20671 22627
rect 20729 22593 20763 22627
rect 21833 22593 21867 22627
rect 24041 22593 24075 22627
rect 24685 22593 24719 22627
rect 25881 22593 25915 22627
rect 27077 22593 27111 22627
rect 27813 22593 27847 22627
rect 31125 22593 31159 22627
rect 32137 22593 32171 22627
rect 33149 22593 33183 22627
rect 33885 22593 33919 22627
rect 35173 22593 35207 22627
rect 37289 22593 37323 22627
rect 39681 22593 39715 22627
rect 40509 22593 40543 22627
rect 41705 22593 41739 22627
rect 41889 22593 41923 22627
rect 42993 22593 43027 22627
rect 44741 22593 44775 22627
rect 47593 22593 47627 22627
rect 11805 22525 11839 22559
rect 17325 22525 17359 22559
rect 17601 22525 17635 22559
rect 31217 22525 31251 22559
rect 39589 22525 39623 22559
rect 42901 22525 42935 22559
rect 43821 22525 43855 22559
rect 45201 22525 45235 22559
rect 45385 22525 45419 22559
rect 46397 22525 46431 22559
rect 44557 22457 44591 22491
rect 12081 22389 12115 22423
rect 13645 22389 13679 22423
rect 15209 22389 15243 22423
rect 20085 22389 20119 22423
rect 27997 22389 28031 22423
rect 31493 22389 31527 22423
rect 32229 22389 32263 22423
rect 33333 22389 33367 22423
rect 34069 22389 34103 22423
rect 34989 22389 35023 22423
rect 40601 22389 40635 22423
rect 40969 22389 41003 22423
rect 41797 22389 41831 22423
rect 47685 22389 47719 22423
rect 11792 22185 11826 22219
rect 17417 22185 17451 22219
rect 31204 22185 31238 22219
rect 34989 22185 35023 22219
rect 35173 22185 35207 22219
rect 35541 22185 35575 22219
rect 40693 22185 40727 22219
rect 45661 22185 45695 22219
rect 45845 22185 45879 22219
rect 42349 22117 42383 22151
rect 13553 22049 13587 22083
rect 15025 22049 15059 22083
rect 15301 22049 15335 22083
rect 19349 22049 19383 22083
rect 19809 22049 19843 22083
rect 30941 22049 30975 22083
rect 32689 22049 32723 22083
rect 34345 22049 34379 22083
rect 46305 22049 46339 22083
rect 46489 22049 46523 22083
rect 46765 22049 46799 22083
rect 11529 21981 11563 22015
rect 14841 21981 14875 22015
rect 17233 21981 17267 22015
rect 19441 21981 19475 22015
rect 24593 21981 24627 22015
rect 25237 21981 25271 22015
rect 27261 21981 27295 22015
rect 27445 21981 27479 22015
rect 28089 21981 28123 22015
rect 29009 21981 29043 22015
rect 29561 21981 29595 22015
rect 32965 21981 32999 22015
rect 34713 21981 34747 22015
rect 37105 21981 37139 22015
rect 39957 21981 39991 22015
rect 40141 21981 40175 22015
rect 40877 21981 40911 22015
rect 42533 21981 42567 22015
rect 42625 21981 42659 22015
rect 44281 21981 44315 22015
rect 44465 21981 44499 22015
rect 45293 21981 45327 22015
rect 45569 21981 45603 22015
rect 33793 21913 33827 21947
rect 36277 21913 36311 21947
rect 37289 21913 37323 21947
rect 38945 21913 38979 21947
rect 40233 21913 40267 21947
rect 42349 21913 42383 21947
rect 24409 21845 24443 21879
rect 25329 21845 25363 21879
rect 27445 21845 27479 21879
rect 28273 21845 28307 21879
rect 28825 21845 28859 21879
rect 29653 21845 29687 21879
rect 36369 21845 36403 21879
rect 44465 21845 44499 21879
rect 11989 21641 12023 21675
rect 13093 21641 13127 21675
rect 22385 21641 22419 21675
rect 36645 21641 36679 21675
rect 45753 21641 45787 21675
rect 14473 21573 14507 21607
rect 24317 21573 24351 21607
rect 28733 21573 28767 21607
rect 33701 21573 33735 21607
rect 35909 21573 35943 21607
rect 37657 21573 37691 21607
rect 45477 21573 45511 21607
rect 45569 21573 45603 21607
rect 47777 21573 47811 21607
rect 11805 21505 11839 21539
rect 13001 21505 13035 21539
rect 16957 21505 16991 21539
rect 17785 21505 17819 21539
rect 18889 21505 18923 21539
rect 22293 21505 22327 21539
rect 23397 21505 23431 21539
rect 27537 21505 27571 21539
rect 28457 21505 28491 21539
rect 32505 21505 32539 21539
rect 35357 21505 35391 21539
rect 35817 21505 35851 21539
rect 36553 21505 36587 21539
rect 42717 21505 42751 21539
rect 42901 21505 42935 21539
rect 43821 21505 43855 21539
rect 44005 21505 44039 21539
rect 45385 21505 45419 21539
rect 46213 21505 46247 21539
rect 47593 21505 47627 21539
rect 14289 21437 14323 21471
rect 14749 21437 14783 21471
rect 23581 21437 23615 21471
rect 24041 21437 24075 21471
rect 30205 21437 30239 21471
rect 32781 21437 32815 21471
rect 33517 21437 33551 21471
rect 46489 21437 46523 21471
rect 45201 21369 45235 21403
rect 47961 21369 47995 21403
rect 17141 21301 17175 21335
rect 17969 21301 18003 21335
rect 18981 21301 19015 21335
rect 25789 21301 25823 21335
rect 27721 21301 27755 21335
rect 38945 21301 38979 21335
rect 42717 21301 42751 21335
rect 43913 21301 43947 21335
rect 44741 21301 44775 21335
rect 42717 21097 42751 21131
rect 24777 21029 24811 21063
rect 25421 21029 25455 21063
rect 11345 20961 11379 20995
rect 16865 20961 16899 20995
rect 22845 20961 22879 20995
rect 24869 20961 24903 20995
rect 25605 20961 25639 20995
rect 25881 20961 25915 20995
rect 27721 20961 27755 20995
rect 31217 20961 31251 20995
rect 33977 20961 34011 20995
rect 46305 20961 46339 20995
rect 48145 20961 48179 20995
rect 10885 20893 10919 20927
rect 13185 20893 13219 20927
rect 14657 20893 14691 20927
rect 15761 20893 15795 20927
rect 16405 20893 16439 20927
rect 19349 20893 19383 20927
rect 20729 20893 20763 20927
rect 22293 20893 22327 20927
rect 25697 20893 25731 20927
rect 25789 20893 25823 20927
rect 26801 20893 26835 20927
rect 26985 20893 27019 20927
rect 27813 20893 27847 20927
rect 28641 20893 28675 20927
rect 29653 20893 29687 20927
rect 33701 20893 33735 20927
rect 37289 20893 37323 20927
rect 38025 20893 38059 20927
rect 42073 20893 42107 20927
rect 42257 20893 42291 20927
rect 42901 20893 42935 20927
rect 42993 20893 43027 20927
rect 43085 20893 43119 20927
rect 43177 20893 43211 20927
rect 43729 20893 43763 20927
rect 43913 20893 43947 20927
rect 45201 20893 45235 20927
rect 45661 20893 45695 20927
rect 11069 20825 11103 20859
rect 15853 20825 15887 20859
rect 16589 20825 16623 20859
rect 21281 20825 21315 20859
rect 24409 20825 24443 20859
rect 31401 20825 31435 20859
rect 33057 20825 33091 20859
rect 34990 20825 35024 20859
rect 35081 20825 35115 20859
rect 36001 20825 36035 20859
rect 42165 20825 42199 20859
rect 45753 20825 45787 20859
rect 46489 20825 46523 20859
rect 13277 20757 13311 20791
rect 14933 20757 14967 20791
rect 19441 20757 19475 20791
rect 27169 20757 27203 20791
rect 28181 20757 28215 20791
rect 28825 20757 28859 20791
rect 29745 20757 29779 20791
rect 43821 20757 43855 20791
rect 45017 20757 45051 20791
rect 10885 20553 10919 20587
rect 23397 20553 23431 20587
rect 25973 20553 26007 20587
rect 26985 20553 27019 20587
rect 28089 20553 28123 20587
rect 30297 20553 30331 20587
rect 31401 20553 31435 20587
rect 41889 20553 41923 20587
rect 44281 20553 44315 20587
rect 47685 20553 47719 20587
rect 15393 20485 15427 20519
rect 18981 20485 19015 20519
rect 25789 20485 25823 20519
rect 25881 20485 25915 20519
rect 28825 20485 28859 20519
rect 33885 20485 33919 20519
rect 35541 20485 35575 20519
rect 36461 20485 36495 20519
rect 45385 20485 45419 20519
rect 10793 20417 10827 20451
rect 13737 20417 13771 20451
rect 15301 20417 15335 20451
rect 16773 20417 16807 20451
rect 17509 20417 17543 20451
rect 22293 20417 22327 20451
rect 23213 20417 23247 20451
rect 23949 20417 23983 20451
rect 27169 20417 27203 20451
rect 27721 20417 27755 20451
rect 27905 20417 27939 20451
rect 28549 20417 28583 20451
rect 31309 20417 31343 20451
rect 33517 20417 33551 20451
rect 41705 20417 41739 20451
rect 41889 20417 41923 20451
rect 42993 20417 43027 20451
rect 44373 20417 44407 20451
rect 44557 20417 44591 20451
rect 47593 20417 47627 20451
rect 11529 20349 11563 20383
rect 11805 20349 11839 20383
rect 18797 20349 18831 20383
rect 19533 20349 19567 20383
rect 22477 20349 22511 20383
rect 35449 20349 35483 20383
rect 42901 20349 42935 20383
rect 43545 20349 43579 20383
rect 45201 20349 45235 20383
rect 46397 20349 46431 20383
rect 13277 20281 13311 20315
rect 25605 20281 25639 20315
rect 44097 20281 44131 20315
rect 13737 20213 13771 20247
rect 16957 20213 16991 20247
rect 17509 20213 17543 20247
rect 24041 20213 24075 20247
rect 26157 20213 26191 20247
rect 11621 20009 11655 20043
rect 12357 20009 12391 20043
rect 15577 20009 15611 20043
rect 19533 20009 19567 20043
rect 19717 20009 19751 20043
rect 44005 20009 44039 20043
rect 13277 19941 13311 19975
rect 25329 19941 25363 19975
rect 26341 19941 26375 19975
rect 16957 19873 16991 19907
rect 20361 19873 20395 19907
rect 22017 19873 22051 19907
rect 2053 19805 2087 19839
rect 11805 19805 11839 19839
rect 12357 19805 12391 19839
rect 12541 19805 12575 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 20177 19805 20211 19839
rect 25697 19805 25731 19839
rect 26617 19805 26651 19839
rect 32413 19805 32447 19839
rect 34713 19805 34747 19839
rect 42441 19805 42475 19839
rect 42809 19805 42843 19839
rect 43637 19805 43671 19839
rect 45845 19805 45879 19839
rect 46305 19805 46339 19839
rect 13277 19737 13311 19771
rect 15393 19737 15427 19771
rect 15609 19737 15643 19771
rect 17233 19737 17267 19771
rect 19349 19737 19383 19771
rect 22569 19737 22603 19771
rect 25513 19737 25547 19771
rect 25881 19737 25915 19771
rect 26709 19737 26743 19771
rect 42625 19737 42659 19771
rect 43821 19737 43855 19771
rect 46489 19737 46523 19771
rect 48145 19737 48179 19771
rect 13461 19669 13495 19703
rect 14197 19669 14231 19703
rect 15761 19669 15795 19703
rect 18705 19669 18739 19703
rect 19559 19669 19593 19703
rect 22661 19669 22695 19703
rect 25605 19669 25639 19703
rect 26525 19669 26559 19703
rect 26893 19669 26927 19703
rect 32229 19669 32263 19703
rect 34805 19669 34839 19703
rect 20085 19465 20119 19499
rect 43085 19465 43119 19499
rect 45569 19465 45603 19499
rect 47685 19465 47719 19499
rect 15393 19397 15427 19431
rect 15593 19397 15627 19431
rect 17417 19397 17451 19431
rect 19993 19397 20027 19431
rect 20913 19397 20947 19431
rect 21833 19397 21867 19431
rect 22033 19397 22067 19431
rect 25973 19397 26007 19431
rect 26173 19397 26207 19431
rect 32229 19397 32263 19431
rect 32321 19397 32355 19431
rect 33517 19397 33551 19431
rect 35173 19397 35207 19431
rect 45017 19397 45051 19431
rect 1777 19329 1811 19363
rect 13185 19329 13219 19363
rect 16773 19329 16807 19363
rect 17601 19329 17635 19363
rect 17877 19329 17911 19363
rect 18061 19329 18095 19363
rect 18881 19329 18915 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 21005 19329 21039 19363
rect 21097 19329 21131 19363
rect 22937 19329 22971 19363
rect 23765 19329 23799 19363
rect 42993 19329 43027 19363
rect 43177 19329 43211 19363
rect 44005 19329 44039 19363
rect 45753 19329 45787 19363
rect 46857 19329 46891 19363
rect 47593 19329 47627 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 13461 19261 13495 19295
rect 14933 19261 14967 19295
rect 21281 19261 21315 19295
rect 23029 19261 23063 19295
rect 24041 19261 24075 19295
rect 32505 19261 32539 19295
rect 33333 19261 33367 19295
rect 15761 19193 15795 19227
rect 18981 19193 19015 19227
rect 20729 19193 20763 19227
rect 22201 19193 22235 19227
rect 23305 19193 23339 19227
rect 26341 19193 26375 19227
rect 15577 19125 15611 19159
rect 16865 19125 16899 19159
rect 20269 19125 20303 19159
rect 22017 19125 22051 19159
rect 25513 19125 25547 19159
rect 26157 19125 26191 19159
rect 46397 19125 46431 19159
rect 46949 19125 46983 19159
rect 2237 18921 2271 18955
rect 14105 18921 14139 18955
rect 14657 18921 14691 18955
rect 22385 18921 22419 18955
rect 25973 18921 26007 18955
rect 28917 18921 28951 18955
rect 30757 18921 30791 18955
rect 32597 18921 32631 18955
rect 33333 18921 33367 18955
rect 45845 18921 45879 18955
rect 31861 18853 31895 18887
rect 14749 18785 14783 18819
rect 21097 18785 21131 18819
rect 21557 18785 21591 18819
rect 22017 18785 22051 18819
rect 29929 18785 29963 18819
rect 31309 18785 31343 18819
rect 32873 18785 32907 18819
rect 34713 18785 34747 18819
rect 34897 18785 34931 18819
rect 45293 18785 45327 18819
rect 46305 18785 46339 18819
rect 46489 18785 46523 18819
rect 47041 18785 47075 18819
rect 2145 18717 2179 18751
rect 14230 18717 14264 18751
rect 15393 18717 15427 18751
rect 15669 18717 15703 18751
rect 16313 18717 16347 18751
rect 17601 18717 17635 18751
rect 21189 18717 21223 18751
rect 22201 18717 22235 18751
rect 25421 18717 25455 18751
rect 25881 18717 25915 18751
rect 26893 18717 26927 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 29561 18717 29595 18751
rect 30389 18717 30423 18751
rect 30573 18717 30607 18751
rect 32413 18717 32447 18751
rect 33517 18717 33551 18751
rect 45477 18717 45511 18751
rect 25145 18649 25179 18683
rect 29745 18649 29779 18683
rect 31401 18649 31435 18683
rect 36553 18649 36587 18683
rect 45661 18649 45695 18683
rect 14289 18581 14323 18615
rect 15209 18581 15243 18615
rect 15577 18581 15611 18615
rect 16129 18581 16163 18615
rect 17693 18581 17727 18615
rect 25243 18581 25277 18615
rect 25329 18581 25363 18615
rect 26985 18581 27019 18615
rect 45569 18581 45603 18615
rect 15117 18309 15151 18343
rect 17693 18309 17727 18343
rect 22109 18309 22143 18343
rect 31585 18309 31619 18343
rect 41797 18309 41831 18343
rect 42625 18309 42659 18343
rect 1869 18241 1903 18275
rect 11897 18241 11931 18275
rect 13001 18241 13035 18275
rect 14381 18241 14415 18275
rect 25145 18241 25179 18275
rect 25789 18241 25823 18275
rect 25973 18241 26007 18275
rect 29009 18241 29043 18275
rect 29193 18241 29227 18275
rect 35081 18241 35115 18275
rect 41705 18241 41739 18275
rect 45109 18241 45143 18275
rect 45569 18241 45603 18275
rect 45845 18241 45879 18275
rect 46121 18241 46155 18275
rect 47593 18241 47627 18275
rect 13093 18173 13127 18207
rect 15577 18173 15611 18207
rect 17509 18173 17543 18207
rect 19165 18173 19199 18207
rect 21833 18173 21867 18207
rect 23857 18173 23891 18207
rect 29745 18173 29779 18207
rect 29929 18173 29963 18207
rect 32781 18173 32815 18207
rect 32965 18173 32999 18207
rect 33977 18173 34011 18207
rect 42441 18173 42475 18207
rect 43913 18173 43947 18207
rect 2053 18105 2087 18139
rect 15393 18105 15427 18139
rect 35541 18105 35575 18139
rect 11989 18037 12023 18071
rect 13369 18037 13403 18071
rect 14473 18037 14507 18071
rect 25053 18037 25087 18071
rect 25789 18037 25823 18071
rect 29101 18037 29135 18071
rect 35357 18037 35391 18071
rect 45569 18037 45603 18071
rect 47041 18037 47075 18071
rect 47685 18037 47719 18071
rect 17141 17833 17175 17867
rect 22109 17833 22143 17867
rect 22753 17833 22787 17867
rect 26801 17833 26835 17867
rect 31217 17833 31251 17867
rect 33885 17833 33919 17867
rect 36093 17833 36127 17867
rect 45661 17833 45695 17867
rect 35265 17765 35299 17799
rect 11713 17697 11747 17731
rect 11897 17697 11931 17731
rect 12173 17697 12207 17731
rect 15669 17697 15703 17731
rect 25053 17697 25087 17731
rect 25329 17697 25363 17731
rect 28733 17697 28767 17731
rect 29837 17697 29871 17731
rect 30665 17697 30699 17731
rect 44465 17697 44499 17731
rect 45017 17697 45051 17731
rect 46305 17697 46339 17731
rect 14841 17629 14875 17663
rect 14933 17629 14967 17663
rect 15393 17629 15427 17663
rect 19257 17629 19291 17663
rect 21925 17629 21959 17663
rect 22661 17629 22695 17663
rect 24409 17629 24443 17663
rect 28365 17629 28399 17663
rect 28457 17629 28491 17663
rect 28641 17629 28675 17663
rect 31125 17629 31159 17663
rect 34069 17629 34103 17663
rect 35173 17629 35207 17663
rect 35357 17629 35391 17663
rect 35449 17629 35483 17663
rect 43453 17629 43487 17663
rect 43637 17629 43671 17663
rect 45385 17629 45419 17663
rect 45477 17629 45511 17663
rect 19533 17561 19567 17595
rect 44097 17561 44131 17595
rect 44281 17561 44315 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 21005 17493 21039 17527
rect 24501 17493 24535 17527
rect 28733 17493 28767 17527
rect 43637 17493 43671 17527
rect 16773 17289 16807 17323
rect 17877 17289 17911 17323
rect 21097 17289 21131 17323
rect 26157 17289 26191 17323
rect 28733 17289 28767 17323
rect 13737 17221 13771 17255
rect 20729 17221 20763 17255
rect 20929 17221 20963 17255
rect 23673 17221 23707 17255
rect 28641 17221 28675 17255
rect 35081 17221 35115 17255
rect 44281 17221 44315 17255
rect 45201 17221 45235 17255
rect 11989 17153 12023 17187
rect 16681 17153 16715 17187
rect 17693 17153 17727 17187
rect 21833 17153 21867 17187
rect 23489 17153 23523 17187
rect 26065 17153 26099 17187
rect 27537 17153 27571 17187
rect 27721 17153 27755 17187
rect 28865 17153 28899 17187
rect 29009 17153 29043 17187
rect 29653 17153 29687 17187
rect 30297 17153 30331 17187
rect 45017 17153 45051 17187
rect 47593 17153 47627 17187
rect 13461 17085 13495 17119
rect 18521 17085 18555 17119
rect 18797 17085 18831 17119
rect 20269 17085 20303 17119
rect 25329 17085 25363 17119
rect 27629 17085 27663 17119
rect 29469 17085 29503 17119
rect 34897 17085 34931 17119
rect 36553 17085 36587 17119
rect 43729 17085 43763 17119
rect 45753 17085 45787 17119
rect 28457 17017 28491 17051
rect 2053 16949 2087 16983
rect 12081 16949 12115 16983
rect 15209 16949 15243 16983
rect 20913 16949 20947 16983
rect 21925 16949 21959 16983
rect 29837 16949 29871 16983
rect 30389 16949 30423 16983
rect 47685 16949 47719 16983
rect 17969 16745 18003 16779
rect 19809 16745 19843 16779
rect 24869 16745 24903 16779
rect 25053 16745 25087 16779
rect 25697 16745 25731 16779
rect 28825 16745 28859 16779
rect 25881 16677 25915 16711
rect 27629 16677 27663 16711
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 11713 16609 11747 16643
rect 11897 16609 11931 16643
rect 12449 16609 12483 16643
rect 19533 16609 19567 16643
rect 21189 16609 21223 16643
rect 21373 16609 21407 16643
rect 30665 16609 30699 16643
rect 32321 16609 32355 16643
rect 46305 16609 46339 16643
rect 48145 16609 48179 16643
rect 14105 16541 14139 16575
rect 14197 16541 14231 16575
rect 16221 16541 16255 16575
rect 17877 16541 17911 16575
rect 19441 16541 19475 16575
rect 20269 16541 20303 16575
rect 20545 16541 20579 16575
rect 23673 16541 23707 16575
rect 27629 16541 27663 16575
rect 27813 16541 27847 16575
rect 29653 16541 29687 16575
rect 29837 16541 29871 16575
rect 45569 16541 45603 16575
rect 45753 16541 45787 16575
rect 1593 16473 1627 16507
rect 23029 16473 23063 16507
rect 24685 16473 24719 16507
rect 25513 16473 25547 16507
rect 28457 16473 28491 16507
rect 28641 16473 28675 16507
rect 32505 16473 32539 16507
rect 34161 16473 34195 16507
rect 45661 16473 45695 16507
rect 46489 16473 46523 16507
rect 16313 16405 16347 16439
rect 20367 16405 20401 16439
rect 20453 16405 20487 16439
rect 23765 16405 23799 16439
rect 24895 16405 24929 16439
rect 25723 16405 25757 16439
rect 2145 16201 2179 16235
rect 19993 16201 20027 16235
rect 23581 16201 23615 16235
rect 25881 16201 25915 16235
rect 28641 16201 28675 16235
rect 29193 16201 29227 16235
rect 32413 16201 32447 16235
rect 16037 16133 16071 16167
rect 16865 16133 16899 16167
rect 19349 16133 19383 16167
rect 2053 16065 2087 16099
rect 15945 16065 15979 16099
rect 19257 16065 19291 16099
rect 19901 16065 19935 16099
rect 21189 16065 21223 16099
rect 26985 16065 27019 16099
rect 28457 16065 28491 16099
rect 28641 16065 28675 16099
rect 29101 16065 29135 16099
rect 29285 16065 29319 16099
rect 31401 16065 31435 16099
rect 32321 16065 32355 16099
rect 44005 16065 44039 16099
rect 47777 16065 47811 16099
rect 16681 15997 16715 16031
rect 18521 15997 18555 16031
rect 21281 15997 21315 16031
rect 21833 15997 21867 16031
rect 22109 15997 22143 16031
rect 24133 15997 24167 16031
rect 24409 15997 24443 16031
rect 44189 15997 44223 16031
rect 45845 15997 45879 16031
rect 27077 15861 27111 15895
rect 31493 15861 31527 15895
rect 19625 15657 19659 15691
rect 21833 15657 21867 15691
rect 23029 15657 23063 15691
rect 24869 15657 24903 15691
rect 44097 15657 44131 15691
rect 16313 15521 16347 15555
rect 16589 15521 16623 15555
rect 23857 15521 23891 15555
rect 24685 15521 24719 15555
rect 25513 15521 25547 15555
rect 25973 15521 26007 15555
rect 26709 15521 26743 15555
rect 28181 15521 28215 15555
rect 30389 15521 30423 15555
rect 30573 15521 30607 15555
rect 30849 15521 30883 15555
rect 2053 15453 2087 15487
rect 16129 15453 16163 15487
rect 19625 15453 19659 15487
rect 19809 15453 19843 15487
rect 22017 15453 22051 15487
rect 22293 15453 22327 15487
rect 22477 15453 22511 15487
rect 22937 15453 22971 15487
rect 23765 15453 23799 15487
rect 24593 15453 24627 15487
rect 25605 15453 25639 15487
rect 26433 15453 26467 15487
rect 44005 15453 44039 15487
rect 25973 15113 26007 15147
rect 27169 15113 27203 15147
rect 23765 15045 23799 15079
rect 1777 14977 1811 15011
rect 25881 14977 25915 15011
rect 26985 14977 27019 15011
rect 43637 14977 43671 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 23581 14909 23615 14943
rect 24041 14909 24075 14943
rect 43821 14909 43855 14943
rect 45109 14909 45143 14943
rect 2329 14569 2363 14603
rect 24777 14569 24811 14603
rect 43821 14569 43855 14603
rect 2237 14365 2271 14399
rect 24685 14365 24719 14399
rect 24869 14365 24903 14399
rect 43729 14365 43763 14399
rect 47593 13889 47627 13923
rect 47685 13685 47719 13719
rect 46489 13345 46523 13379
rect 46305 13277 46339 13311
rect 48145 13209 48179 13243
rect 1409 12801 1443 12835
rect 47777 12801 47811 12835
rect 1593 12597 1627 12631
rect 47685 11101 47719 11135
rect 47593 10625 47627 10659
rect 47685 10421 47719 10455
rect 24409 10081 24443 10115
rect 26157 10081 26191 10115
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 24593 9945 24627 9979
rect 24593 9673 24627 9707
rect 24501 9537 24535 9571
rect 47869 9537 47903 9571
rect 48053 9401 48087 9435
rect 47777 8857 47811 8891
rect 47869 8789 47903 8823
rect 44833 8585 44867 8619
rect 45201 8449 45235 8483
rect 45293 8245 45327 8279
rect 45661 8245 45695 8279
rect 46581 7905 46615 7939
rect 45385 7837 45419 7871
rect 45937 7769 45971 7803
rect 46029 7769 46063 7803
rect 45201 7701 45235 7735
rect 47961 7497 47995 7531
rect 45661 7429 45695 7463
rect 46581 7429 46615 7463
rect 48145 7361 48179 7395
rect 45569 7293 45603 7327
rect 42349 6817 42383 6851
rect 47317 6817 47351 6851
rect 47593 6749 47627 6783
rect 41337 6681 41371 6715
rect 41429 6681 41463 6715
rect 40877 6613 40911 6647
rect 41245 6409 41279 6443
rect 48053 6409 48087 6443
rect 42625 6341 42659 6375
rect 41429 6273 41463 6307
rect 47961 6273 47995 6307
rect 42533 6205 42567 6239
rect 42809 6205 42843 6239
rect 40969 5865 41003 5899
rect 41337 5865 41371 5899
rect 40877 5661 40911 5695
rect 38669 5321 38703 5355
rect 37381 5253 37415 5287
rect 37473 5253 37507 5287
rect 39681 5185 39715 5219
rect 47777 5185 47811 5219
rect 38393 5117 38427 5151
rect 47961 5049 47995 5083
rect 39773 4981 39807 5015
rect 47593 4641 47627 4675
rect 7941 4573 7975 4607
rect 8953 4573 8987 4607
rect 15669 4573 15703 4607
rect 16313 4573 16347 4607
rect 20453 4573 20487 4607
rect 21097 4573 21131 4607
rect 21189 4573 21223 4607
rect 21741 4573 21775 4607
rect 22477 4573 22511 4607
rect 39129 4573 39163 4607
rect 39221 4573 39255 4607
rect 39865 4573 39899 4607
rect 46673 4573 46707 4607
rect 47317 4573 47351 4607
rect 15761 4505 15795 4539
rect 40049 4505 40083 4539
rect 41705 4505 41739 4539
rect 9045 4437 9079 4471
rect 16405 4437 16439 4471
rect 20545 4437 20579 4471
rect 21833 4437 21867 4471
rect 22569 4437 22603 4471
rect 46765 4437 46799 4471
rect 21925 4233 21959 4267
rect 22845 4233 22879 4267
rect 40601 4233 40635 4267
rect 27629 4165 27663 4199
rect 37381 4165 37415 4199
rect 37473 4165 37507 4199
rect 38393 4165 38427 4199
rect 39773 4165 39807 4199
rect 46581 4165 46615 4199
rect 47777 4165 47811 4199
rect 2053 4097 2087 4131
rect 7665 4097 7699 4131
rect 12081 4097 12115 4131
rect 13737 4097 13771 4131
rect 14381 4097 14415 4131
rect 15025 4097 15059 4131
rect 15669 4097 15703 4131
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 17969 4097 18003 4131
rect 18613 4097 18647 4131
rect 19257 4097 19291 4131
rect 19901 4097 19935 4131
rect 20545 4097 20579 4131
rect 21833 4097 21867 4131
rect 22753 4097 22787 4131
rect 23581 4097 23615 4131
rect 36737 4097 36771 4131
rect 39129 4097 39163 4131
rect 39957 4097 39991 4131
rect 40141 4097 40175 4131
rect 40785 4097 40819 4131
rect 41245 4097 41279 4131
rect 41337 4097 41371 4131
rect 42441 4097 42475 4131
rect 7849 4029 7883 4063
rect 9137 4029 9171 4063
rect 27537 4029 27571 4063
rect 28549 4029 28583 4063
rect 39221 4029 39255 4063
rect 47961 3961 47995 3995
rect 2145 3893 2179 3927
rect 2881 3893 2915 3927
rect 10149 3893 10183 3927
rect 12173 3893 12207 3927
rect 13829 3893 13863 3927
rect 14473 3893 14507 3927
rect 15117 3893 15151 3927
rect 15761 3893 15795 3927
rect 16773 3893 16807 3927
rect 17417 3893 17451 3927
rect 18061 3893 18095 3927
rect 18705 3893 18739 3927
rect 19349 3893 19383 3927
rect 19993 3893 20027 3927
rect 20637 3893 20671 3927
rect 23673 3893 23707 3927
rect 36553 3893 36587 3927
rect 42533 3893 42567 3927
rect 46029 3893 46063 3927
rect 46673 3893 46707 3927
rect 17325 3689 17359 3723
rect 18613 3689 18647 3723
rect 20821 3689 20855 3723
rect 27905 3689 27939 3723
rect 16681 3621 16715 3655
rect 3985 3553 4019 3587
rect 9229 3553 9263 3587
rect 9689 3553 9723 3587
rect 14289 3553 14323 3587
rect 14565 3553 14599 3587
rect 17969 3553 18003 3587
rect 22937 3553 22971 3587
rect 33793 3553 33827 3587
rect 46305 3553 46339 3587
rect 2697 3485 2731 3519
rect 6929 3485 6963 3519
rect 7389 3485 7423 3519
rect 8033 3485 8067 3519
rect 11713 3485 11747 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 16589 3485 16623 3519
rect 17233 3485 17267 3519
rect 17877 3485 17911 3519
rect 18521 3485 18555 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 20729 3485 20763 3519
rect 22293 3485 22327 3519
rect 22661 3485 22695 3519
rect 23765 3485 23799 3519
rect 24685 3485 24719 3519
rect 25513 3485 25547 3519
rect 27629 3485 27663 3519
rect 32965 3485 32999 3519
rect 40417 3485 40451 3519
rect 40877 3485 40911 3519
rect 43361 3485 43395 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 1869 3417 1903 3451
rect 2237 3417 2271 3451
rect 9413 3417 9447 3451
rect 24777 3417 24811 3451
rect 41061 3417 41095 3451
rect 42717 3417 42751 3451
rect 45753 3417 45787 3451
rect 46489 3417 46523 3451
rect 48145 3417 48179 3451
rect 2789 3349 2823 3383
rect 7481 3349 7515 3383
rect 8125 3349 8159 3383
rect 19533 3349 19567 3383
rect 28089 3349 28123 3383
rect 33057 3349 33091 3383
rect 40233 3349 40267 3383
rect 14933 3145 14967 3179
rect 15577 3145 15611 3179
rect 16773 3145 16807 3179
rect 17417 3145 17451 3179
rect 18889 3145 18923 3179
rect 36737 3145 36771 3179
rect 39865 3145 39899 3179
rect 41061 3145 41095 3179
rect 48053 3145 48087 3179
rect 2053 3077 2087 3111
rect 7481 3077 7515 3111
rect 10057 3077 10091 3111
rect 11713 3077 11747 3111
rect 19625 3077 19659 3111
rect 22937 3077 22971 3111
rect 25329 3077 25363 3111
rect 27537 3077 27571 3111
rect 27629 3077 27663 3111
rect 28549 3077 28583 3111
rect 33057 3077 33091 3111
rect 42625 3077 42659 3111
rect 45385 3077 45419 3111
rect 1869 3009 1903 3043
rect 7297 3009 7331 3043
rect 9965 3009 9999 3043
rect 11529 3009 11563 3043
rect 14013 3009 14047 3043
rect 14841 3009 14875 3043
rect 15485 3009 15519 3043
rect 16681 3009 16715 3043
rect 17325 3009 17359 3043
rect 18797 3009 18831 3043
rect 21833 3009 21867 3043
rect 21925 3009 21959 3043
rect 22753 3009 22787 3043
rect 25145 3009 25179 3043
rect 29193 3009 29227 3043
rect 32873 3009 32907 3043
rect 36277 3009 36311 3043
rect 39221 3009 39255 3043
rect 41705 3009 41739 3043
rect 42441 3009 42475 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2329 2941 2363 2975
rect 7757 2941 7791 2975
rect 12265 2941 12299 2975
rect 13921 2941 13955 2975
rect 14381 2941 14415 2975
rect 19441 2941 19475 2975
rect 20361 2941 20395 2975
rect 23213 2941 23247 2975
rect 33517 2941 33551 2975
rect 39405 2941 39439 2975
rect 40417 2941 40451 2975
rect 40601 2941 40635 2975
rect 43177 2941 43211 2975
rect 47041 2941 47075 2975
rect 6837 2805 6871 2839
rect 29009 2805 29043 2839
rect 36369 2805 36403 2839
rect 41521 2805 41555 2839
rect 5273 2601 5307 2635
rect 14657 2601 14691 2635
rect 19901 2601 19935 2635
rect 20913 2601 20947 2635
rect 22385 2601 22419 2635
rect 23397 2601 23431 2635
rect 28641 2601 28675 2635
rect 35541 2601 35575 2635
rect 36369 2601 36403 2635
rect 40233 2601 40267 2635
rect 40509 2601 40543 2635
rect 41153 2601 41187 2635
rect 17325 2533 17359 2567
rect 30205 2533 30239 2567
rect 38301 2533 38335 2567
rect 41705 2533 41739 2567
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2881 2465 2915 2499
rect 6561 2465 6595 2499
rect 7021 2465 7055 2499
rect 9689 2465 9723 2499
rect 24593 2465 24627 2499
rect 24777 2465 24811 2499
rect 25145 2465 25179 2499
rect 27261 2465 27295 2499
rect 39313 2465 39347 2499
rect 40233 2465 40267 2499
rect 43913 2465 43947 2499
rect 46489 2465 46523 2499
rect 47869 2465 47903 2499
rect 3801 2397 3835 2431
rect 5457 2397 5491 2431
rect 14565 2397 14599 2431
rect 15301 2397 15335 2431
rect 15577 2397 15611 2431
rect 19809 2397 19843 2431
rect 23581 2397 23615 2431
rect 26985 2397 27019 2431
rect 28457 2397 28491 2431
rect 30849 2397 30883 2431
rect 35725 2397 35759 2431
rect 38117 2397 38151 2431
rect 39957 2397 39991 2431
rect 41889 2397 41923 2431
rect 43637 2397 43671 2431
rect 46213 2397 46247 2431
rect 47685 2397 47719 2431
rect 6745 2329 6779 2363
rect 9413 2329 9447 2363
rect 17141 2329 17175 2363
rect 20821 2329 20855 2363
rect 22293 2329 22327 2363
rect 30021 2329 30055 2363
rect 36277 2329 36311 2363
rect 39129 2329 39163 2363
rect 41061 2329 41095 2363
rect 45385 2329 45419 2363
rect 3985 2261 4019 2295
rect 30665 2261 30699 2295
rect 45477 2261 45511 2295
<< metal1 >>
rect 12618 47404 12624 47456
rect 12676 47444 12682 47456
rect 15838 47444 15844 47456
rect 12676 47416 15844 47444
rect 12676 47404 12682 47416
rect 15838 47404 15844 47416
rect 15896 47404 15902 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 40586 47240 40592 47252
rect 2056 47212 40592 47240
rect 2056 47113 2084 47212
rect 40586 47200 40592 47212
rect 40644 47200 40650 47252
rect 3053 47175 3111 47181
rect 3053 47141 3065 47175
rect 3099 47172 3111 47175
rect 3099 47144 26234 47172
rect 3099 47141 3111 47144
rect 3053 47135 3111 47141
rect 2041 47107 2099 47113
rect 2041 47073 2053 47107
rect 2087 47073 2099 47107
rect 2041 47067 2099 47073
rect 12250 47064 12256 47116
rect 12308 47104 12314 47116
rect 12345 47107 12403 47113
rect 12345 47104 12357 47107
rect 12308 47076 12357 47104
rect 12308 47064 12314 47076
rect 12345 47073 12357 47076
rect 12391 47073 12403 47107
rect 12618 47104 12624 47116
rect 12579 47076 12624 47104
rect 12345 47067 12403 47073
rect 12618 47064 12624 47076
rect 12676 47064 12682 47116
rect 13814 47064 13820 47116
rect 13872 47104 13878 47116
rect 16945 47107 17003 47113
rect 13872 47076 14964 47104
rect 13872 47064 13878 47076
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47036 1823 47039
rect 1946 47036 1952 47048
rect 1811 47008 1952 47036
rect 1811 47005 1823 47008
rect 1765 46999 1823 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4798 47036 4804 47048
rect 4759 47008 4804 47036
rect 3789 46999 3847 47005
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 5868 47008 6377 47036
rect 5868 46996 5874 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 7282 47036 7288 47048
rect 7243 47008 7288 47036
rect 6365 46999 6423 47005
rect 7282 46996 7288 47008
rect 7340 46996 7346 47048
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 14936 47045 14964 47076
rect 15212 47076 16896 47104
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 9401 46999 9459 47005
rect 14093 47039 14151 47045
rect 14093 47005 14105 47039
rect 14139 47005 14151 47039
rect 14093 46999 14151 47005
rect 14921 47039 14979 47045
rect 14921 47005 14933 47039
rect 14967 47005 14979 47039
rect 14921 46999 14979 47005
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 2777 46931 2835 46937
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 2792 46900 2820 46931
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 6638 46968 6644 46980
rect 6599 46940 6644 46968
rect 6638 46928 6644 46940
rect 6696 46928 6702 46980
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 9585 46931 9643 46937
rect 4890 46900 4896 46912
rect 2648 46872 2820 46900
rect 4851 46872 4896 46900
rect 2648 46860 2654 46872
rect 4890 46860 4896 46872
rect 4948 46860 4954 46912
rect 7466 46900 7472 46912
rect 7427 46872 7472 46900
rect 7466 46860 7472 46872
rect 7524 46860 7530 46912
rect 12894 46860 12900 46912
rect 12952 46900 12958 46912
rect 14108 46900 14136 46999
rect 14292 46940 14964 46968
rect 14292 46909 14320 46940
rect 12952 46872 14136 46900
rect 14277 46903 14335 46909
rect 12952 46860 12958 46872
rect 14277 46869 14289 46903
rect 14323 46869 14335 46903
rect 14936 46900 14964 46940
rect 15010 46928 15016 46980
rect 15068 46968 15074 46980
rect 15105 46971 15163 46977
rect 15105 46968 15117 46971
rect 15068 46940 15117 46968
rect 15068 46928 15074 46940
rect 15105 46937 15117 46940
rect 15151 46937 15163 46971
rect 15105 46931 15163 46937
rect 15212 46900 15240 47076
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 16868 46968 16896 47076
rect 16945 47073 16957 47107
rect 16991 47104 17003 47107
rect 21174 47104 21180 47116
rect 16991 47076 21180 47104
rect 16991 47073 17003 47076
rect 16945 47067 17003 47073
rect 21174 47064 21180 47076
rect 21232 47064 21238 47116
rect 26206 47104 26234 47144
rect 29086 47132 29092 47184
rect 29144 47172 29150 47184
rect 29917 47175 29975 47181
rect 29917 47172 29929 47175
rect 29144 47144 29929 47172
rect 29144 47132 29150 47144
rect 29917 47141 29929 47144
rect 29963 47141 29975 47175
rect 29917 47135 29975 47141
rect 30374 47132 30380 47184
rect 30432 47172 30438 47184
rect 31021 47175 31079 47181
rect 31021 47172 31033 47175
rect 30432 47144 31033 47172
rect 30432 47132 30438 47144
rect 31021 47141 31033 47144
rect 31067 47141 31079 47175
rect 31021 47135 31079 47141
rect 47949 47175 48007 47181
rect 47949 47141 47961 47175
rect 47995 47172 48007 47175
rect 48038 47172 48044 47184
rect 47995 47144 48044 47172
rect 47995 47141 48007 47144
rect 47949 47135 48007 47141
rect 48038 47132 48044 47144
rect 48096 47132 48102 47184
rect 35434 47104 35440 47116
rect 26206 47076 35440 47104
rect 35434 47064 35440 47076
rect 35492 47064 35498 47116
rect 43162 47104 43168 47116
rect 43123 47076 43168 47104
rect 43162 47064 43168 47076
rect 43220 47064 43226 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 18690 46996 18696 47048
rect 18748 47036 18754 47048
rect 19245 47039 19303 47045
rect 19245 47036 19257 47039
rect 18748 47008 19257 47036
rect 18748 46996 18754 47008
rect 19245 47005 19257 47008
rect 19291 47005 19303 47039
rect 20346 47036 20352 47048
rect 19245 46999 19303 47005
rect 19352 47008 20352 47036
rect 19352 46968 19380 47008
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 20898 47036 20904 47048
rect 20859 47008 20904 47036
rect 20898 46996 20904 47008
rect 20956 46996 20962 47048
rect 22005 47039 22063 47045
rect 22005 47036 22017 47039
rect 21008 47008 22017 47036
rect 19518 46968 19524 46980
rect 16868 46940 19380 46968
rect 19479 46940 19524 46968
rect 19518 46928 19524 46940
rect 19576 46928 19582 46980
rect 14936 46872 15240 46900
rect 14277 46863 14335 46869
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 21008 46900 21036 47008
rect 22005 47005 22017 47008
rect 22051 47005 22063 47039
rect 24854 47036 24860 47048
rect 24815 47008 24860 47036
rect 22005 46999 22063 47005
rect 24854 46996 24860 47008
rect 24912 46996 24918 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28537 47039 28595 47045
rect 28537 47036 28549 47039
rect 28408 47008 28549 47036
rect 28408 46996 28414 47008
rect 28537 47005 28549 47008
rect 28583 47005 28595 47039
rect 28537 46999 28595 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 30926 46996 30932 47048
rect 30984 47036 30990 47048
rect 31205 47039 31263 47045
rect 31205 47036 31217 47039
rect 30984 47008 31217 47036
rect 30984 46996 30990 47008
rect 31205 47005 31217 47008
rect 31251 47005 31263 47039
rect 31205 46999 31263 47005
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 38381 46999 38439 47005
rect 40218 46996 40224 47048
rect 40276 47036 40282 47048
rect 40497 47039 40555 47045
rect 40497 47036 40509 47039
rect 40276 47008 40509 47036
rect 40276 46996 40282 47008
rect 40497 47005 40509 47008
rect 40543 47005 40555 47039
rect 40497 46999 40555 47005
rect 41877 47039 41935 47045
rect 41877 47005 41889 47039
rect 41923 47036 41935 47039
rect 42613 47039 42671 47045
rect 42613 47036 42625 47039
rect 41923 47008 42625 47036
rect 41923 47005 41935 47008
rect 41877 46999 41935 47005
rect 42613 47005 42625 47008
rect 42659 47005 42671 47039
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 42613 46999 42671 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 28721 46971 28779 46977
rect 28721 46937 28733 46971
rect 28767 46968 28779 46971
rect 28810 46968 28816 46980
rect 28767 46940 28816 46968
rect 28767 46937 28779 46940
rect 28721 46931 28779 46937
rect 28810 46928 28816 46940
rect 28868 46928 28874 46980
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 42797 46971 42855 46977
rect 42797 46937 42809 46971
rect 42843 46968 42855 46971
rect 43162 46968 43168 46980
rect 42843 46940 43168 46968
rect 42843 46937 42855 46940
rect 42797 46931 42855 46937
rect 21818 46900 21824 46912
rect 20036 46872 21036 46900
rect 21779 46872 21824 46900
rect 20036 46860 20042 46872
rect 21818 46860 21824 46872
rect 21876 46860 21882 46912
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 43162 46928 43168 46940
rect 43220 46928 43226 46980
rect 45370 46968 45376 46980
rect 45331 46940 45376 46968
rect 45370 46928 45376 46940
rect 45428 46928 45434 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 41230 46860 41236 46912
rect 41288 46900 41294 46912
rect 41782 46900 41788 46912
rect 41288 46872 41788 46900
rect 41288 46860 41294 46872
rect 41782 46860 41788 46872
rect 41840 46860 41846 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 3878 46588 3884 46640
rect 3936 46628 3942 46640
rect 5813 46631 5871 46637
rect 5813 46628 5825 46631
rect 3936 46600 5825 46628
rect 3936 46588 3942 46600
rect 5813 46597 5825 46600
rect 5859 46597 5871 46631
rect 5813 46591 5871 46597
rect 10962 46588 10968 46640
rect 11020 46628 11026 46640
rect 13357 46631 13415 46637
rect 13357 46628 13369 46631
rect 11020 46600 13369 46628
rect 11020 46588 11026 46600
rect 13357 46597 13369 46600
rect 13403 46597 13415 46631
rect 24854 46628 24860 46640
rect 13357 46591 13415 46597
rect 24596 46600 24860 46628
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 24596 46569 24624 46600
rect 24854 46588 24860 46600
rect 24912 46588 24918 46640
rect 24581 46563 24639 46569
rect 24581 46529 24593 46563
rect 24627 46529 24639 46563
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 24581 46523 24639 46529
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 47946 46560 47952 46572
rect 47907 46532 47952 46560
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 3970 46492 3976 46504
rect 3931 46464 3976 46492
rect 3970 46452 3976 46464
rect 4028 46452 4034 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46492 4215 46495
rect 5350 46492 5356 46504
rect 4203 46464 5356 46492
rect 4203 46461 4215 46464
rect 4157 46455 4215 46461
rect 5350 46452 5356 46464
rect 5408 46452 5414 46504
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11517 46455 11575 46461
rect 11701 46495 11759 46501
rect 11701 46461 11713 46495
rect 11747 46492 11759 46495
rect 13078 46492 13084 46504
rect 11747 46464 13084 46492
rect 11747 46461 11759 46464
rect 11701 46455 11759 46461
rect 13078 46452 13084 46464
rect 13136 46452 13142 46504
rect 13814 46492 13820 46504
rect 13775 46464 13820 46492
rect 13814 46452 13820 46464
rect 13872 46452 13878 46504
rect 14001 46495 14059 46501
rect 14001 46461 14013 46495
rect 14047 46492 14059 46495
rect 14182 46492 14188 46504
rect 14047 46464 14188 46492
rect 14047 46461 14059 46464
rect 14001 46455 14059 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 19429 46495 19487 46501
rect 14332 46464 14377 46492
rect 14332 46452 14338 46464
rect 19429 46461 19441 46495
rect 19475 46461 19487 46495
rect 19429 46455 19487 46461
rect 19613 46495 19671 46501
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 20162 46492 20168 46504
rect 19659 46464 20168 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 19444 46424 19472 46455
rect 20162 46452 20168 46464
rect 20220 46452 20226 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 31573 46495 31631 46501
rect 31573 46461 31585 46495
rect 31619 46492 31631 46495
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 31619 46464 32137 46492
rect 31619 46461 31631 46464
rect 31573 46455 31631 46461
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32306 46492 32312 46504
rect 32267 46464 32312 46492
rect 32125 46455 32183 46461
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46461 32643 46495
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 32585 46455 32643 46461
rect 22005 46427 22063 46433
rect 22005 46424 22017 46427
rect 19444 46396 22017 46424
rect 22005 46393 22017 46396
rect 22051 46393 22063 46427
rect 22005 46387 22063 46393
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 32600 46424 32628 46455
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 42889 46455 42947 46461
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45189 46455 45247 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46658 46492 46664 46504
rect 45419 46464 46664 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 32272 46396 32628 46424
rect 32272 46384 32278 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 42576 46396 42932 46424
rect 45204 46424 45232 46455
rect 46658 46452 46664 46464
rect 46716 46452 46722 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 45462 46424 45468 46436
rect 45204 46396 45468 46424
rect 42576 46384 42582 46396
rect 45462 46384 45468 46396
rect 45520 46384 45526 46436
rect 1486 46316 1492 46368
rect 1544 46356 1550 46368
rect 1581 46359 1639 46365
rect 1581 46356 1593 46359
rect 1544 46328 1593 46356
rect 1544 46316 1550 46328
rect 1581 46325 1593 46328
rect 1627 46325 1639 46359
rect 1581 46319 1639 46325
rect 41233 46359 41291 46365
rect 41233 46325 41245 46359
rect 41279 46356 41291 46359
rect 41322 46356 41328 46368
rect 41279 46328 41328 46356
rect 41279 46325 41291 46328
rect 41233 46319 41291 46325
rect 41322 46316 41328 46328
rect 41380 46316 41386 46368
rect 47762 46316 47768 46368
rect 47820 46356 47826 46368
rect 48041 46359 48099 46365
rect 48041 46356 48053 46359
rect 47820 46328 48053 46356
rect 47820 46316 47826 46328
rect 48041 46325 48053 46328
rect 48087 46325 48099 46359
rect 48041 46319 48099 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3970 46112 3976 46164
rect 4028 46152 4034 46164
rect 4617 46155 4675 46161
rect 4617 46152 4629 46155
rect 4028 46124 4629 46152
rect 4028 46112 4034 46124
rect 4617 46121 4629 46124
rect 4663 46121 4675 46155
rect 5350 46152 5356 46164
rect 5311 46124 5356 46152
rect 4617 46115 4675 46121
rect 5350 46112 5356 46124
rect 5408 46112 5414 46164
rect 13078 46152 13084 46164
rect 13039 46124 13084 46152
rect 13078 46112 13084 46124
rect 13136 46112 13142 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 20162 46152 20168 46164
rect 20123 46124 20168 46152
rect 20162 46112 20168 46124
rect 20220 46112 20226 46164
rect 20714 46152 20720 46164
rect 20272 46124 20720 46152
rect 6886 46056 14044 46084
rect 1762 45908 1768 45960
rect 1820 45948 1826 45960
rect 2041 45951 2099 45957
rect 2041 45948 2053 45951
rect 1820 45920 2053 45948
rect 1820 45908 1826 45920
rect 2041 45917 2053 45920
rect 2087 45917 2099 45951
rect 2041 45911 2099 45917
rect 5261 45951 5319 45957
rect 5261 45917 5273 45951
rect 5307 45948 5319 45951
rect 6886 45948 6914 46056
rect 11606 45976 11612 46028
rect 11664 46016 11670 46028
rect 11701 46019 11759 46025
rect 11701 46016 11713 46019
rect 11664 45988 11713 46016
rect 11664 45976 11670 45988
rect 11701 45985 11713 45988
rect 11747 45985 11759 46019
rect 14016 46016 14044 46056
rect 14090 46044 14096 46096
rect 14148 46084 14154 46096
rect 20272 46084 20300 46124
rect 20714 46112 20720 46124
rect 20772 46112 20778 46164
rect 24762 46152 24768 46164
rect 24723 46124 24768 46152
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 31849 46155 31907 46161
rect 31849 46121 31861 46155
rect 31895 46152 31907 46155
rect 32306 46152 32312 46164
rect 31895 46124 32312 46152
rect 31895 46121 31907 46124
rect 31849 46115 31907 46121
rect 32306 46112 32312 46124
rect 32364 46112 32370 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 14148 46056 20300 46084
rect 20640 46056 31800 46084
rect 14148 46044 14154 46056
rect 20640 46016 20668 46056
rect 14016 45988 20668 46016
rect 20717 46019 20775 46025
rect 11701 45979 11759 45985
rect 20717 45985 20729 46019
rect 20763 46016 20775 46019
rect 20898 46016 20904 46028
rect 20763 45988 20904 46016
rect 20763 45985 20775 45988
rect 20717 45979 20775 45985
rect 20898 45976 20904 45988
rect 20956 45976 20962 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 5307 45920 6914 45948
rect 11977 45951 12035 45957
rect 5307 45917 5319 45920
rect 5261 45911 5319 45917
rect 11977 45917 11989 45951
rect 12023 45917 12035 45951
rect 11977 45911 12035 45917
rect 12989 45951 13047 45957
rect 12989 45917 13001 45951
rect 13035 45948 13047 45951
rect 13906 45948 13912 45960
rect 13035 45920 13912 45948
rect 13035 45917 13047 45920
rect 12989 45911 13047 45917
rect 11992 45880 12020 45911
rect 13906 45908 13912 45920
rect 13964 45908 13970 45960
rect 14090 45948 14096 45960
rect 14051 45920 14096 45948
rect 14090 45908 14096 45920
rect 14148 45908 14154 45960
rect 24688 45957 24716 46056
rect 25317 46019 25375 46025
rect 25317 45985 25329 46019
rect 25363 46016 25375 46019
rect 26234 46016 26240 46028
rect 25363 45988 26240 46016
rect 25363 45985 25375 45988
rect 25317 45979 25375 45985
rect 26234 45976 26240 45988
rect 26292 45976 26298 46028
rect 26697 46019 26755 46025
rect 26697 45985 26709 46019
rect 26743 45985 26755 46019
rect 26697 45979 26755 45985
rect 20073 45951 20131 45957
rect 20073 45917 20085 45951
rect 20119 45917 20131 45951
rect 20073 45911 20131 45917
rect 24673 45951 24731 45957
rect 24673 45917 24685 45951
rect 24719 45917 24731 45951
rect 24673 45911 24731 45917
rect 17310 45880 17316 45892
rect 11992 45852 17316 45880
rect 17310 45840 17316 45852
rect 17368 45840 17374 45892
rect 20088 45824 20116 45911
rect 20898 45880 20904 45892
rect 20859 45852 20904 45880
rect 20898 45840 20904 45852
rect 20956 45840 20962 45892
rect 25498 45880 25504 45892
rect 25459 45852 25504 45880
rect 25498 45840 25504 45852
rect 25556 45840 25562 45892
rect 14090 45772 14096 45824
rect 14148 45812 14154 45824
rect 20070 45812 20076 45824
rect 14148 45784 20076 45812
rect 14148 45772 14154 45784
rect 20070 45772 20076 45784
rect 20128 45772 20134 45824
rect 25774 45772 25780 45824
rect 25832 45812 25838 45824
rect 26712 45812 26740 45979
rect 31772 45960 31800 46056
rect 39390 46044 39396 46096
rect 39448 46084 39454 46096
rect 42978 46084 42984 46096
rect 39448 46056 42984 46084
rect 39448 46044 39454 46056
rect 42978 46044 42984 46056
rect 43036 46044 43042 46096
rect 41322 46016 41328 46028
rect 41283 45988 41328 46016
rect 41322 45976 41328 45988
rect 41380 45976 41386 46028
rect 41874 46016 41880 46028
rect 41835 45988 41880 46016
rect 41874 45976 41880 45988
rect 41932 45976 41938 46028
rect 45830 45976 45836 46028
rect 45888 46016 45894 46028
rect 46293 46019 46351 46025
rect 46293 46016 46305 46019
rect 45888 45988 46305 46016
rect 45888 45976 45894 45988
rect 46293 45985 46305 45988
rect 46339 45985 46351 46019
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 46293 45979 46351 45985
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 31754 45948 31760 45960
rect 31667 45920 31760 45948
rect 31754 45908 31760 45920
rect 31812 45908 31818 45960
rect 38194 45948 38200 45960
rect 38155 45920 38200 45948
rect 38194 45908 38200 45920
rect 38252 45908 38258 45960
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43901 45951 43959 45957
rect 43901 45948 43913 45951
rect 43864 45920 43913 45948
rect 43864 45908 43870 45920
rect 43901 45917 43913 45920
rect 43947 45917 43959 45951
rect 43901 45911 43959 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 41506 45880 41512 45892
rect 41467 45852 41512 45880
rect 41506 45840 41512 45852
rect 41564 45840 41570 45892
rect 45833 45883 45891 45889
rect 45833 45880 45845 45883
rect 43272 45852 45845 45880
rect 25832 45784 26740 45812
rect 25832 45772 25838 45784
rect 31018 45772 31024 45824
rect 31076 45812 31082 45824
rect 43272 45812 43300 45852
rect 45833 45849 45845 45852
rect 45879 45849 45891 45883
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 45833 45843 45891 45849
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 44082 45812 44088 45824
rect 31076 45784 43300 45812
rect 44043 45784 44088 45812
rect 31076 45772 31082 45784
rect 44082 45772 44088 45784
rect 44140 45772 44146 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 20809 45611 20867 45617
rect 20809 45577 20821 45611
rect 20855 45608 20867 45611
rect 20898 45608 20904 45620
rect 20855 45580 20904 45608
rect 20855 45577 20867 45580
rect 20809 45571 20867 45577
rect 20898 45568 20904 45580
rect 20956 45568 20962 45620
rect 24762 45568 24768 45620
rect 24820 45608 24826 45620
rect 25498 45608 25504 45620
rect 24820 45580 25360 45608
rect 25459 45580 25504 45608
rect 24820 45568 24826 45580
rect 25332 45540 25360 45580
rect 25498 45568 25504 45580
rect 25556 45568 25562 45620
rect 31018 45608 31024 45620
rect 25608 45580 31024 45608
rect 25608 45540 25636 45580
rect 31018 45568 31024 45580
rect 31076 45568 31082 45620
rect 31754 45568 31760 45620
rect 31812 45608 31818 45620
rect 39390 45608 39396 45620
rect 31812 45580 39396 45608
rect 31812 45568 31818 45580
rect 39390 45568 39396 45580
rect 39448 45568 39454 45620
rect 41417 45611 41475 45617
rect 41417 45577 41429 45611
rect 41463 45608 41475 45611
rect 41506 45608 41512 45620
rect 41463 45580 41512 45608
rect 41463 45577 41475 45580
rect 41417 45571 41475 45577
rect 41506 45568 41512 45580
rect 41564 45568 41570 45620
rect 42521 45611 42579 45617
rect 42521 45577 42533 45611
rect 42567 45608 42579 45611
rect 42610 45608 42616 45620
rect 42567 45580 42616 45608
rect 42567 45577 42579 45580
rect 42521 45571 42579 45577
rect 42610 45568 42616 45580
rect 42668 45568 42674 45620
rect 45094 45568 45100 45620
rect 45152 45608 45158 45620
rect 45152 45580 45876 45608
rect 45152 45568 45158 45580
rect 43162 45540 43168 45552
rect 25332 45512 25636 45540
rect 43123 45512 43168 45540
rect 43162 45500 43168 45512
rect 43220 45500 43226 45552
rect 43809 45543 43867 45549
rect 43809 45509 43821 45543
rect 43855 45540 43867 45543
rect 44174 45540 44180 45552
rect 43855 45512 44180 45540
rect 43855 45509 43867 45512
rect 43809 45503 43867 45509
rect 44174 45500 44180 45512
rect 44232 45500 44238 45552
rect 45646 45540 45652 45552
rect 44284 45512 45652 45540
rect 1762 45472 1768 45484
rect 1723 45444 1768 45472
rect 1762 45432 1768 45444
rect 1820 45432 1826 45484
rect 13814 45432 13820 45484
rect 13872 45472 13878 45484
rect 13909 45475 13967 45481
rect 13909 45472 13921 45475
rect 13872 45444 13921 45472
rect 13872 45432 13878 45444
rect 13909 45441 13921 45444
rect 13955 45441 13967 45475
rect 20714 45472 20720 45484
rect 20675 45444 20720 45472
rect 13909 45435 13967 45441
rect 20714 45432 20720 45444
rect 20772 45432 20778 45484
rect 25409 45475 25467 45481
rect 25409 45441 25421 45475
rect 25455 45472 25467 45475
rect 38654 45472 38660 45484
rect 25455 45444 38660 45472
rect 25455 45441 25467 45444
rect 25409 45435 25467 45441
rect 38654 45432 38660 45444
rect 38712 45432 38718 45484
rect 41322 45472 41328 45484
rect 41283 45444 41328 45472
rect 41322 45432 41328 45444
rect 41380 45432 41386 45484
rect 42429 45475 42487 45481
rect 42429 45441 42441 45475
rect 42475 45441 42487 45475
rect 43070 45472 43076 45484
rect 43031 45444 43076 45472
rect 42429 45435 42487 45441
rect 1949 45407 2007 45413
rect 1949 45373 1961 45407
rect 1995 45404 2007 45407
rect 2222 45404 2228 45416
rect 1995 45376 2228 45404
rect 1995 45373 2007 45376
rect 1949 45367 2007 45373
rect 2222 45364 2228 45376
rect 2280 45364 2286 45416
rect 2774 45404 2780 45416
rect 2735 45376 2780 45404
rect 2774 45364 2780 45376
rect 2832 45364 2838 45416
rect 26234 45364 26240 45416
rect 26292 45404 26298 45416
rect 42444 45404 42472 45435
rect 43070 45432 43076 45444
rect 43128 45432 43134 45484
rect 44284 45404 44312 45512
rect 45646 45500 45652 45512
rect 45704 45500 45710 45552
rect 44450 45404 44456 45416
rect 26292 45376 26337 45404
rect 42444 45376 44312 45404
rect 44411 45376 44456 45404
rect 26292 45364 26298 45376
rect 44450 45364 44456 45376
rect 44508 45364 44514 45416
rect 44637 45407 44695 45413
rect 44637 45373 44649 45407
rect 44683 45404 44695 45407
rect 45094 45404 45100 45416
rect 44683 45376 45100 45404
rect 44683 45373 44695 45376
rect 44637 45367 44695 45373
rect 45094 45364 45100 45376
rect 45152 45364 45158 45416
rect 45848 45413 45876 45580
rect 46658 45500 46664 45552
rect 46716 45540 46722 45552
rect 47673 45543 47731 45549
rect 47673 45540 47685 45543
rect 46716 45512 47685 45540
rect 46716 45500 46722 45512
rect 47673 45509 47685 45512
rect 47719 45509 47731 45543
rect 47673 45503 47731 45509
rect 46750 45472 46756 45484
rect 46711 45444 46756 45472
rect 46750 45432 46756 45444
rect 46808 45432 46814 45484
rect 47581 45475 47639 45481
rect 47581 45441 47593 45475
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 45833 45407 45891 45413
rect 45833 45373 45845 45407
rect 45879 45373 45891 45407
rect 45833 45367 45891 45373
rect 38194 45296 38200 45348
rect 38252 45336 38258 45348
rect 47596 45336 47624 45435
rect 38252 45308 47624 45336
rect 38252 45296 38258 45308
rect 43898 45268 43904 45280
rect 43859 45240 43904 45268
rect 43898 45228 43904 45240
rect 43956 45228 43962 45280
rect 46937 45271 46995 45277
rect 46937 45237 46949 45271
rect 46983 45268 46995 45271
rect 47302 45268 47308 45280
rect 46983 45240 47308 45268
rect 46983 45237 46995 45240
rect 46937 45231 46995 45237
rect 47302 45228 47308 45240
rect 47360 45228 47366 45280
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 2222 45064 2228 45076
rect 2183 45036 2228 45064
rect 2222 45024 2228 45036
rect 2280 45024 2286 45076
rect 43809 45067 43867 45073
rect 43809 45033 43821 45067
rect 43855 45064 43867 45067
rect 44450 45064 44456 45076
rect 43855 45036 44456 45064
rect 43855 45033 43867 45036
rect 43809 45027 43867 45033
rect 44450 45024 44456 45036
rect 44508 45024 44514 45076
rect 45094 45064 45100 45076
rect 45055 45036 45100 45064
rect 45094 45024 45100 45036
rect 45152 45024 45158 45076
rect 45741 45067 45799 45073
rect 45741 45033 45753 45067
rect 45787 45064 45799 45067
rect 46474 45064 46480 45076
rect 45787 45036 46480 45064
rect 45787 45033 45799 45036
rect 45741 45027 45799 45033
rect 46474 45024 46480 45036
rect 46532 45024 46538 45076
rect 43070 44956 43076 45008
rect 43128 44996 43134 45008
rect 47486 44996 47492 45008
rect 43128 44968 47492 44996
rect 43128 44956 43134 44968
rect 47486 44956 47492 44968
rect 47544 44956 47550 45008
rect 44453 44931 44511 44937
rect 44453 44897 44465 44931
rect 44499 44928 44511 44931
rect 45186 44928 45192 44940
rect 44499 44900 45192 44928
rect 44499 44897 44511 44900
rect 44453 44891 44511 44897
rect 45186 44888 45192 44900
rect 45244 44888 45250 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 2038 44820 2044 44872
rect 2096 44860 2102 44872
rect 2133 44863 2191 44869
rect 2133 44860 2145 44863
rect 2096 44832 2145 44860
rect 2096 44820 2102 44832
rect 2133 44829 2145 44832
rect 2179 44829 2191 44863
rect 45002 44860 45008 44872
rect 44963 44832 45008 44860
rect 2133 44823 2191 44829
rect 45002 44820 45008 44832
rect 45060 44820 45066 44872
rect 45646 44860 45652 44872
rect 45559 44832 45652 44860
rect 45646 44820 45652 44832
rect 45704 44820 45710 44872
rect 46290 44860 46296 44872
rect 46251 44832 46296 44860
rect 46290 44820 46296 44832
rect 46348 44820 46354 44872
rect 45664 44792 45692 44820
rect 46477 44795 46535 44801
rect 45664 44764 45784 44792
rect 45756 44724 45784 44764
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 47670 44792 47676 44804
rect 46523 44764 47676 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 47670 44752 47676 44764
rect 47728 44752 47734 44804
rect 46658 44724 46664 44736
rect 45756 44696 46664 44724
rect 46658 44684 46664 44696
rect 46716 44684 46722 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 45370 44480 45376 44532
rect 45428 44520 45434 44532
rect 46293 44523 46351 44529
rect 46293 44520 46305 44523
rect 45428 44492 46305 44520
rect 45428 44480 45434 44492
rect 46293 44489 46305 44492
rect 46339 44489 46351 44523
rect 47670 44520 47676 44532
rect 47631 44492 47676 44520
rect 46293 44483 46351 44489
rect 47670 44480 47676 44492
rect 47728 44480 47734 44532
rect 41322 44412 41328 44464
rect 41380 44452 41386 44464
rect 45554 44452 45560 44464
rect 41380 44424 45560 44452
rect 41380 44412 41386 44424
rect 45554 44412 45560 44424
rect 45612 44452 45618 44464
rect 45612 44424 46888 44452
rect 45612 44412 45618 44424
rect 45738 44384 45744 44396
rect 45699 44356 45744 44384
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46198 44384 46204 44396
rect 46159 44356 46204 44384
rect 46198 44344 46204 44356
rect 46256 44344 46262 44396
rect 46860 44393 46888 44424
rect 46845 44387 46903 44393
rect 46845 44353 46857 44387
rect 46891 44384 46903 44387
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 46891 44356 47593 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 31754 44276 31760 44328
rect 31812 44316 31818 44328
rect 38565 44319 38623 44325
rect 38565 44316 38577 44319
rect 31812 44288 38577 44316
rect 31812 44276 31818 44288
rect 38565 44285 38577 44288
rect 38611 44285 38623 44319
rect 38746 44316 38752 44328
rect 38707 44288 38752 44316
rect 38565 44279 38623 44285
rect 38746 44276 38752 44288
rect 38804 44276 38810 44328
rect 40034 44316 40040 44328
rect 39995 44288 40040 44316
rect 40034 44276 40040 44288
rect 40092 44276 40098 44328
rect 45097 44183 45155 44189
rect 45097 44149 45109 44183
rect 45143 44180 45155 44183
rect 45922 44180 45928 44192
rect 45143 44152 45928 44180
rect 45143 44149 45155 44152
rect 45097 44143 45155 44149
rect 45922 44140 45928 44152
rect 45980 44140 45986 44192
rect 46934 44180 46940 44192
rect 46895 44152 46940 44180
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 28169 43979 28227 43985
rect 28169 43945 28181 43979
rect 28215 43976 28227 43979
rect 31754 43976 31760 43988
rect 28215 43948 31760 43976
rect 28215 43945 28227 43948
rect 28169 43939 28227 43945
rect 31754 43936 31760 43948
rect 31812 43936 31818 43988
rect 38746 43976 38752 43988
rect 38707 43948 38752 43976
rect 38746 43936 38752 43948
rect 38804 43936 38810 43988
rect 45833 43979 45891 43985
rect 45833 43945 45845 43979
rect 45879 43976 45891 43979
rect 46290 43976 46296 43988
rect 45879 43948 46296 43976
rect 45879 43945 45891 43948
rect 45833 43939 45891 43945
rect 46290 43936 46296 43948
rect 46348 43936 46354 43988
rect 45922 43800 45928 43852
rect 45980 43840 45986 43852
rect 46293 43843 46351 43849
rect 46293 43840 46305 43843
rect 45980 43812 46305 43840
rect 45980 43800 45986 43812
rect 46293 43809 46305 43812
rect 46339 43809 46351 43843
rect 46293 43803 46351 43809
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 46934 43840 46940 43852
rect 46523 43812 46940 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 46934 43800 46940 43812
rect 46992 43800 46998 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 25774 43732 25780 43784
rect 25832 43772 25838 43784
rect 28077 43775 28135 43781
rect 28077 43772 28089 43775
rect 25832 43744 28089 43772
rect 25832 43732 25838 43744
rect 28077 43741 28089 43744
rect 28123 43741 28135 43775
rect 38654 43772 38660 43784
rect 38615 43744 38660 43772
rect 28077 43735 28135 43741
rect 38654 43732 38660 43744
rect 38712 43732 38718 43784
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 45462 43256 45468 43308
rect 45520 43296 45526 43308
rect 46845 43299 46903 43305
rect 46845 43296 46857 43299
rect 45520 43268 46857 43296
rect 45520 43256 45526 43268
rect 46845 43265 46857 43268
rect 46891 43265 46903 43299
rect 46845 43259 46903 43265
rect 1673 43231 1731 43237
rect 1673 43197 1685 43231
rect 1719 43228 1731 43231
rect 35710 43228 35716 43240
rect 1719 43200 35716 43228
rect 1719 43197 1731 43200
rect 1673 43191 1731 43197
rect 35710 43188 35716 43200
rect 35768 43188 35774 43240
rect 46934 43052 46940 43104
rect 46992 43092 46998 43104
rect 47765 43095 47823 43101
rect 47765 43092 47777 43095
rect 46992 43064 47777 43092
rect 46992 43052 46998 43064
rect 47765 43061 47777 43064
rect 47811 43061 47823 43095
rect 47765 43055 47823 43061
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46293 42755 46351 42761
rect 46293 42721 46305 42755
rect 46339 42752 46351 42755
rect 46934 42752 46940 42764
rect 46339 42724 46940 42752
rect 46339 42721 46351 42724
rect 46293 42715 46351 42721
rect 46934 42712 46940 42724
rect 46992 42712 46998 42764
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 47486 42168 47492 42220
rect 47544 42208 47550 42220
rect 47581 42211 47639 42217
rect 47581 42208 47593 42211
rect 47544 42180 47593 42208
rect 47544 42168 47550 42180
rect 47581 42177 47593 42180
rect 47627 42177 47639 42211
rect 47581 42171 47639 42177
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46477 41531 46535 41537
rect 46477 41497 46489 41531
rect 46523 41528 46535 41531
rect 46934 41528 46940 41540
rect 46523 41500 46940 41528
rect 46523 41497 46535 41500
rect 46477 41491 46535 41497
rect 46934 41488 46940 41500
rect 46992 41488 46998 41540
rect 48130 41528 48136 41540
rect 48091 41500 48136 41528
rect 48130 41488 48136 41500
rect 48188 41488 48194 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 46934 41256 46940 41268
rect 46895 41228 46940 41256
rect 2133 41219 2191 41225
rect 46934 41216 46940 41228
rect 46992 41216 46998 41268
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 46658 41080 46664 41132
rect 46716 41120 46722 41132
rect 46845 41123 46903 41129
rect 46845 41120 46857 41123
rect 46716 41092 46857 41120
rect 46716 41080 46722 41092
rect 46845 41089 46857 41092
rect 46891 41089 46903 41123
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 46845 41083 46903 41089
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 48133 40987 48191 40993
rect 48133 40984 48145 40987
rect 45526 40956 48145 40984
rect 38930 40876 38936 40928
rect 38988 40916 38994 40928
rect 45526 40916 45554 40956
rect 48133 40953 48145 40956
rect 48179 40953 48191 40987
rect 48133 40947 48191 40953
rect 38988 40888 45554 40916
rect 38988 40876 38994 40888
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 1946 40372 1952 40384
rect 1907 40344 1952 40372
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 23566 39448 23572 39500
rect 23624 39488 23630 39500
rect 24949 39491 25007 39497
rect 24949 39488 24961 39491
rect 23624 39460 24961 39488
rect 23624 39448 23630 39460
rect 24949 39457 24961 39460
rect 24995 39457 25007 39491
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 24949 39451 25007 39457
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 23385 39423 23443 39429
rect 23385 39389 23397 39423
rect 23431 39420 23443 39423
rect 24762 39420 24768 39432
rect 23431 39392 24440 39420
rect 24723 39392 24768 39420
rect 23431 39389 23443 39392
rect 23385 39383 23443 39389
rect 22738 39244 22744 39296
rect 22796 39284 22802 39296
rect 24412 39293 24440 39392
rect 24762 39380 24768 39392
rect 24820 39380 24826 39432
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 46842 39352 46848 39364
rect 46523 39324 46848 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 46842 39312 46848 39324
rect 46900 39312 46906 39364
rect 23201 39287 23259 39293
rect 23201 39284 23213 39287
rect 22796 39256 23213 39284
rect 22796 39244 22802 39256
rect 23201 39253 23213 39256
rect 23247 39253 23259 39287
rect 23201 39247 23259 39253
rect 24397 39287 24455 39293
rect 24397 39253 24409 39287
rect 24443 39253 24455 39287
rect 24397 39247 24455 39253
rect 24486 39244 24492 39296
rect 24544 39284 24550 39296
rect 24857 39287 24915 39293
rect 24857 39284 24869 39287
rect 24544 39256 24869 39284
rect 24544 39244 24550 39256
rect 24857 39253 24869 39256
rect 24903 39253 24915 39287
rect 24857 39247 24915 39253
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 23566 39080 23572 39092
rect 22066 39052 23572 39080
rect 20257 39015 20315 39021
rect 20257 38981 20269 39015
rect 20303 39012 20315 39015
rect 21818 39012 21824 39024
rect 20303 38984 21824 39012
rect 20303 38981 20315 38984
rect 20257 38975 20315 38981
rect 21818 38972 21824 38984
rect 21876 38972 21882 39024
rect 20441 38947 20499 38953
rect 20441 38913 20453 38947
rect 20487 38944 20499 38947
rect 22066 38944 22094 39052
rect 23566 39040 23572 39052
rect 23624 39040 23630 39092
rect 46842 39080 46848 39092
rect 46803 39052 46848 39080
rect 46842 39040 46848 39052
rect 46900 39040 46906 39092
rect 22738 39012 22744 39024
rect 22699 38984 22744 39012
rect 22738 38972 22744 38984
rect 22796 38972 22802 39024
rect 23474 38972 23480 39024
rect 23532 38972 23538 39024
rect 44266 38944 44272 38956
rect 20487 38916 22094 38944
rect 44227 38916 44272 38944
rect 20487 38913 20499 38916
rect 20441 38907 20499 38913
rect 44266 38904 44272 38916
rect 44324 38904 44330 38956
rect 45830 38904 45836 38956
rect 45888 38944 45894 38956
rect 46753 38947 46811 38953
rect 46753 38944 46765 38947
rect 45888 38916 46765 38944
rect 45888 38904 45894 38916
rect 46753 38913 46765 38916
rect 46799 38913 46811 38947
rect 47854 38944 47860 38956
rect 47815 38916 47860 38944
rect 46753 38907 46811 38913
rect 47854 38904 47860 38916
rect 47912 38904 47918 38956
rect 21910 38836 21916 38888
rect 21968 38876 21974 38888
rect 22465 38879 22523 38885
rect 22465 38876 22477 38879
rect 21968 38848 22477 38876
rect 21968 38836 21974 38848
rect 22465 38845 22477 38848
rect 22511 38845 22523 38879
rect 22465 38839 22523 38845
rect 44726 38836 44732 38888
rect 44784 38876 44790 38888
rect 45005 38879 45063 38885
rect 45005 38876 45017 38879
rect 44784 38848 45017 38876
rect 44784 38836 44790 38848
rect 45005 38845 45017 38848
rect 45051 38876 45063 38879
rect 46658 38876 46664 38888
rect 45051 38848 46664 38876
rect 45051 38845 45063 38848
rect 45005 38839 45063 38845
rect 46658 38836 46664 38848
rect 46716 38836 46722 38888
rect 48041 38811 48099 38817
rect 48041 38808 48053 38811
rect 45526 38780 48053 38808
rect 20530 38700 20536 38752
rect 20588 38740 20594 38752
rect 20625 38743 20683 38749
rect 20625 38740 20637 38743
rect 20588 38712 20637 38740
rect 20588 38700 20594 38712
rect 20625 38709 20637 38712
rect 20671 38709 20683 38743
rect 24210 38740 24216 38752
rect 24171 38712 24216 38740
rect 20625 38703 20683 38709
rect 24210 38700 24216 38712
rect 24268 38700 24274 38752
rect 44174 38700 44180 38752
rect 44232 38740 44238 38752
rect 45526 38740 45554 38780
rect 48041 38777 48053 38780
rect 48087 38777 48099 38811
rect 48041 38771 48099 38777
rect 44232 38712 45554 38740
rect 44232 38700 44238 38712
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 22741 38539 22799 38545
rect 22741 38505 22753 38539
rect 22787 38536 22799 38539
rect 23474 38536 23480 38548
rect 22787 38508 23480 38536
rect 22787 38505 22799 38508
rect 22741 38499 22799 38505
rect 23474 38496 23480 38508
rect 23532 38496 23538 38548
rect 38654 38496 38660 38548
rect 38712 38536 38718 38548
rect 46750 38536 46756 38548
rect 38712 38508 46756 38536
rect 38712 38496 38718 38508
rect 46750 38496 46756 38508
rect 46808 38496 46814 38548
rect 20533 38471 20591 38477
rect 20533 38437 20545 38471
rect 20579 38468 20591 38471
rect 21082 38468 21088 38480
rect 20579 38440 21088 38468
rect 20579 38437 20591 38440
rect 20533 38431 20591 38437
rect 21082 38428 21088 38440
rect 21140 38468 21146 38480
rect 23845 38471 23903 38477
rect 21140 38440 22094 38468
rect 21140 38428 21146 38440
rect 15838 38292 15844 38344
rect 15896 38332 15902 38344
rect 17129 38335 17187 38341
rect 17129 38332 17141 38335
rect 15896 38304 17141 38332
rect 15896 38292 15902 38304
rect 17129 38301 17141 38304
rect 17175 38301 17187 38335
rect 17129 38295 17187 38301
rect 17218 38292 17224 38344
rect 17276 38332 17282 38344
rect 17313 38335 17371 38341
rect 17313 38332 17325 38335
rect 17276 38304 17325 38332
rect 17276 38292 17282 38304
rect 17313 38301 17325 38304
rect 17359 38301 17371 38335
rect 20346 38332 20352 38344
rect 20259 38304 20352 38332
rect 17313 38295 17371 38301
rect 20346 38292 20352 38304
rect 20404 38332 20410 38344
rect 20622 38332 20628 38344
rect 20404 38304 20628 38332
rect 20404 38292 20410 38304
rect 20622 38292 20628 38304
rect 20680 38292 20686 38344
rect 22066 38332 22094 38440
rect 23845 38437 23857 38471
rect 23891 38468 23903 38471
rect 24486 38468 24492 38480
rect 23891 38440 24492 38468
rect 23891 38437 23903 38440
rect 23845 38431 23903 38437
rect 24486 38428 24492 38440
rect 24544 38428 24550 38480
rect 23385 38403 23443 38409
rect 23385 38369 23397 38403
rect 23431 38400 23443 38403
rect 23658 38400 23664 38412
rect 23431 38372 23664 38400
rect 23431 38369 23443 38372
rect 23385 38363 23443 38369
rect 23658 38360 23664 38372
rect 23716 38360 23722 38412
rect 42978 38400 42984 38412
rect 42939 38372 42984 38400
rect 42978 38360 42984 38372
rect 43036 38360 43042 38412
rect 44361 38403 44419 38409
rect 44361 38369 44373 38403
rect 44407 38400 44419 38403
rect 45002 38400 45008 38412
rect 44407 38372 45008 38400
rect 44407 38369 44419 38372
rect 44361 38363 44419 38369
rect 45002 38360 45008 38372
rect 45060 38360 45066 38412
rect 45465 38403 45523 38409
rect 45465 38369 45477 38403
rect 45511 38369 45523 38403
rect 45465 38363 45523 38369
rect 22649 38335 22707 38341
rect 22649 38332 22661 38335
rect 22066 38304 22661 38332
rect 22649 38301 22661 38304
rect 22695 38301 22707 38335
rect 22649 38295 22707 38301
rect 23477 38335 23535 38341
rect 23477 38301 23489 38335
rect 23523 38332 23535 38335
rect 23566 38332 23572 38344
rect 23523 38304 23572 38332
rect 23523 38301 23535 38304
rect 23477 38295 23535 38301
rect 23566 38292 23572 38304
rect 23624 38332 23630 38344
rect 24210 38332 24216 38344
rect 23624 38304 24216 38332
rect 23624 38292 23630 38304
rect 24210 38292 24216 38304
rect 24268 38292 24274 38344
rect 42613 38335 42671 38341
rect 42613 38301 42625 38335
rect 42659 38332 42671 38335
rect 43809 38335 43867 38341
rect 43809 38332 43821 38335
rect 42659 38304 43821 38332
rect 42659 38301 42671 38304
rect 42613 38295 42671 38301
rect 43809 38301 43821 38304
rect 43855 38332 43867 38335
rect 44266 38332 44272 38344
rect 43855 38304 44272 38332
rect 43855 38301 43867 38304
rect 43809 38295 43867 38301
rect 44266 38292 44272 38304
rect 44324 38332 44330 38344
rect 45097 38335 45155 38341
rect 45097 38332 45109 38335
rect 44324 38304 45109 38332
rect 44324 38292 44330 38304
rect 45097 38301 45109 38304
rect 45143 38301 45155 38335
rect 45097 38295 45155 38301
rect 45480 38276 45508 38363
rect 46290 38332 46296 38344
rect 46251 38304 46296 38332
rect 46290 38292 46296 38304
rect 46348 38292 46354 38344
rect 45462 38224 45468 38276
rect 45520 38264 45526 38276
rect 45554 38264 45560 38276
rect 45520 38236 45560 38264
rect 45520 38224 45526 38236
rect 45554 38224 45560 38236
rect 45612 38224 45618 38276
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 46842 38264 46848 38276
rect 46523 38236 46848 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 46842 38224 46848 38236
rect 46900 38224 46906 38276
rect 48130 38264 48136 38276
rect 48091 38236 48136 38264
rect 48130 38224 48136 38236
rect 48188 38224 48194 38276
rect 17221 38199 17279 38205
rect 17221 38165 17233 38199
rect 17267 38196 17279 38199
rect 19242 38196 19248 38208
rect 17267 38168 19248 38196
rect 17267 38165 17279 38168
rect 17221 38159 17279 38165
rect 19242 38156 19248 38168
rect 19300 38156 19306 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 26421 37995 26479 38001
rect 26421 37992 26433 37995
rect 24412 37964 26433 37992
rect 21913 37927 21971 37933
rect 21913 37924 21925 37927
rect 21022 37896 21925 37924
rect 21913 37893 21925 37896
rect 21959 37893 21971 37927
rect 21913 37887 21971 37893
rect 23293 37927 23351 37933
rect 23293 37893 23305 37927
rect 23339 37924 23351 37927
rect 23842 37924 23848 37936
rect 23339 37896 23848 37924
rect 23339 37893 23351 37896
rect 23293 37887 23351 37893
rect 23842 37884 23848 37896
rect 23900 37884 23906 37936
rect 21818 37856 21824 37868
rect 21779 37828 21824 37856
rect 21818 37816 21824 37828
rect 21876 37816 21882 37868
rect 23566 37856 23572 37868
rect 23527 37828 23572 37856
rect 23566 37816 23572 37828
rect 23624 37816 23630 37868
rect 19518 37788 19524 37800
rect 19479 37760 19524 37788
rect 19518 37748 19524 37760
rect 19576 37748 19582 37800
rect 19794 37788 19800 37800
rect 19755 37760 19800 37788
rect 19794 37748 19800 37760
rect 19852 37748 19858 37800
rect 23477 37791 23535 37797
rect 23477 37757 23489 37791
rect 23523 37788 23535 37791
rect 23750 37788 23756 37800
rect 23523 37760 23756 37788
rect 23523 37757 23535 37760
rect 23477 37751 23535 37757
rect 23750 37748 23756 37760
rect 23808 37788 23814 37800
rect 24412 37788 24440 37964
rect 26421 37961 26433 37964
rect 26467 37961 26479 37995
rect 46842 37992 46848 38004
rect 46803 37964 46848 37992
rect 26421 37955 26479 37961
rect 46842 37952 46848 37964
rect 46900 37952 46906 38004
rect 25958 37884 25964 37936
rect 26016 37884 26022 37936
rect 46290 37884 46296 37936
rect 46348 37924 46354 37936
rect 46348 37896 47808 37924
rect 46348 37884 46354 37896
rect 27798 37856 27804 37868
rect 27759 37828 27804 37856
rect 27798 37816 27804 37828
rect 27856 37816 27862 37868
rect 44266 37856 44272 37868
rect 44227 37828 44272 37856
rect 44266 37816 44272 37828
rect 44324 37816 44330 37868
rect 46750 37856 46756 37868
rect 46711 37828 46756 37856
rect 46750 37816 46756 37828
rect 46808 37816 46814 37868
rect 47780 37865 47808 37896
rect 47765 37859 47823 37865
rect 47765 37825 47777 37859
rect 47811 37825 47823 37859
rect 47765 37819 47823 37825
rect 23808 37760 24440 37788
rect 24673 37791 24731 37797
rect 23808 37748 23814 37760
rect 24673 37757 24685 37791
rect 24719 37757 24731 37791
rect 24946 37788 24952 37800
rect 24907 37760 24952 37788
rect 24673 37751 24731 37757
rect 21269 37723 21327 37729
rect 21269 37689 21281 37723
rect 21315 37720 21327 37723
rect 22094 37720 22100 37732
rect 21315 37692 22100 37720
rect 21315 37689 21327 37692
rect 21269 37683 21327 37689
rect 22094 37680 22100 37692
rect 22152 37720 22158 37732
rect 22152 37692 23336 37720
rect 22152 37680 22158 37692
rect 23308 37661 23336 37692
rect 23293 37655 23351 37661
rect 23293 37621 23305 37655
rect 23339 37621 23351 37655
rect 23293 37615 23351 37621
rect 23382 37612 23388 37664
rect 23440 37652 23446 37664
rect 23753 37655 23811 37661
rect 23753 37652 23765 37655
rect 23440 37624 23765 37652
rect 23440 37612 23446 37624
rect 23753 37621 23765 37624
rect 23799 37621 23811 37655
rect 24688 37652 24716 37751
rect 24946 37748 24952 37760
rect 25004 37748 25010 37800
rect 45097 37791 45155 37797
rect 45097 37757 45109 37791
rect 45143 37788 45155 37791
rect 45554 37788 45560 37800
rect 45143 37760 45560 37788
rect 45143 37757 45155 37760
rect 45097 37751 45155 37757
rect 45554 37748 45560 37760
rect 45612 37788 45618 37800
rect 46198 37788 46204 37800
rect 45612 37760 46204 37788
rect 45612 37748 45618 37760
rect 46198 37748 46204 37760
rect 46256 37748 46262 37800
rect 26326 37652 26332 37664
rect 24688 37624 26332 37652
rect 23753 37615 23811 37621
rect 26326 37612 26332 37624
rect 26384 37612 26390 37664
rect 27893 37655 27951 37661
rect 27893 37621 27905 37655
rect 27939 37652 27951 37655
rect 27982 37652 27988 37664
rect 27939 37624 27988 37652
rect 27939 37621 27951 37624
rect 27893 37615 27951 37621
rect 27982 37612 27988 37624
rect 28040 37612 28046 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 19794 37408 19800 37460
rect 19852 37448 19858 37460
rect 20441 37451 20499 37457
rect 20441 37448 20453 37451
rect 19852 37420 20453 37448
rect 19852 37408 19858 37420
rect 20441 37417 20453 37420
rect 20487 37417 20499 37451
rect 20441 37411 20499 37417
rect 21085 37451 21143 37457
rect 21085 37417 21097 37451
rect 21131 37448 21143 37451
rect 21818 37448 21824 37460
rect 21131 37420 21824 37448
rect 21131 37417 21143 37420
rect 21085 37411 21143 37417
rect 21818 37408 21824 37420
rect 21876 37408 21882 37460
rect 24946 37408 24952 37460
rect 25004 37448 25010 37460
rect 25133 37451 25191 37457
rect 25133 37448 25145 37451
rect 25004 37420 25145 37448
rect 25004 37408 25010 37420
rect 25133 37417 25145 37420
rect 25179 37417 25191 37451
rect 44266 37448 44272 37460
rect 44227 37420 44272 37448
rect 25133 37411 25191 37417
rect 44266 37408 44272 37420
rect 44324 37408 44330 37460
rect 19904 37284 20208 37312
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 2041 37207 2099 37213
rect 19242 37204 19248 37256
rect 19300 37244 19306 37256
rect 19904 37244 19932 37284
rect 20070 37244 20076 37256
rect 19300 37216 19932 37244
rect 20031 37216 20076 37244
rect 19300 37204 19306 37216
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 20180 37244 20208 37284
rect 20254 37272 20260 37324
rect 20312 37312 20318 37324
rect 21836 37312 21864 37408
rect 42978 37340 42984 37392
rect 43036 37380 43042 37392
rect 47026 37380 47032 37392
rect 43036 37352 47032 37380
rect 43036 37340 43042 37352
rect 47026 37340 47032 37352
rect 47084 37340 47090 37392
rect 20312 37284 20357 37312
rect 21836 37284 23428 37312
rect 20312 37272 20318 37284
rect 20441 37247 20499 37253
rect 20441 37244 20453 37247
rect 20180 37216 20453 37244
rect 20441 37213 20453 37216
rect 20487 37213 20499 37247
rect 20441 37207 20499 37213
rect 20622 37204 20628 37256
rect 20680 37244 20686 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20680 37216 20913 37244
rect 20680 37204 20686 37216
rect 20901 37213 20913 37216
rect 20947 37213 20959 37247
rect 21910 37244 21916 37256
rect 21871 37216 21916 37244
rect 20901 37207 20959 37213
rect 21910 37204 21916 37216
rect 21968 37204 21974 37256
rect 23400 37244 23428 37284
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 23400 37216 24409 37244
rect 24397 37213 24409 37216
rect 24443 37244 24455 37247
rect 24443 37216 25084 37244
rect 24443 37213 24455 37216
rect 24397 37207 24455 37213
rect 17310 37136 17316 37188
rect 17368 37176 17374 37188
rect 19518 37176 19524 37188
rect 17368 37148 19524 37176
rect 17368 37136 17374 37148
rect 19518 37136 19524 37148
rect 19576 37176 19582 37188
rect 19978 37176 19984 37188
rect 19576 37148 19984 37176
rect 19576 37136 19582 37148
rect 19978 37136 19984 37148
rect 20036 37176 20042 37188
rect 21928 37176 21956 37204
rect 22186 37176 22192 37188
rect 20036 37148 21956 37176
rect 22147 37148 22192 37176
rect 20036 37136 20042 37148
rect 22186 37136 22192 37148
rect 22244 37136 22250 37188
rect 24489 37179 24547 37185
rect 24489 37176 24501 37179
rect 23414 37148 24501 37176
rect 24489 37145 24501 37148
rect 24535 37145 24547 37179
rect 25056 37176 25084 37216
rect 25130 37204 25136 37256
rect 25188 37244 25194 37256
rect 25317 37247 25375 37253
rect 25317 37244 25329 37247
rect 25188 37216 25329 37244
rect 25188 37204 25194 37216
rect 25317 37213 25329 37216
rect 25363 37213 25375 37247
rect 25317 37207 25375 37213
rect 25869 37247 25927 37253
rect 25869 37213 25881 37247
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 25884 37176 25912 37207
rect 25958 37204 25964 37256
rect 26016 37244 26022 37256
rect 26016 37216 26061 37244
rect 26016 37204 26022 37216
rect 26326 37204 26332 37256
rect 26384 37244 26390 37256
rect 26697 37247 26755 37253
rect 26697 37244 26709 37247
rect 26384 37216 26709 37244
rect 26384 37204 26390 37216
rect 26697 37213 26709 37216
rect 26743 37213 26755 37247
rect 26697 37207 26755 37213
rect 43622 37204 43628 37256
rect 43680 37244 43686 37256
rect 44174 37244 44180 37256
rect 43680 37216 44180 37244
rect 43680 37204 43686 37216
rect 44174 37204 44180 37216
rect 44232 37204 44238 37256
rect 26970 37176 26976 37188
rect 25056 37148 25912 37176
rect 26931 37148 26976 37176
rect 24489 37139 24547 37145
rect 20165 37111 20223 37117
rect 20165 37077 20177 37111
rect 20211 37108 20223 37111
rect 23566 37108 23572 37120
rect 20211 37080 23572 37108
rect 20211 37077 20223 37080
rect 20165 37071 20223 37077
rect 23566 37068 23572 37080
rect 23624 37068 23630 37120
rect 23661 37111 23719 37117
rect 23661 37077 23673 37111
rect 23707 37108 23719 37111
rect 23842 37108 23848 37120
rect 23707 37080 23848 37108
rect 23707 37077 23719 37080
rect 23661 37071 23719 37077
rect 23842 37068 23848 37080
rect 23900 37068 23906 37120
rect 25884 37108 25912 37148
rect 26970 37136 26976 37148
rect 27028 37136 27034 37188
rect 27982 37136 27988 37188
rect 28040 37136 28046 37188
rect 27798 37108 27804 37120
rect 25884 37080 27804 37108
rect 27798 37068 27804 37080
rect 27856 37068 27862 37120
rect 28442 37108 28448 37120
rect 28403 37080 28448 37108
rect 28442 37068 28448 37080
rect 28500 37068 28506 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 9490 36864 9496 36916
rect 9548 36904 9554 36916
rect 9548 36876 18920 36904
rect 9548 36864 9554 36876
rect 18322 36796 18328 36848
rect 18380 36796 18386 36848
rect 18892 36836 18920 36876
rect 20070 36864 20076 36916
rect 20128 36904 20134 36916
rect 22097 36907 22155 36913
rect 22097 36904 22109 36907
rect 20128 36876 22109 36904
rect 20128 36864 20134 36876
rect 22097 36873 22109 36876
rect 22143 36873 22155 36907
rect 22097 36867 22155 36873
rect 23477 36907 23535 36913
rect 23477 36873 23489 36907
rect 23523 36904 23535 36907
rect 23658 36904 23664 36916
rect 23523 36876 23664 36904
rect 23523 36873 23535 36876
rect 23477 36867 23535 36873
rect 23658 36864 23664 36876
rect 23716 36864 23722 36916
rect 25774 36904 25780 36916
rect 25735 36876 25780 36904
rect 25774 36864 25780 36876
rect 25832 36864 25838 36916
rect 26970 36904 26976 36916
rect 26931 36876 26976 36904
rect 26970 36864 26976 36876
rect 27028 36864 27034 36916
rect 27798 36864 27804 36916
rect 27856 36904 27862 36916
rect 27856 36876 28488 36904
rect 27856 36864 27862 36876
rect 28353 36839 28411 36845
rect 28353 36836 28365 36839
rect 18892 36808 24808 36836
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 15749 36771 15807 36777
rect 15749 36737 15761 36771
rect 15795 36768 15807 36771
rect 16022 36768 16028 36780
rect 15795 36740 16028 36768
rect 15795 36737 15807 36740
rect 15749 36731 15807 36737
rect 16022 36728 16028 36740
rect 16080 36728 16086 36780
rect 17310 36768 17316 36780
rect 17271 36740 17316 36768
rect 17310 36728 17316 36740
rect 17368 36728 17374 36780
rect 20438 36728 20444 36780
rect 20496 36768 20502 36780
rect 20622 36768 20628 36780
rect 20496 36740 20628 36768
rect 20496 36728 20502 36740
rect 20622 36728 20628 36740
rect 20680 36728 20686 36780
rect 21818 36768 21824 36780
rect 21779 36740 21824 36768
rect 21818 36728 21824 36740
rect 21876 36728 21882 36780
rect 23293 36771 23351 36777
rect 23293 36737 23305 36771
rect 23339 36768 23351 36771
rect 23474 36768 23480 36780
rect 23339 36740 23480 36768
rect 23339 36737 23351 36740
rect 23293 36731 23351 36737
rect 23474 36728 23480 36740
rect 23532 36728 23538 36780
rect 23661 36771 23719 36777
rect 23661 36737 23673 36771
rect 23707 36737 23719 36771
rect 23661 36731 23719 36737
rect 23845 36771 23903 36777
rect 23845 36737 23857 36771
rect 23891 36737 23903 36771
rect 23845 36731 23903 36737
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 17589 36703 17647 36709
rect 17589 36669 17601 36703
rect 17635 36700 17647 36703
rect 18230 36700 18236 36712
rect 17635 36672 18236 36700
rect 17635 36669 17647 36672
rect 17589 36663 17647 36669
rect 18230 36660 18236 36672
rect 18288 36660 18294 36712
rect 22094 36660 22100 36712
rect 22152 36700 22158 36712
rect 23676 36700 23704 36731
rect 22152 36672 23704 36700
rect 22152 36660 22158 36672
rect 21913 36635 21971 36641
rect 21913 36601 21925 36635
rect 21959 36632 21971 36635
rect 23198 36632 23204 36644
rect 21959 36604 23204 36632
rect 21959 36601 21971 36604
rect 21913 36595 21971 36601
rect 23198 36592 23204 36604
rect 23256 36632 23262 36644
rect 23860 36632 23888 36731
rect 24780 36700 24808 36808
rect 27172 36808 28365 36836
rect 25222 36728 25228 36780
rect 25280 36768 25286 36780
rect 27172 36777 27200 36808
rect 28353 36805 28365 36808
rect 28399 36805 28411 36839
rect 28353 36799 28411 36805
rect 25593 36771 25651 36777
rect 25593 36768 25605 36771
rect 25280 36740 25605 36768
rect 25280 36728 25286 36740
rect 25593 36737 25605 36740
rect 25639 36737 25651 36771
rect 25593 36731 25651 36737
rect 27157 36771 27215 36777
rect 27157 36737 27169 36771
rect 27203 36737 27215 36771
rect 27157 36731 27215 36737
rect 27246 36728 27252 36780
rect 27304 36768 27310 36780
rect 27522 36768 27528 36780
rect 27304 36740 27349 36768
rect 27483 36740 27528 36768
rect 27304 36728 27310 36740
rect 27522 36728 27528 36740
rect 27580 36728 27586 36780
rect 28169 36771 28227 36777
rect 28169 36768 28181 36771
rect 27632 36740 28181 36768
rect 27433 36703 27491 36709
rect 27433 36700 27445 36703
rect 24780 36672 27445 36700
rect 27433 36669 27445 36672
rect 27479 36669 27491 36703
rect 27632 36700 27660 36740
rect 28169 36737 28181 36740
rect 28215 36737 28227 36771
rect 28460 36768 28488 36876
rect 28997 36771 29055 36777
rect 28997 36768 29009 36771
rect 28460 36740 29009 36768
rect 28169 36731 28227 36737
rect 28997 36737 29009 36740
rect 29043 36737 29055 36771
rect 28997 36731 29055 36737
rect 27982 36700 27988 36712
rect 27433 36663 27491 36669
rect 27540 36672 27660 36700
rect 27895 36672 27988 36700
rect 27540 36644 27568 36672
rect 27982 36660 27988 36672
rect 28040 36700 28046 36712
rect 28442 36700 28448 36712
rect 28040 36672 28448 36700
rect 28040 36660 28046 36672
rect 28442 36660 28448 36672
rect 28500 36660 28506 36712
rect 23256 36604 23888 36632
rect 23256 36592 23262 36604
rect 27522 36592 27528 36644
rect 27580 36592 27586 36644
rect 15746 36524 15752 36576
rect 15804 36564 15810 36576
rect 15841 36567 15899 36573
rect 15841 36564 15853 36567
rect 15804 36536 15853 36564
rect 15804 36524 15810 36536
rect 15841 36533 15853 36536
rect 15887 36533 15899 36567
rect 19058 36564 19064 36576
rect 19019 36536 19064 36564
rect 15841 36527 15899 36533
rect 19058 36524 19064 36536
rect 19116 36524 19122 36576
rect 23753 36567 23811 36573
rect 23753 36533 23765 36567
rect 23799 36564 23811 36567
rect 24854 36564 24860 36576
rect 23799 36536 24860 36564
rect 23799 36533 23811 36536
rect 23753 36527 23811 36533
rect 24854 36524 24860 36536
rect 24912 36524 24918 36576
rect 29089 36567 29147 36573
rect 29089 36533 29101 36567
rect 29135 36564 29147 36567
rect 29362 36564 29368 36576
rect 29135 36536 29368 36564
rect 29135 36533 29147 36536
rect 29089 36527 29147 36533
rect 29362 36524 29368 36536
rect 29420 36524 29426 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 45554 36360 45560 36372
rect 6886 36332 45560 36360
rect 2133 36159 2191 36165
rect 2133 36125 2145 36159
rect 2179 36156 2191 36159
rect 2314 36156 2320 36168
rect 2179 36128 2320 36156
rect 2179 36125 2191 36128
rect 2133 36119 2191 36125
rect 2314 36116 2320 36128
rect 2372 36156 2378 36168
rect 6886 36156 6914 36332
rect 45554 36320 45560 36332
rect 45612 36320 45618 36372
rect 18230 36292 18236 36304
rect 18191 36264 18236 36292
rect 18230 36252 18236 36264
rect 18288 36252 18294 36304
rect 18616 36264 22140 36292
rect 14737 36227 14795 36233
rect 14737 36193 14749 36227
rect 14783 36224 14795 36227
rect 17310 36224 17316 36236
rect 14783 36196 17316 36224
rect 14783 36193 14795 36196
rect 14737 36187 14795 36193
rect 17310 36184 17316 36196
rect 17368 36184 17374 36236
rect 17402 36184 17408 36236
rect 17460 36224 17466 36236
rect 17460 36196 18552 36224
rect 17460 36184 17466 36196
rect 2372 36128 6914 36156
rect 18417 36159 18475 36165
rect 2372 36116 2378 36128
rect 18417 36125 18429 36159
rect 18463 36125 18475 36159
rect 18417 36119 18475 36125
rect 15013 36091 15071 36097
rect 15013 36057 15025 36091
rect 15059 36088 15071 36091
rect 15286 36088 15292 36100
rect 15059 36060 15292 36088
rect 15059 36057 15071 36060
rect 15013 36051 15071 36057
rect 15286 36048 15292 36060
rect 15344 36048 15350 36100
rect 15746 36048 15752 36100
rect 15804 36048 15810 36100
rect 16390 35980 16396 36032
rect 16448 36020 16454 36032
rect 16485 36023 16543 36029
rect 16485 36020 16497 36023
rect 16448 35992 16497 36020
rect 16448 35980 16454 35992
rect 16485 35989 16497 35992
rect 16531 35989 16543 36023
rect 18432 36020 18460 36119
rect 18524 36088 18552 36196
rect 18616 36165 18644 36264
rect 19521 36227 19579 36233
rect 19521 36193 19533 36227
rect 19567 36224 19579 36227
rect 20070 36224 20076 36236
rect 19567 36196 20076 36224
rect 19567 36193 19579 36196
rect 19521 36187 19579 36193
rect 20070 36184 20076 36196
rect 20128 36184 20134 36236
rect 22112 36224 22140 36264
rect 22186 36252 22192 36304
rect 22244 36292 22250 36304
rect 22649 36295 22707 36301
rect 22649 36292 22661 36295
rect 22244 36264 22661 36292
rect 22244 36252 22250 36264
rect 22649 36261 22661 36264
rect 22695 36261 22707 36295
rect 22649 36255 22707 36261
rect 23474 36252 23480 36304
rect 23532 36252 23538 36304
rect 24946 36292 24952 36304
rect 24907 36264 24952 36292
rect 24946 36252 24952 36264
rect 25004 36252 25010 36304
rect 25130 36292 25136 36304
rect 25091 36264 25136 36292
rect 25130 36252 25136 36264
rect 25188 36252 25194 36304
rect 22922 36224 22928 36236
rect 22112 36196 22928 36224
rect 22922 36184 22928 36196
rect 22980 36184 22986 36236
rect 23014 36184 23020 36236
rect 23072 36224 23078 36236
rect 23492 36224 23520 36252
rect 25222 36224 25228 36236
rect 23072 36196 23336 36224
rect 23492 36196 25228 36224
rect 23072 36184 23078 36196
rect 18601 36159 18659 36165
rect 18601 36125 18613 36159
rect 18647 36125 18659 36159
rect 18601 36119 18659 36125
rect 18693 36159 18751 36165
rect 18693 36125 18705 36159
rect 18739 36125 18751 36159
rect 18693 36119 18751 36125
rect 18708 36088 18736 36119
rect 19058 36116 19064 36168
rect 19116 36156 19122 36168
rect 19242 36156 19248 36168
rect 19116 36128 19248 36156
rect 19116 36116 19122 36128
rect 19242 36116 19248 36128
rect 19300 36156 19306 36168
rect 19429 36159 19487 36165
rect 19429 36156 19441 36159
rect 19300 36128 19441 36156
rect 19300 36116 19306 36128
rect 19429 36125 19441 36128
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 22554 36116 22560 36168
rect 22612 36156 22618 36168
rect 22833 36159 22891 36165
rect 22833 36156 22845 36159
rect 22612 36128 22845 36156
rect 22612 36116 22618 36128
rect 22833 36125 22845 36128
rect 22879 36125 22891 36159
rect 22833 36119 22891 36125
rect 23109 36159 23167 36165
rect 23109 36125 23121 36159
rect 23155 36156 23167 36159
rect 23308 36156 23336 36196
rect 25222 36184 25228 36196
rect 25280 36184 25286 36236
rect 23569 36159 23627 36165
rect 23569 36156 23581 36159
rect 23155 36128 23244 36156
rect 23308 36128 23581 36156
rect 23155 36125 23167 36128
rect 23109 36119 23167 36125
rect 18524 36060 18736 36088
rect 18966 36048 18972 36100
rect 19024 36088 19030 36100
rect 23216 36088 23244 36128
rect 23569 36125 23581 36128
rect 23615 36156 23627 36159
rect 23842 36156 23848 36168
rect 23615 36128 23848 36156
rect 23615 36125 23627 36128
rect 23569 36119 23627 36125
rect 23842 36116 23848 36128
rect 23900 36116 23906 36168
rect 27617 36159 27675 36165
rect 27617 36125 27629 36159
rect 27663 36156 27675 36159
rect 27982 36156 27988 36168
rect 27663 36128 27988 36156
rect 27663 36125 27675 36128
rect 27617 36119 27675 36125
rect 27982 36116 27988 36128
rect 28040 36116 28046 36168
rect 23474 36088 23480 36100
rect 19024 36060 19840 36088
rect 23216 36060 23480 36088
rect 19024 36048 19030 36060
rect 19334 36020 19340 36032
rect 18432 35992 19340 36020
rect 16485 35983 16543 35989
rect 19334 35980 19340 35992
rect 19392 35980 19398 36032
rect 19812 36029 19840 36060
rect 23474 36048 23480 36060
rect 23532 36048 23538 36100
rect 24673 36091 24731 36097
rect 24673 36057 24685 36091
rect 24719 36088 24731 36091
rect 25130 36088 25136 36100
rect 24719 36060 25136 36088
rect 24719 36057 24731 36060
rect 24673 36051 24731 36057
rect 25130 36048 25136 36060
rect 25188 36048 25194 36100
rect 27433 36091 27491 36097
rect 27433 36057 27445 36091
rect 27479 36088 27491 36091
rect 27522 36088 27528 36100
rect 27479 36060 27528 36088
rect 27479 36057 27491 36060
rect 27433 36051 27491 36057
rect 27522 36048 27528 36060
rect 27580 36048 27586 36100
rect 19797 36023 19855 36029
rect 19797 35989 19809 36023
rect 19843 35989 19855 36023
rect 23014 36020 23020 36032
rect 22975 35992 23020 36020
rect 19797 35983 19855 35989
rect 23014 35980 23020 35992
rect 23072 35980 23078 36032
rect 23661 36023 23719 36029
rect 23661 35989 23673 36023
rect 23707 36020 23719 36023
rect 24026 36020 24032 36032
rect 23707 35992 24032 36020
rect 23707 35989 23719 35992
rect 23661 35983 23719 35989
rect 24026 35980 24032 35992
rect 24084 35980 24090 36032
rect 27798 36020 27804 36032
rect 27759 35992 27804 36020
rect 27798 35980 27804 35992
rect 27856 35980 27862 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 18322 35816 18328 35828
rect 18283 35788 18328 35816
rect 18322 35776 18328 35788
rect 18380 35776 18386 35828
rect 19334 35776 19340 35828
rect 19392 35816 19398 35828
rect 19521 35819 19579 35825
rect 19521 35816 19533 35819
rect 19392 35788 19533 35816
rect 19392 35776 19398 35788
rect 19521 35785 19533 35788
rect 19567 35785 19579 35819
rect 23198 35816 23204 35828
rect 23159 35788 23204 35816
rect 19521 35779 19579 35785
rect 23198 35776 23204 35788
rect 23256 35776 23262 35828
rect 23661 35819 23719 35825
rect 23661 35785 23673 35819
rect 23707 35816 23719 35819
rect 23750 35816 23756 35828
rect 23707 35788 23756 35816
rect 23707 35785 23719 35788
rect 23661 35779 23719 35785
rect 23750 35776 23756 35788
rect 23808 35776 23814 35828
rect 24305 35819 24363 35825
rect 24305 35785 24317 35819
rect 24351 35816 24363 35819
rect 24965 35819 25023 35825
rect 24965 35816 24977 35819
rect 24351 35788 24977 35816
rect 24351 35785 24363 35788
rect 24305 35779 24363 35785
rect 24965 35785 24977 35788
rect 25011 35785 25023 35819
rect 25130 35816 25136 35828
rect 25091 35788 25136 35816
rect 24965 35779 25023 35785
rect 25130 35776 25136 35788
rect 25188 35776 25194 35828
rect 27246 35816 27252 35828
rect 27207 35788 27252 35816
rect 27246 35776 27252 35788
rect 27304 35776 27310 35828
rect 27433 35819 27491 35825
rect 27433 35785 27445 35819
rect 27479 35816 27491 35819
rect 27798 35816 27804 35828
rect 27479 35788 27804 35816
rect 27479 35785 27491 35788
rect 27433 35779 27491 35785
rect 27798 35776 27804 35788
rect 27856 35776 27862 35828
rect 16022 35708 16028 35760
rect 16080 35748 16086 35760
rect 19242 35757 19248 35760
rect 16080 35720 18276 35748
rect 16080 35708 16086 35720
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 15565 35683 15623 35689
rect 15565 35649 15577 35683
rect 15611 35680 15623 35683
rect 15611 35652 16160 35680
rect 15611 35649 15623 35652
rect 15565 35643 15623 35649
rect 16132 35624 16160 35652
rect 16574 35640 16580 35692
rect 16632 35680 16638 35692
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16632 35652 16865 35680
rect 16632 35640 16638 35652
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 16945 35683 17003 35689
rect 16945 35649 16957 35683
rect 16991 35649 17003 35683
rect 17218 35680 17224 35692
rect 17131 35652 17224 35680
rect 16945 35643 17003 35649
rect 15657 35615 15715 35621
rect 15657 35581 15669 35615
rect 15703 35612 15715 35615
rect 15746 35612 15752 35624
rect 15703 35584 15752 35612
rect 15703 35581 15715 35584
rect 15657 35575 15715 35581
rect 15746 35572 15752 35584
rect 15804 35572 15810 35624
rect 16114 35572 16120 35624
rect 16172 35612 16178 35624
rect 16390 35612 16396 35624
rect 16172 35584 16396 35612
rect 16172 35572 16178 35584
rect 16390 35572 16396 35584
rect 16448 35612 16454 35624
rect 16960 35612 16988 35643
rect 17218 35640 17224 35652
rect 17276 35640 17282 35692
rect 18248 35689 18276 35720
rect 19241 35711 19248 35757
rect 19300 35748 19306 35760
rect 19300 35720 19341 35748
rect 19242 35708 19248 35711
rect 19300 35708 19306 35720
rect 20254 35708 20260 35760
rect 20312 35748 20318 35760
rect 21910 35748 21916 35760
rect 20312 35720 21916 35748
rect 20312 35708 20318 35720
rect 21910 35708 21916 35720
rect 21968 35708 21974 35760
rect 22741 35751 22799 35757
rect 22741 35717 22753 35751
rect 22787 35748 22799 35751
rect 22787 35720 24532 35748
rect 22787 35717 22799 35720
rect 22741 35711 22799 35717
rect 18233 35683 18291 35689
rect 18233 35649 18245 35683
rect 18279 35680 18291 35683
rect 18322 35680 18328 35692
rect 18279 35652 18328 35680
rect 18279 35649 18291 35652
rect 18233 35643 18291 35649
rect 18322 35640 18328 35652
rect 18380 35640 18386 35692
rect 18966 35680 18972 35692
rect 18927 35652 18972 35680
rect 18966 35640 18972 35652
rect 19024 35640 19030 35692
rect 19153 35683 19211 35689
rect 19153 35649 19165 35683
rect 19199 35649 19211 35683
rect 19153 35643 19211 35649
rect 19337 35683 19395 35689
rect 19337 35649 19349 35683
rect 19383 35680 19395 35683
rect 21818 35680 21824 35692
rect 19383 35652 21824 35680
rect 19383 35649 19395 35652
rect 19337 35643 19395 35649
rect 17126 35612 17132 35624
rect 16448 35584 16988 35612
rect 17087 35584 17132 35612
rect 16448 35572 16454 35584
rect 17126 35572 17132 35584
rect 17184 35572 17190 35624
rect 16942 35504 16948 35556
rect 17000 35544 17006 35556
rect 17236 35544 17264 35640
rect 19168 35612 19196 35643
rect 21818 35640 21824 35652
rect 21876 35680 21882 35692
rect 22646 35680 22652 35692
rect 21876 35652 22652 35680
rect 21876 35640 21882 35652
rect 22646 35640 22652 35652
rect 22704 35640 22710 35692
rect 23017 35683 23075 35689
rect 23017 35649 23029 35683
rect 23063 35680 23075 35683
rect 23750 35680 23756 35692
rect 23063 35652 23756 35680
rect 23063 35649 23075 35652
rect 23017 35643 23075 35649
rect 23750 35640 23756 35652
rect 23808 35680 23814 35692
rect 24504 35680 24532 35720
rect 24578 35708 24584 35760
rect 24636 35748 24642 35760
rect 24765 35751 24823 35757
rect 24765 35748 24777 35751
rect 24636 35720 24777 35748
rect 24636 35708 24642 35720
rect 24765 35717 24777 35720
rect 24811 35717 24823 35751
rect 24765 35711 24823 35717
rect 26326 35708 26332 35760
rect 26384 35748 26390 35760
rect 27522 35748 27528 35760
rect 26384 35720 27528 35748
rect 26384 35708 26390 35720
rect 27522 35708 27528 35720
rect 27580 35748 27586 35760
rect 27580 35720 28672 35748
rect 27580 35708 27586 35720
rect 26237 35683 26295 35689
rect 26237 35680 26249 35683
rect 23808 35652 24472 35680
rect 24504 35652 26249 35680
rect 23808 35640 23814 35652
rect 22925 35615 22983 35621
rect 19168 35584 22876 35612
rect 20254 35544 20260 35556
rect 17000 35516 20260 35544
rect 17000 35504 17006 35516
rect 20254 35504 20260 35516
rect 20312 35504 20318 35556
rect 22848 35544 22876 35584
rect 22925 35581 22937 35615
rect 22971 35612 22983 35615
rect 23566 35612 23572 35624
rect 22971 35584 23572 35612
rect 22971 35581 22983 35584
rect 22925 35575 22983 35581
rect 23566 35572 23572 35584
rect 23624 35572 23630 35624
rect 24026 35612 24032 35624
rect 23987 35584 24032 35612
rect 24026 35572 24032 35584
rect 24084 35572 24090 35624
rect 24118 35572 24124 35624
rect 24176 35612 24182 35624
rect 24444 35612 24472 35652
rect 26237 35649 26249 35652
rect 26283 35649 26295 35683
rect 26237 35643 26295 35649
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35680 26479 35683
rect 26970 35680 26976 35692
rect 26467 35652 26976 35680
rect 26467 35649 26479 35652
rect 26421 35643 26479 35649
rect 24762 35612 24768 35624
rect 24176 35584 24221 35612
rect 24444 35584 24768 35612
rect 24176 35572 24182 35584
rect 24762 35572 24768 35584
rect 24820 35572 24826 35624
rect 26252 35612 26280 35643
rect 26970 35640 26976 35652
rect 27028 35640 27034 35692
rect 27374 35683 27432 35689
rect 27374 35680 27386 35683
rect 27080 35652 27386 35680
rect 26326 35612 26332 35624
rect 26252 35584 26332 35612
rect 26326 35572 26332 35584
rect 26384 35572 26390 35624
rect 23106 35544 23112 35556
rect 22848 35516 23112 35544
rect 23106 35504 23112 35516
rect 23164 35544 23170 35556
rect 24670 35544 24676 35556
rect 23164 35516 24676 35544
rect 23164 35504 23170 35516
rect 24670 35504 24676 35516
rect 24728 35544 24734 35556
rect 27080 35544 27108 35652
rect 27374 35649 27386 35652
rect 27420 35649 27432 35683
rect 27374 35643 27432 35649
rect 27893 35683 27951 35689
rect 27893 35649 27905 35683
rect 27939 35680 27951 35683
rect 27982 35680 27988 35692
rect 27939 35652 27988 35680
rect 27939 35649 27951 35652
rect 27893 35643 27951 35649
rect 27982 35640 27988 35652
rect 28040 35640 28046 35692
rect 28644 35689 28672 35720
rect 29362 35708 29368 35760
rect 29420 35708 29426 35760
rect 28629 35683 28687 35689
rect 28629 35649 28641 35683
rect 28675 35649 28687 35683
rect 48130 35680 48136 35692
rect 48091 35652 48136 35680
rect 28629 35643 28687 35649
rect 48130 35640 48136 35652
rect 48188 35640 48194 35692
rect 28905 35615 28963 35621
rect 28905 35581 28917 35615
rect 28951 35612 28963 35615
rect 29362 35612 29368 35624
rect 28951 35584 29368 35612
rect 28951 35581 28963 35584
rect 28905 35575 28963 35581
rect 29362 35572 29368 35584
rect 29420 35572 29426 35624
rect 24728 35516 27108 35544
rect 24728 35504 24734 35516
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 2222 35476 2228 35488
rect 1443 35448 2228 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 2222 35436 2228 35448
rect 2280 35436 2286 35488
rect 15841 35479 15899 35485
rect 15841 35445 15853 35479
rect 15887 35476 15899 35479
rect 15930 35476 15936 35488
rect 15887 35448 15936 35476
rect 15887 35445 15899 35448
rect 15841 35439 15899 35445
rect 15930 35436 15936 35448
rect 15988 35436 15994 35488
rect 16666 35476 16672 35488
rect 16627 35448 16672 35476
rect 16666 35436 16672 35448
rect 16724 35436 16730 35488
rect 23014 35476 23020 35488
rect 22975 35448 23020 35476
rect 23014 35436 23020 35448
rect 23072 35436 23078 35488
rect 23198 35436 23204 35488
rect 23256 35476 23262 35488
rect 24949 35479 25007 35485
rect 24949 35476 24961 35479
rect 23256 35448 24961 35476
rect 23256 35436 23262 35448
rect 24949 35445 24961 35448
rect 24995 35445 25007 35479
rect 26234 35476 26240 35488
rect 26195 35448 26240 35476
rect 24949 35439 25007 35445
rect 26234 35436 26240 35448
rect 26292 35436 26298 35488
rect 26418 35436 26424 35488
rect 26476 35476 26482 35488
rect 27801 35479 27859 35485
rect 27801 35476 27813 35479
rect 26476 35448 27813 35476
rect 26476 35436 26482 35448
rect 27801 35445 27813 35448
rect 27847 35476 27859 35479
rect 28350 35476 28356 35488
rect 27847 35448 28356 35476
rect 27847 35445 27859 35448
rect 27801 35439 27859 35445
rect 28350 35436 28356 35448
rect 28408 35436 28414 35488
rect 28902 35436 28908 35488
rect 28960 35476 28966 35488
rect 30377 35479 30435 35485
rect 30377 35476 30389 35479
rect 28960 35448 30389 35476
rect 28960 35436 28966 35448
rect 30377 35445 30389 35448
rect 30423 35445 30435 35479
rect 30377 35439 30435 35445
rect 47118 35436 47124 35488
rect 47176 35476 47182 35488
rect 47949 35479 48007 35485
rect 47949 35476 47961 35479
rect 47176 35448 47961 35476
rect 47176 35436 47182 35448
rect 47949 35445 47961 35448
rect 47995 35445 48007 35479
rect 47949 35439 48007 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 15286 35232 15292 35284
rect 15344 35272 15350 35284
rect 15565 35275 15623 35281
rect 15565 35272 15577 35275
rect 15344 35244 15577 35272
rect 15344 35232 15350 35244
rect 15565 35241 15577 35244
rect 15611 35241 15623 35275
rect 15930 35272 15936 35284
rect 15891 35244 15936 35272
rect 15565 35235 15623 35241
rect 15930 35232 15936 35244
rect 15988 35232 15994 35284
rect 20717 35275 20775 35281
rect 20717 35241 20729 35275
rect 20763 35272 20775 35275
rect 20806 35272 20812 35284
rect 20763 35244 20812 35272
rect 20763 35241 20775 35244
rect 20717 35235 20775 35241
rect 20806 35232 20812 35244
rect 20864 35272 20870 35284
rect 22554 35272 22560 35284
rect 20864 35244 22560 35272
rect 20864 35232 20870 35244
rect 22554 35232 22560 35244
rect 22612 35232 22618 35284
rect 22646 35232 22652 35284
rect 22704 35272 22710 35284
rect 22833 35275 22891 35281
rect 22833 35272 22845 35275
rect 22704 35244 22845 35272
rect 22704 35232 22710 35244
rect 22833 35241 22845 35244
rect 22879 35241 22891 35275
rect 22833 35235 22891 35241
rect 23474 35232 23480 35284
rect 23532 35272 23538 35284
rect 24581 35275 24639 35281
rect 24581 35272 24593 35275
rect 23532 35244 24593 35272
rect 23532 35232 23538 35244
rect 24581 35241 24593 35244
rect 24627 35241 24639 35275
rect 24581 35235 24639 35241
rect 24946 35232 24952 35284
rect 25004 35272 25010 35284
rect 25225 35275 25283 35281
rect 25225 35272 25237 35275
rect 25004 35244 25237 35272
rect 25004 35232 25010 35244
rect 25225 35241 25237 35244
rect 25271 35241 25283 35275
rect 25225 35235 25283 35241
rect 25406 35232 25412 35284
rect 25464 35272 25470 35284
rect 26418 35272 26424 35284
rect 25464 35244 26424 35272
rect 25464 35232 25470 35244
rect 26418 35232 26424 35244
rect 26476 35232 26482 35284
rect 27249 35275 27307 35281
rect 27249 35241 27261 35275
rect 27295 35272 27307 35275
rect 27982 35272 27988 35284
rect 27295 35244 27988 35272
rect 27295 35241 27307 35244
rect 27249 35235 27307 35241
rect 27982 35232 27988 35244
rect 28040 35232 28046 35284
rect 24118 35204 24124 35216
rect 20548 35176 22968 35204
rect 16666 35136 16672 35148
rect 15764 35108 16672 35136
rect 15764 35077 15792 35108
rect 16666 35096 16672 35108
rect 16724 35096 16730 35148
rect 15749 35071 15807 35077
rect 15749 35037 15761 35071
rect 15795 35037 15807 35071
rect 15749 35031 15807 35037
rect 15930 35028 15936 35080
rect 15988 35068 15994 35080
rect 16025 35071 16083 35077
rect 16025 35068 16037 35071
rect 15988 35040 16037 35068
rect 15988 35028 15994 35040
rect 16025 35037 16037 35040
rect 16071 35037 16083 35071
rect 18322 35068 18328 35080
rect 18283 35040 18328 35068
rect 16025 35031 16083 35037
rect 18322 35028 18328 35040
rect 18380 35028 18386 35080
rect 20548 35077 20576 35176
rect 21450 35096 21456 35148
rect 21508 35136 21514 35148
rect 22738 35136 22744 35148
rect 21508 35108 22744 35136
rect 21508 35096 21514 35108
rect 22738 35096 22744 35108
rect 22796 35096 22802 35148
rect 20533 35071 20591 35077
rect 20533 35037 20545 35071
rect 20579 35037 20591 35071
rect 21726 35068 21732 35080
rect 21687 35040 21732 35068
rect 20533 35031 20591 35037
rect 16574 34960 16580 35012
rect 16632 35000 16638 35012
rect 20548 35000 20576 35031
rect 21726 35028 21732 35040
rect 21784 35028 21790 35080
rect 21913 35071 21971 35077
rect 21913 35037 21925 35071
rect 21959 35037 21971 35071
rect 21913 35031 21971 35037
rect 22005 35071 22063 35077
rect 22005 35037 22017 35071
rect 22051 35068 22063 35071
rect 22830 35068 22836 35080
rect 22051 35040 22836 35068
rect 22051 35037 22063 35040
rect 22005 35031 22063 35037
rect 16632 34972 20576 35000
rect 21928 35000 21956 35031
rect 22830 35028 22836 35040
rect 22888 35028 22894 35080
rect 22094 35000 22100 35012
rect 21928 34972 22100 35000
rect 16632 34960 16638 34972
rect 22094 34960 22100 34972
rect 22152 34960 22158 35012
rect 18414 34932 18420 34944
rect 18375 34904 18420 34932
rect 18414 34892 18420 34904
rect 18472 34892 18478 34944
rect 21545 34935 21603 34941
rect 21545 34901 21557 34935
rect 21591 34932 21603 34935
rect 22278 34932 22284 34944
rect 21591 34904 22284 34932
rect 21591 34901 21603 34904
rect 21545 34895 21603 34901
rect 22278 34892 22284 34904
rect 22336 34892 22342 34944
rect 22940 34932 22968 35176
rect 23124 35176 24124 35204
rect 23017 35071 23075 35077
rect 23017 35037 23029 35071
rect 23063 35068 23075 35071
rect 23124 35068 23152 35176
rect 24118 35164 24124 35176
rect 24176 35204 24182 35216
rect 24489 35207 24547 35213
rect 24489 35204 24501 35207
rect 24176 35176 24501 35204
rect 24176 35164 24182 35176
rect 24489 35173 24501 35176
rect 24535 35204 24547 35207
rect 24535 35176 26280 35204
rect 24535 35173 24547 35176
rect 24489 35167 24547 35173
rect 26252 35148 26280 35176
rect 26326 35164 26332 35216
rect 26384 35204 26390 35216
rect 27433 35207 27491 35213
rect 27433 35204 27445 35207
rect 26384 35176 27445 35204
rect 26384 35164 26390 35176
rect 27433 35173 27445 35176
rect 27479 35173 27491 35207
rect 27433 35167 27491 35173
rect 24026 35136 24032 35148
rect 23216 35108 24032 35136
rect 23216 35077 23244 35108
rect 24026 35096 24032 35108
rect 24084 35096 24090 35148
rect 24673 35139 24731 35145
rect 24673 35105 24685 35139
rect 24719 35105 24731 35139
rect 24673 35099 24731 35105
rect 24398 35081 24456 35087
rect 23063 35040 23152 35068
rect 23201 35071 23259 35077
rect 23063 35037 23075 35040
rect 23017 35031 23075 35037
rect 23201 35037 23213 35071
rect 23247 35037 23259 35071
rect 23201 35031 23259 35037
rect 23477 35071 23535 35077
rect 23477 35037 23489 35071
rect 23523 35068 23535 35071
rect 23934 35068 23940 35080
rect 23523 35040 23940 35068
rect 23523 35037 23535 35040
rect 23477 35031 23535 35037
rect 23934 35028 23940 35040
rect 23992 35028 23998 35080
rect 24398 35078 24410 35081
rect 24320 35068 24410 35078
rect 24044 35050 24410 35068
rect 24044 35040 24348 35050
rect 24398 35047 24410 35050
rect 24444 35068 24456 35081
rect 24486 35068 24492 35080
rect 24444 35047 24492 35068
rect 24398 35041 24492 35047
rect 24428 35040 24492 35041
rect 23106 35000 23112 35012
rect 23067 34972 23112 35000
rect 23106 34960 23112 34972
rect 23164 34960 23170 35012
rect 23290 34960 23296 35012
rect 23348 35009 23354 35012
rect 23348 35003 23377 35009
rect 23365 35000 23377 35003
rect 24044 35000 24072 35040
rect 24486 35028 24492 35040
rect 24544 35028 24550 35080
rect 23365 34972 24072 35000
rect 23365 34969 23377 34972
rect 23348 34963 23377 34969
rect 23348 34960 23354 34963
rect 24688 34932 24716 35099
rect 24946 35096 24952 35148
rect 25004 35136 25010 35148
rect 25685 35139 25743 35145
rect 25685 35136 25697 35139
rect 25004 35108 25697 35136
rect 25004 35096 25010 35108
rect 25685 35105 25697 35108
rect 25731 35105 25743 35139
rect 25685 35099 25743 35105
rect 26234 35096 26240 35148
rect 26292 35136 26298 35148
rect 26292 35108 28396 35136
rect 26292 35096 26298 35108
rect 25406 35068 25412 35080
rect 25367 35040 25412 35068
rect 25406 35028 25412 35040
rect 25464 35028 25470 35080
rect 25501 35071 25559 35077
rect 25501 35037 25513 35071
rect 25547 35037 25559 35071
rect 25501 35031 25559 35037
rect 24762 34960 24768 35012
rect 24820 35000 24826 35012
rect 25516 35000 25544 35031
rect 25590 35028 25596 35080
rect 25648 35068 25654 35080
rect 25777 35071 25835 35077
rect 25777 35068 25789 35071
rect 25648 35040 25789 35068
rect 25648 35028 25654 35040
rect 25777 35037 25789 35040
rect 25823 35037 25835 35071
rect 25777 35031 25835 35037
rect 26329 35071 26387 35077
rect 26329 35037 26341 35071
rect 26375 35068 26387 35071
rect 26418 35068 26424 35080
rect 26375 35040 26424 35068
rect 26375 35037 26387 35040
rect 26329 35031 26387 35037
rect 26418 35028 26424 35040
rect 26476 35028 26482 35080
rect 27154 35068 27160 35080
rect 27115 35040 27160 35068
rect 27154 35028 27160 35040
rect 27212 35028 27218 35080
rect 27249 35071 27307 35077
rect 27249 35037 27261 35071
rect 27295 35037 27307 35071
rect 27249 35031 27307 35037
rect 24820 34972 25544 35000
rect 26973 35003 27031 35009
rect 24820 34960 24826 34972
rect 26973 34969 26985 35003
rect 27019 35000 27031 35003
rect 27062 35000 27068 35012
rect 27019 34972 27068 35000
rect 27019 34969 27031 34972
rect 26973 34963 27031 34969
rect 27062 34960 27068 34972
rect 27120 34960 27126 35012
rect 27264 35000 27292 35031
rect 27798 35028 27804 35080
rect 27856 35068 27862 35080
rect 28368 35077 28396 35108
rect 28077 35071 28135 35077
rect 28077 35068 28089 35071
rect 27856 35040 28089 35068
rect 27856 35028 27862 35040
rect 28077 35037 28089 35040
rect 28123 35037 28135 35071
rect 28077 35031 28135 35037
rect 28169 35071 28227 35077
rect 28169 35037 28181 35071
rect 28215 35037 28227 35071
rect 28169 35031 28227 35037
rect 28353 35071 28411 35077
rect 28353 35037 28365 35071
rect 28399 35037 28411 35071
rect 28353 35031 28411 35037
rect 28184 35000 28212 35031
rect 28442 35028 28448 35080
rect 28500 35068 28506 35080
rect 28500 35040 28545 35068
rect 28500 35028 28506 35040
rect 29822 35028 29828 35080
rect 29880 35068 29886 35080
rect 30009 35071 30067 35077
rect 30009 35068 30021 35071
rect 29880 35040 30021 35068
rect 29880 35028 29886 35040
rect 30009 35037 30021 35040
rect 30055 35037 30067 35071
rect 30374 35068 30380 35080
rect 30335 35040 30380 35068
rect 30009 35031 30067 35037
rect 30374 35028 30380 35040
rect 30432 35028 30438 35080
rect 48133 35071 48191 35077
rect 48133 35037 48145 35071
rect 48179 35068 48191 35071
rect 48222 35068 48228 35080
rect 48179 35040 48228 35068
rect 48179 35037 48191 35040
rect 48133 35031 48191 35037
rect 48222 35028 48228 35040
rect 48280 35028 48286 35080
rect 28902 35000 28908 35012
rect 27264 34972 28908 35000
rect 28902 34960 28908 34972
rect 28960 34960 28966 35012
rect 28994 34960 29000 35012
rect 29052 35000 29058 35012
rect 30193 35003 30251 35009
rect 30193 35000 30205 35003
rect 29052 34972 30205 35000
rect 29052 34960 29058 34972
rect 30193 34969 30205 34972
rect 30239 34969 30251 35003
rect 30193 34963 30251 34969
rect 30285 35003 30343 35009
rect 30285 34969 30297 35003
rect 30331 34969 30343 35003
rect 30285 34963 30343 34969
rect 26142 34932 26148 34944
rect 22940 34904 26148 34932
rect 26142 34892 26148 34904
rect 26200 34932 26206 34944
rect 26421 34935 26479 34941
rect 26421 34932 26433 34935
rect 26200 34904 26433 34932
rect 26200 34892 26206 34904
rect 26421 34901 26433 34904
rect 26467 34901 26479 34935
rect 26421 34895 26479 34901
rect 27893 34935 27951 34941
rect 27893 34901 27905 34935
rect 27939 34932 27951 34935
rect 28626 34932 28632 34944
rect 27939 34904 28632 34932
rect 27939 34901 27951 34904
rect 27893 34895 27951 34901
rect 28626 34892 28632 34904
rect 28684 34892 28690 34944
rect 29454 34892 29460 34944
rect 29512 34932 29518 34944
rect 30300 34932 30328 34963
rect 29512 34904 30328 34932
rect 30561 34935 30619 34941
rect 29512 34892 29518 34904
rect 30561 34901 30573 34935
rect 30607 34932 30619 34935
rect 30742 34932 30748 34944
rect 30607 34904 30748 34932
rect 30607 34901 30619 34904
rect 30561 34895 30619 34901
rect 30742 34892 30748 34904
rect 30800 34892 30806 34944
rect 47854 34892 47860 34944
rect 47912 34932 47918 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47912 34904 47961 34932
rect 47912 34892 47918 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 22094 34728 22100 34740
rect 21836 34700 22100 34728
rect 18414 34620 18420 34672
rect 18472 34620 18478 34672
rect 21266 34660 21272 34672
rect 20364 34632 21272 34660
rect 15289 34595 15347 34601
rect 15289 34561 15301 34595
rect 15335 34592 15347 34595
rect 16022 34592 16028 34604
rect 15335 34564 16028 34592
rect 15335 34561 15347 34564
rect 15289 34555 15347 34561
rect 16022 34552 16028 34564
rect 16080 34552 16086 34604
rect 17310 34552 17316 34604
rect 17368 34592 17374 34604
rect 20364 34601 20392 34632
rect 21266 34620 21272 34632
rect 21324 34620 21330 34672
rect 21836 34669 21864 34700
rect 22094 34688 22100 34700
rect 22152 34728 22158 34740
rect 23477 34731 23535 34737
rect 23477 34728 23489 34731
rect 22152 34700 23489 34728
rect 22152 34688 22158 34700
rect 23477 34697 23489 34700
rect 23523 34697 23535 34731
rect 26326 34728 26332 34740
rect 23477 34691 23535 34697
rect 24964 34700 26332 34728
rect 21821 34663 21879 34669
rect 21821 34629 21833 34663
rect 21867 34629 21879 34663
rect 21821 34623 21879 34629
rect 21910 34620 21916 34672
rect 21968 34660 21974 34672
rect 23109 34663 23167 34669
rect 21968 34632 23060 34660
rect 21968 34620 21974 34632
rect 17405 34595 17463 34601
rect 17405 34592 17417 34595
rect 17368 34564 17417 34592
rect 17368 34552 17374 34564
rect 17405 34561 17417 34564
rect 17451 34561 17463 34595
rect 17405 34555 17463 34561
rect 20349 34595 20407 34601
rect 20349 34561 20361 34595
rect 20395 34561 20407 34595
rect 20349 34555 20407 34561
rect 20533 34595 20591 34601
rect 20533 34561 20545 34595
rect 20579 34592 20591 34595
rect 20806 34592 20812 34604
rect 20579 34564 20812 34592
rect 20579 34561 20591 34564
rect 20533 34555 20591 34561
rect 20806 34552 20812 34564
rect 20864 34552 20870 34604
rect 20901 34595 20959 34601
rect 20901 34561 20913 34595
rect 20947 34592 20959 34595
rect 21450 34592 21456 34604
rect 20947 34564 21456 34592
rect 20947 34561 20959 34564
rect 20901 34555 20959 34561
rect 21450 34552 21456 34564
rect 21508 34552 21514 34604
rect 22097 34595 22155 34601
rect 22097 34592 22109 34595
rect 21744 34564 22109 34592
rect 17678 34524 17684 34536
rect 17639 34496 17684 34524
rect 17678 34484 17684 34496
rect 17736 34484 17742 34536
rect 20625 34527 20683 34533
rect 20625 34493 20637 34527
rect 20671 34493 20683 34527
rect 20625 34487 20683 34493
rect 20717 34527 20775 34533
rect 20717 34493 20729 34527
rect 20763 34524 20775 34527
rect 21174 34524 21180 34536
rect 20763 34496 21180 34524
rect 20763 34493 20775 34496
rect 20717 34487 20775 34493
rect 20640 34456 20668 34487
rect 21174 34484 21180 34496
rect 21232 34484 21238 34536
rect 21744 34468 21772 34564
rect 22097 34561 22109 34564
rect 22143 34561 22155 34595
rect 22097 34555 22155 34561
rect 22005 34527 22063 34533
rect 22005 34493 22017 34527
rect 22051 34524 22063 34527
rect 22051 34496 22140 34524
rect 22051 34493 22063 34496
rect 22005 34487 22063 34493
rect 22112 34468 22140 34496
rect 22830 34484 22836 34536
rect 22888 34524 22894 34536
rect 23032 34524 23060 34632
rect 23109 34629 23121 34663
rect 23155 34660 23167 34663
rect 23382 34660 23388 34672
rect 23155 34632 23388 34660
rect 23155 34629 23167 34632
rect 23109 34623 23167 34629
rect 23382 34620 23388 34632
rect 23440 34620 23446 34672
rect 23566 34620 23572 34672
rect 23624 34660 23630 34672
rect 24029 34663 24087 34669
rect 24029 34660 24041 34663
rect 23624 34632 24041 34660
rect 23624 34620 23630 34632
rect 24029 34629 24041 34632
rect 24075 34629 24087 34663
rect 24029 34623 24087 34629
rect 23293 34595 23351 34601
rect 23293 34561 23305 34595
rect 23339 34592 23351 34595
rect 24964 34592 24992 34700
rect 26326 34688 26332 34700
rect 26384 34688 26390 34740
rect 27062 34728 27068 34740
rect 26436 34700 27068 34728
rect 25038 34620 25044 34672
rect 25096 34660 25102 34672
rect 25225 34663 25283 34669
rect 25225 34660 25237 34663
rect 25096 34632 25237 34660
rect 25096 34620 25102 34632
rect 25225 34629 25237 34632
rect 25271 34660 25283 34663
rect 25590 34660 25596 34672
rect 25271 34632 25596 34660
rect 25271 34629 25283 34632
rect 25225 34623 25283 34629
rect 25590 34620 25596 34632
rect 25648 34620 25654 34672
rect 26436 34660 26464 34700
rect 27062 34688 27068 34700
rect 27120 34688 27126 34740
rect 27341 34731 27399 34737
rect 27341 34697 27353 34731
rect 27387 34728 27399 34731
rect 27430 34728 27436 34740
rect 27387 34700 27436 34728
rect 27387 34697 27399 34700
rect 27341 34691 27399 34697
rect 27430 34688 27436 34700
rect 27488 34688 27494 34740
rect 29362 34728 29368 34740
rect 29323 34700 29368 34728
rect 29362 34688 29368 34700
rect 29420 34688 29426 34740
rect 26160 34632 26464 34660
rect 26160 34601 26188 34632
rect 26510 34620 26516 34672
rect 26568 34660 26574 34672
rect 29454 34660 29460 34672
rect 26568 34632 29460 34660
rect 26568 34620 26574 34632
rect 29454 34620 29460 34632
rect 29512 34620 29518 34672
rect 30929 34663 30987 34669
rect 30929 34629 30941 34663
rect 30975 34660 30987 34663
rect 31386 34660 31392 34672
rect 30975 34632 31392 34660
rect 30975 34629 30987 34632
rect 30929 34623 30987 34629
rect 31386 34620 31392 34632
rect 31444 34620 31450 34672
rect 23339 34564 24992 34592
rect 26145 34595 26203 34601
rect 23339 34561 23351 34564
rect 23293 34555 23351 34561
rect 26145 34561 26157 34595
rect 26191 34561 26203 34595
rect 26970 34592 26976 34604
rect 26931 34564 26976 34592
rect 26145 34555 26203 34561
rect 26970 34552 26976 34564
rect 27028 34552 27034 34604
rect 27154 34592 27160 34604
rect 27115 34564 27160 34592
rect 27154 34552 27160 34564
rect 27212 34552 27218 34604
rect 28626 34592 28632 34604
rect 28587 34564 28632 34592
rect 28626 34552 28632 34564
rect 28684 34552 28690 34604
rect 28813 34595 28871 34601
rect 28813 34561 28825 34595
rect 28859 34561 28871 34595
rect 28813 34555 28871 34561
rect 25406 34524 25412 34536
rect 22888 34496 22968 34524
rect 23032 34496 25412 34524
rect 22888 34484 22894 34496
rect 21726 34456 21732 34468
rect 20640 34428 21732 34456
rect 21726 34416 21732 34428
rect 21784 34416 21790 34468
rect 22094 34416 22100 34468
rect 22152 34416 22158 34468
rect 22940 34456 22968 34496
rect 25406 34484 25412 34496
rect 25464 34484 25470 34536
rect 25516 34496 26188 34524
rect 24213 34459 24271 34465
rect 24213 34456 24225 34459
rect 22940 34428 24225 34456
rect 24213 34425 24225 34428
rect 24259 34456 24271 34459
rect 25516 34456 25544 34496
rect 24259 34428 25544 34456
rect 26160 34456 26188 34496
rect 26234 34484 26240 34536
rect 26292 34524 26298 34536
rect 26421 34527 26479 34533
rect 26421 34524 26433 34527
rect 26292 34496 26433 34524
rect 26292 34484 26298 34496
rect 26421 34493 26433 34496
rect 26467 34524 26479 34527
rect 27172 34524 27200 34552
rect 26467 34496 27200 34524
rect 26467 34493 26479 34496
rect 26421 34487 26479 34493
rect 28534 34484 28540 34536
rect 28592 34524 28598 34536
rect 28828 34524 28856 34555
rect 28902 34552 28908 34604
rect 28960 34592 28966 34604
rect 29178 34592 29184 34604
rect 28960 34564 29005 34592
rect 29139 34564 29184 34592
rect 28960 34552 28966 34564
rect 29178 34552 29184 34564
rect 29236 34552 29242 34604
rect 30742 34592 30748 34604
rect 30703 34564 30748 34592
rect 30742 34552 30748 34564
rect 30800 34552 30806 34604
rect 31018 34552 31024 34604
rect 31076 34592 31082 34604
rect 47762 34592 47768 34604
rect 31076 34564 31121 34592
rect 47723 34564 47768 34592
rect 31076 34552 31082 34564
rect 47762 34552 47768 34564
rect 47820 34552 47826 34604
rect 28592 34496 28856 34524
rect 28997 34527 29055 34533
rect 28592 34484 28598 34496
rect 28997 34493 29009 34527
rect 29043 34524 29055 34527
rect 29270 34524 29276 34536
rect 29043 34496 29276 34524
rect 29043 34493 29055 34496
rect 28997 34487 29055 34493
rect 29270 34484 29276 34496
rect 29328 34484 29334 34536
rect 26510 34456 26516 34468
rect 26160 34428 26516 34456
rect 24259 34425 24271 34428
rect 24213 34419 24271 34425
rect 15381 34391 15439 34397
rect 15381 34357 15393 34391
rect 15427 34388 15439 34391
rect 15470 34388 15476 34400
rect 15427 34360 15476 34388
rect 15427 34357 15439 34360
rect 15381 34351 15439 34357
rect 15470 34348 15476 34360
rect 15528 34348 15534 34400
rect 19058 34348 19064 34400
rect 19116 34388 19122 34400
rect 19153 34391 19211 34397
rect 19153 34388 19165 34391
rect 19116 34360 19165 34388
rect 19116 34348 19122 34360
rect 19153 34357 19165 34360
rect 19199 34357 19211 34391
rect 19153 34351 19211 34357
rect 20714 34348 20720 34400
rect 20772 34388 20778 34400
rect 21085 34391 21143 34397
rect 21085 34388 21097 34391
rect 20772 34360 21097 34388
rect 20772 34348 20778 34360
rect 21085 34357 21097 34360
rect 21131 34357 21143 34391
rect 21818 34388 21824 34400
rect 21779 34360 21824 34388
rect 21085 34351 21143 34357
rect 21818 34348 21824 34360
rect 21876 34348 21882 34400
rect 22186 34348 22192 34400
rect 22244 34388 22250 34400
rect 26252 34397 26280 34428
rect 26510 34416 26516 34428
rect 26568 34456 26574 34468
rect 26970 34456 26976 34468
rect 26568 34428 26976 34456
rect 26568 34416 26574 34428
rect 26970 34416 26976 34428
rect 27028 34416 27034 34468
rect 22281 34391 22339 34397
rect 22281 34388 22293 34391
rect 22244 34360 22293 34388
rect 22244 34348 22250 34360
rect 22281 34357 22293 34360
rect 22327 34357 22339 34391
rect 22281 34351 22339 34357
rect 26237 34391 26295 34397
rect 26237 34357 26249 34391
rect 26283 34357 26295 34391
rect 26237 34351 26295 34357
rect 26329 34391 26387 34397
rect 26329 34357 26341 34391
rect 26375 34388 26387 34391
rect 26878 34388 26884 34400
rect 26375 34360 26884 34388
rect 26375 34357 26387 34360
rect 26329 34351 26387 34357
rect 26878 34348 26884 34360
rect 26936 34348 26942 34400
rect 27062 34388 27068 34400
rect 27023 34360 27068 34388
rect 27062 34348 27068 34360
rect 27120 34348 27126 34400
rect 30558 34388 30564 34400
rect 30519 34360 30564 34388
rect 30558 34348 30564 34360
rect 30616 34348 30622 34400
rect 47210 34348 47216 34400
rect 47268 34388 47274 34400
rect 47581 34391 47639 34397
rect 47581 34388 47593 34391
rect 47268 34360 47593 34388
rect 47268 34348 47274 34360
rect 47581 34357 47593 34360
rect 47627 34357 47639 34391
rect 47581 34351 47639 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1946 34144 1952 34196
rect 2004 34184 2010 34196
rect 2004 34156 17448 34184
rect 2004 34144 2010 34156
rect 17310 34116 17316 34128
rect 16776 34088 17316 34116
rect 14185 34051 14243 34057
rect 14185 34017 14197 34051
rect 14231 34048 14243 34051
rect 16776 34048 16804 34088
rect 17310 34076 17316 34088
rect 17368 34076 17374 34128
rect 17420 34116 17448 34156
rect 17678 34144 17684 34196
rect 17736 34184 17742 34196
rect 18509 34187 18567 34193
rect 18509 34184 18521 34187
rect 17736 34156 18521 34184
rect 17736 34144 17742 34156
rect 18509 34153 18521 34156
rect 18555 34153 18567 34187
rect 21726 34184 21732 34196
rect 21687 34156 21732 34184
rect 18509 34147 18567 34153
rect 21726 34144 21732 34156
rect 21784 34144 21790 34196
rect 22278 34184 22284 34196
rect 22239 34156 22284 34184
rect 22278 34144 22284 34156
rect 22336 34144 22342 34196
rect 23566 34184 23572 34196
rect 23527 34156 23572 34184
rect 23566 34144 23572 34156
rect 23624 34144 23630 34196
rect 24486 34144 24492 34196
rect 24544 34184 24550 34196
rect 24581 34187 24639 34193
rect 24581 34184 24593 34187
rect 24544 34156 24593 34184
rect 24544 34144 24550 34156
rect 24581 34153 24593 34156
rect 24627 34184 24639 34187
rect 24670 34184 24676 34196
rect 24627 34156 24676 34184
rect 24627 34153 24639 34156
rect 24581 34147 24639 34153
rect 24670 34144 24676 34156
rect 24728 34144 24734 34196
rect 30374 34184 30380 34196
rect 27448 34156 30380 34184
rect 17420 34088 18184 34116
rect 14231 34020 16804 34048
rect 14231 34017 14243 34020
rect 14185 34011 14243 34017
rect 16850 34008 16856 34060
rect 16908 34048 16914 34060
rect 18156 34057 18184 34088
rect 21266 34076 21272 34128
rect 21324 34116 21330 34128
rect 22741 34119 22799 34125
rect 22741 34116 22753 34119
rect 21324 34088 22753 34116
rect 21324 34076 21330 34088
rect 22741 34085 22753 34088
rect 22787 34085 22799 34119
rect 27448 34116 27476 34156
rect 30374 34144 30380 34156
rect 30432 34144 30438 34196
rect 30558 34144 30564 34196
rect 30616 34184 30622 34196
rect 31094 34187 31152 34193
rect 31094 34184 31106 34187
rect 30616 34156 31106 34184
rect 30616 34144 30622 34156
rect 31094 34153 31106 34156
rect 31140 34153 31152 34187
rect 31094 34147 31152 34153
rect 22741 34079 22799 34085
rect 23400 34088 27476 34116
rect 18141 34051 18199 34057
rect 16908 34020 16953 34048
rect 16908 34008 16914 34020
rect 18141 34017 18153 34051
rect 18187 34017 18199 34051
rect 19978 34048 19984 34060
rect 19939 34020 19984 34048
rect 18141 34011 18199 34017
rect 19978 34008 19984 34020
rect 20036 34008 20042 34060
rect 20257 34051 20315 34057
rect 20257 34017 20269 34051
rect 20303 34048 20315 34051
rect 20714 34048 20720 34060
rect 20303 34020 20720 34048
rect 20303 34017 20315 34020
rect 20257 34011 20315 34017
rect 20714 34008 20720 34020
rect 20772 34008 20778 34060
rect 21818 34048 21824 34060
rect 21731 34020 21824 34048
rect 1578 33980 1584 33992
rect 1539 33952 1584 33980
rect 1578 33940 1584 33952
rect 1636 33940 1642 33992
rect 16574 33980 16580 33992
rect 16535 33952 16580 33980
rect 16574 33940 16580 33952
rect 16632 33940 16638 33992
rect 16669 33983 16727 33989
rect 16669 33949 16681 33983
rect 16715 33949 16727 33983
rect 16942 33980 16948 33992
rect 16903 33952 16948 33980
rect 16669 33943 16727 33949
rect 14458 33912 14464 33924
rect 14419 33884 14464 33912
rect 14458 33872 14464 33884
rect 14516 33872 14522 33924
rect 15470 33872 15476 33924
rect 15528 33872 15534 33924
rect 16298 33912 16304 33924
rect 15948 33884 16304 33912
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 1946 33844 1952 33856
rect 1443 33816 1952 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 1946 33804 1952 33816
rect 2004 33804 2010 33856
rect 15948 33853 15976 33884
rect 16298 33872 16304 33884
rect 16356 33912 16362 33924
rect 16684 33912 16712 33943
rect 16942 33940 16948 33952
rect 17000 33940 17006 33992
rect 17770 33980 17776 33992
rect 17731 33952 17776 33980
rect 17770 33940 17776 33952
rect 17828 33940 17834 33992
rect 17954 33980 17960 33992
rect 17915 33952 17960 33980
rect 17954 33940 17960 33952
rect 18012 33940 18018 33992
rect 18049 33983 18107 33989
rect 18049 33949 18061 33983
rect 18095 33949 18107 33983
rect 18322 33980 18328 33992
rect 18283 33952 18328 33980
rect 18049 33943 18107 33949
rect 16356 33884 16712 33912
rect 18064 33912 18092 33943
rect 18322 33940 18328 33952
rect 18380 33940 18386 33992
rect 19058 33912 19064 33924
rect 18064 33884 19064 33912
rect 16356 33872 16362 33884
rect 19058 33872 19064 33884
rect 19116 33872 19122 33924
rect 20990 33872 20996 33924
rect 21048 33872 21054 33924
rect 15933 33847 15991 33853
rect 15933 33813 15945 33847
rect 15979 33813 15991 33847
rect 16390 33844 16396 33856
rect 16351 33816 16396 33844
rect 15933 33807 15991 33813
rect 16390 33804 16396 33816
rect 16448 33804 16454 33856
rect 20070 33804 20076 33856
rect 20128 33844 20134 33856
rect 21744 33844 21772 34020
rect 21818 34008 21824 34020
rect 21876 34048 21882 34060
rect 23400 34048 23428 34088
rect 27522 34076 27528 34128
rect 27580 34116 27586 34128
rect 27580 34088 30880 34116
rect 27580 34076 27586 34088
rect 21876 34020 23428 34048
rect 21876 34008 21882 34020
rect 22002 33940 22008 33992
rect 22060 33980 22066 33992
rect 22189 33983 22247 33989
rect 22189 33980 22201 33983
rect 22060 33952 22201 33980
rect 22060 33940 22066 33952
rect 22189 33949 22201 33952
rect 22235 33949 22247 33983
rect 22462 33980 22468 33992
rect 22423 33952 22468 33980
rect 22189 33943 22247 33949
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 22094 33872 22100 33924
rect 22152 33912 22158 33924
rect 23400 33921 23428 34020
rect 26421 34051 26479 34057
rect 26421 34017 26433 34051
rect 26467 34048 26479 34051
rect 27338 34048 27344 34060
rect 26467 34020 27344 34048
rect 26467 34017 26479 34020
rect 26421 34011 26479 34017
rect 27338 34008 27344 34020
rect 27396 34008 27402 34060
rect 29914 34048 29920 34060
rect 29875 34020 29920 34048
rect 29914 34008 29920 34020
rect 29972 34008 29978 34060
rect 30852 34057 30880 34088
rect 30837 34051 30895 34057
rect 30837 34017 30849 34051
rect 30883 34048 30895 34051
rect 32122 34048 32128 34060
rect 30883 34020 32128 34048
rect 30883 34017 30895 34020
rect 30837 34011 30895 34017
rect 32122 34008 32128 34020
rect 32180 34008 32186 34060
rect 47118 34048 47124 34060
rect 47079 34020 47124 34048
rect 47118 34008 47124 34020
rect 47176 34008 47182 34060
rect 47394 34048 47400 34060
rect 47355 34020 47400 34048
rect 47394 34008 47400 34020
rect 47452 34008 47458 34060
rect 24397 33983 24455 33989
rect 24397 33949 24409 33983
rect 24443 33980 24455 33983
rect 24578 33980 24584 33992
rect 24443 33952 24584 33980
rect 24443 33949 24455 33952
rect 24397 33943 24455 33949
rect 24578 33940 24584 33952
rect 24636 33940 24642 33992
rect 26142 33980 26148 33992
rect 26103 33952 26148 33980
rect 26142 33940 26148 33952
rect 26200 33940 26206 33992
rect 26234 33940 26240 33992
rect 26292 33980 26298 33992
rect 26513 33983 26571 33989
rect 26292 33952 26337 33980
rect 26292 33940 26298 33952
rect 26513 33949 26525 33983
rect 26559 33949 26571 33983
rect 26513 33943 26571 33949
rect 23201 33915 23259 33921
rect 23201 33912 23213 33915
rect 22152 33884 23213 33912
rect 22152 33872 22158 33884
rect 23201 33881 23213 33884
rect 23247 33881 23259 33915
rect 23201 33875 23259 33881
rect 23385 33915 23443 33921
rect 23385 33881 23397 33915
rect 23431 33881 23443 33915
rect 23385 33875 23443 33881
rect 25406 33872 25412 33924
rect 25464 33912 25470 33924
rect 26528 33912 26556 33943
rect 26878 33940 26884 33992
rect 26936 33980 26942 33992
rect 26973 33983 27031 33989
rect 26973 33980 26985 33983
rect 26936 33952 26985 33980
rect 26936 33940 26942 33952
rect 26973 33949 26985 33952
rect 27019 33949 27031 33983
rect 26973 33943 27031 33949
rect 27157 33983 27215 33989
rect 27157 33949 27169 33983
rect 27203 33980 27215 33983
rect 27430 33980 27436 33992
rect 27203 33952 27436 33980
rect 27203 33949 27215 33952
rect 27157 33943 27215 33949
rect 27430 33940 27436 33952
rect 27488 33940 27494 33992
rect 29822 33940 29828 33992
rect 29880 33980 29886 33992
rect 30009 33983 30067 33989
rect 30009 33980 30021 33983
rect 29880 33952 30021 33980
rect 29880 33940 29886 33952
rect 30009 33949 30021 33952
rect 30055 33949 30067 33983
rect 30009 33943 30067 33949
rect 25464 33884 26556 33912
rect 30024 33912 30052 33943
rect 32858 33912 32864 33924
rect 30024 33884 31156 33912
rect 32338 33884 32864 33912
rect 25464 33872 25470 33884
rect 25958 33844 25964 33856
rect 20128 33816 21772 33844
rect 25919 33816 25964 33844
rect 20128 33804 20134 33816
rect 25958 33804 25964 33816
rect 26016 33804 26022 33856
rect 26142 33804 26148 33856
rect 26200 33844 26206 33856
rect 27065 33847 27123 33853
rect 27065 33844 27077 33847
rect 26200 33816 27077 33844
rect 26200 33804 26206 33816
rect 27065 33813 27077 33816
rect 27111 33813 27123 33847
rect 27065 33807 27123 33813
rect 30377 33847 30435 33853
rect 30377 33813 30389 33847
rect 30423 33844 30435 33847
rect 31018 33844 31024 33856
rect 30423 33816 31024 33844
rect 30423 33813 30435 33816
rect 30377 33807 30435 33813
rect 31018 33804 31024 33816
rect 31076 33804 31082 33856
rect 31128 33844 31156 33884
rect 32858 33872 32864 33884
rect 32916 33872 32922 33924
rect 47210 33872 47216 33924
rect 47268 33912 47274 33924
rect 47268 33884 47313 33912
rect 47268 33872 47274 33884
rect 32582 33844 32588 33856
rect 31128 33816 32588 33844
rect 32582 33804 32588 33816
rect 32640 33804 32646 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 14458 33600 14464 33652
rect 14516 33640 14522 33652
rect 15105 33643 15163 33649
rect 15105 33640 15117 33643
rect 14516 33612 15117 33640
rect 14516 33600 14522 33612
rect 15105 33609 15117 33612
rect 15151 33609 15163 33643
rect 15105 33603 15163 33609
rect 17770 33600 17776 33652
rect 17828 33640 17834 33652
rect 18417 33643 18475 33649
rect 18417 33640 18429 33643
rect 17828 33612 18429 33640
rect 17828 33600 17834 33612
rect 18417 33609 18429 33612
rect 18463 33609 18475 33643
rect 18417 33603 18475 33609
rect 19978 33600 19984 33652
rect 20036 33640 20042 33652
rect 20622 33640 20628 33652
rect 20036 33612 20628 33640
rect 20036 33600 20042 33612
rect 20622 33600 20628 33612
rect 20680 33640 20686 33652
rect 20717 33643 20775 33649
rect 20717 33640 20729 33643
rect 20680 33612 20729 33640
rect 20680 33600 20686 33612
rect 20717 33609 20729 33612
rect 20763 33609 20775 33643
rect 27433 33643 27491 33649
rect 20717 33603 20775 33609
rect 20824 33612 26004 33640
rect 15746 33572 15752 33584
rect 14660 33544 15752 33572
rect 14458 33504 14464 33516
rect 14419 33476 14464 33504
rect 14458 33464 14464 33476
rect 14516 33464 14522 33516
rect 14660 33513 14688 33544
rect 15746 33532 15752 33544
rect 15804 33532 15810 33584
rect 20824 33572 20852 33612
rect 22186 33572 22192 33584
rect 17880 33544 20852 33572
rect 21928 33544 22192 33572
rect 17880 33516 17908 33544
rect 14645 33507 14703 33513
rect 14645 33473 14657 33507
rect 14691 33473 14703 33507
rect 14645 33467 14703 33473
rect 15289 33507 15347 33513
rect 15289 33473 15301 33507
rect 15335 33504 15347 33507
rect 16390 33504 16396 33516
rect 15335 33476 16396 33504
rect 15335 33473 15347 33476
rect 15289 33467 15347 33473
rect 16390 33464 16396 33476
rect 16448 33464 16454 33516
rect 17862 33504 17868 33516
rect 17775 33476 17868 33504
rect 17862 33464 17868 33476
rect 17920 33464 17926 33516
rect 18233 33507 18291 33513
rect 18233 33473 18245 33507
rect 18279 33504 18291 33507
rect 18877 33507 18935 33513
rect 18877 33504 18889 33507
rect 18279 33476 18889 33504
rect 18279 33473 18291 33476
rect 18233 33467 18291 33473
rect 18877 33473 18889 33476
rect 18923 33473 18935 33507
rect 19058 33504 19064 33516
rect 19019 33476 19064 33504
rect 18877 33467 18935 33473
rect 19058 33464 19064 33476
rect 19116 33464 19122 33516
rect 19242 33464 19248 33516
rect 19300 33504 19306 33516
rect 19337 33507 19395 33513
rect 19337 33504 19349 33507
rect 19300 33476 19349 33504
rect 19300 33464 19306 33476
rect 19337 33473 19349 33476
rect 19383 33473 19395 33507
rect 20346 33504 20352 33516
rect 19337 33467 19395 33473
rect 19444 33476 20352 33504
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 1854 33436 1860 33448
rect 1719 33408 1860 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 1854 33396 1860 33408
rect 1912 33396 1918 33448
rect 15565 33439 15623 33445
rect 15565 33405 15577 33439
rect 15611 33436 15623 33439
rect 15930 33436 15936 33448
rect 15611 33408 15936 33436
rect 15611 33405 15623 33408
rect 15565 33399 15623 33405
rect 15930 33396 15936 33408
rect 15988 33436 15994 33448
rect 19444 33436 19472 33476
rect 20346 33464 20352 33476
rect 20404 33464 20410 33516
rect 20625 33507 20683 33513
rect 20625 33473 20637 33507
rect 20671 33504 20683 33507
rect 21634 33504 21640 33516
rect 20671 33476 21640 33504
rect 20671 33473 20683 33476
rect 20625 33467 20683 33473
rect 21634 33464 21640 33476
rect 21692 33464 21698 33516
rect 21821 33507 21879 33513
rect 21821 33473 21833 33507
rect 21867 33504 21879 33507
rect 21928 33504 21956 33544
rect 22186 33532 22192 33544
rect 22244 33532 22250 33584
rect 25976 33572 26004 33612
rect 27433 33609 27445 33643
rect 27479 33640 27491 33643
rect 27522 33640 27528 33652
rect 27479 33612 27528 33640
rect 27479 33609 27491 33612
rect 27433 33603 27491 33609
rect 27522 33600 27528 33612
rect 27580 33600 27586 33652
rect 30009 33643 30067 33649
rect 30009 33640 30021 33643
rect 28966 33612 30021 33640
rect 28966 33572 28994 33612
rect 30009 33609 30021 33612
rect 30055 33609 30067 33643
rect 32858 33640 32864 33652
rect 32819 33612 32864 33640
rect 30009 33603 30067 33609
rect 32858 33600 32864 33612
rect 32916 33600 32922 33652
rect 47762 33600 47768 33652
rect 47820 33640 47826 33652
rect 48041 33643 48099 33649
rect 48041 33640 48053 33643
rect 47820 33612 48053 33640
rect 47820 33600 47826 33612
rect 48041 33609 48053 33612
rect 48087 33609 48099 33643
rect 48041 33603 48099 33609
rect 25976 33544 28994 33572
rect 29362 33532 29368 33584
rect 29420 33572 29426 33584
rect 29420 33544 29465 33572
rect 29420 33532 29426 33544
rect 21867 33476 21956 33504
rect 21867 33473 21879 33476
rect 21821 33467 21879 33473
rect 22002 33464 22008 33516
rect 22060 33504 22066 33516
rect 22097 33507 22155 33513
rect 22097 33504 22109 33507
rect 22060 33476 22109 33504
rect 22060 33464 22066 33476
rect 22097 33473 22109 33476
rect 22143 33473 22155 33507
rect 22097 33467 22155 33473
rect 24213 33507 24271 33513
rect 24213 33473 24225 33507
rect 24259 33504 24271 33507
rect 24578 33504 24584 33516
rect 24259 33476 24584 33504
rect 24259 33473 24271 33476
rect 24213 33467 24271 33473
rect 24578 33464 24584 33476
rect 24636 33464 24642 33516
rect 25958 33504 25964 33516
rect 25919 33476 25964 33504
rect 25958 33464 25964 33476
rect 26016 33464 26022 33516
rect 26142 33504 26148 33516
rect 26103 33476 26148 33504
rect 26142 33464 26148 33476
rect 26200 33464 26206 33516
rect 27341 33507 27399 33513
rect 27341 33473 27353 33507
rect 27387 33504 27399 33507
rect 27522 33504 27528 33516
rect 27387 33476 27528 33504
rect 27387 33473 27399 33476
rect 27341 33467 27399 33473
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 27985 33507 28043 33513
rect 27985 33473 27997 33507
rect 28031 33504 28043 33507
rect 28350 33504 28356 33516
rect 28031 33476 28356 33504
rect 28031 33473 28043 33476
rect 27985 33467 28043 33473
rect 28350 33464 28356 33476
rect 28408 33464 28414 33516
rect 29704 33507 29762 33513
rect 29704 33473 29716 33507
rect 29750 33504 29762 33507
rect 30006 33504 30012 33516
rect 29750 33502 29776 33504
rect 29840 33502 30012 33504
rect 29750 33476 30012 33502
rect 29750 33474 29868 33476
rect 29750 33473 29762 33474
rect 29704 33467 29762 33473
rect 30006 33464 30012 33476
rect 30064 33464 30070 33516
rect 32125 33507 32183 33513
rect 32125 33473 32137 33507
rect 32171 33504 32183 33507
rect 32306 33504 32312 33516
rect 32171 33476 32312 33504
rect 32171 33473 32183 33476
rect 32125 33467 32183 33473
rect 32306 33464 32312 33476
rect 32364 33464 32370 33516
rect 32769 33507 32827 33513
rect 32769 33473 32781 33507
rect 32815 33504 32827 33507
rect 32858 33504 32864 33516
rect 32815 33476 32864 33504
rect 32815 33473 32827 33476
rect 32769 33467 32827 33473
rect 32858 33464 32864 33476
rect 32916 33464 32922 33516
rect 46842 33504 46848 33516
rect 46803 33476 46848 33504
rect 46842 33464 46848 33476
rect 46900 33464 46906 33516
rect 47581 33507 47639 33513
rect 47581 33473 47593 33507
rect 47627 33473 47639 33507
rect 47581 33467 47639 33473
rect 15988 33408 19472 33436
rect 15988 33396 15994 33408
rect 19978 33396 19984 33448
rect 20036 33436 20042 33448
rect 20036 33408 24440 33436
rect 20036 33396 20042 33408
rect 14553 33371 14611 33377
rect 14553 33337 14565 33371
rect 14599 33368 14611 33371
rect 15473 33371 15531 33377
rect 15473 33368 15485 33371
rect 14599 33340 15485 33368
rect 14599 33337 14611 33340
rect 14553 33331 14611 33337
rect 15473 33337 15485 33340
rect 15519 33337 15531 33371
rect 22462 33368 22468 33380
rect 15473 33331 15531 33337
rect 18248 33340 22468 33368
rect 18248 33312 18276 33340
rect 22462 33328 22468 33340
rect 22520 33368 22526 33380
rect 23106 33368 23112 33380
rect 22520 33340 23112 33368
rect 22520 33328 22526 33340
rect 23106 33328 23112 33340
rect 23164 33328 23170 33380
rect 24412 33377 24440 33408
rect 25590 33396 25596 33448
rect 25648 33436 25654 33448
rect 25648 33408 25968 33436
rect 25648 33396 25654 33408
rect 24397 33371 24455 33377
rect 24397 33337 24409 33371
rect 24443 33368 24455 33371
rect 25940 33368 25968 33408
rect 26050 33396 26056 33448
rect 26108 33436 26114 33448
rect 26237 33439 26295 33445
rect 26237 33436 26249 33439
rect 26108 33408 26249 33436
rect 26108 33396 26114 33408
rect 26237 33405 26249 33408
rect 26283 33405 26295 33439
rect 26237 33399 26295 33405
rect 46658 33396 46664 33448
rect 46716 33436 46722 33448
rect 47596 33436 47624 33467
rect 46716 33408 47624 33436
rect 46716 33396 46722 33408
rect 28169 33371 28227 33377
rect 28169 33368 28181 33371
rect 24443 33340 25912 33368
rect 25940 33340 28181 33368
rect 24443 33337 24455 33340
rect 24397 33331 24455 33337
rect 18230 33300 18236 33312
rect 18143 33272 18236 33300
rect 18230 33260 18236 33272
rect 18288 33260 18294 33312
rect 19245 33303 19303 33309
rect 19245 33269 19257 33303
rect 19291 33300 19303 33303
rect 20070 33300 20076 33312
rect 19291 33272 20076 33300
rect 19291 33269 19303 33272
rect 19245 33263 19303 33269
rect 20070 33260 20076 33272
rect 20128 33260 20134 33312
rect 21542 33260 21548 33312
rect 21600 33300 21606 33312
rect 25590 33300 25596 33312
rect 21600 33272 25596 33300
rect 21600 33260 21606 33272
rect 25590 33260 25596 33272
rect 25648 33260 25654 33312
rect 25682 33260 25688 33312
rect 25740 33300 25746 33312
rect 25777 33303 25835 33309
rect 25777 33300 25789 33303
rect 25740 33272 25789 33300
rect 25740 33260 25746 33272
rect 25777 33269 25789 33272
rect 25823 33269 25835 33303
rect 25884 33300 25912 33340
rect 28169 33337 28181 33340
rect 28215 33368 28227 33371
rect 28626 33368 28632 33380
rect 28215 33340 28632 33368
rect 28215 33337 28227 33340
rect 28169 33331 28227 33337
rect 28626 33328 28632 33340
rect 28684 33328 28690 33380
rect 31386 33368 31392 33380
rect 29472 33340 31392 33368
rect 29472 33300 29500 33340
rect 31386 33328 31392 33340
rect 31444 33328 31450 33380
rect 29546 33309 29552 33312
rect 25884 33272 29500 33300
rect 29530 33303 29552 33309
rect 25777 33263 25835 33269
rect 29530 33269 29542 33303
rect 29530 33263 29552 33269
rect 29546 33260 29552 33263
rect 29604 33260 29610 33312
rect 29641 33303 29699 33309
rect 29641 33269 29653 33303
rect 29687 33300 29699 33303
rect 29914 33300 29920 33312
rect 29687 33272 29920 33300
rect 29687 33269 29699 33272
rect 29641 33263 29699 33269
rect 29914 33260 29920 33272
rect 29972 33260 29978 33312
rect 32214 33300 32220 33312
rect 32175 33272 32220 33300
rect 32214 33260 32220 33272
rect 32272 33260 32278 33312
rect 44174 33260 44180 33312
rect 44232 33300 44238 33312
rect 46937 33303 46995 33309
rect 46937 33300 46949 33303
rect 44232 33272 46949 33300
rect 44232 33260 44238 33272
rect 46937 33269 46949 33272
rect 46983 33269 46995 33303
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 46937 33263 46995 33269
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1946 33096 1952 33108
rect 1907 33068 1952 33096
rect 1946 33056 1952 33068
rect 2004 33056 2010 33108
rect 14458 33056 14464 33108
rect 14516 33096 14522 33108
rect 14829 33099 14887 33105
rect 14829 33096 14841 33099
rect 14516 33068 14841 33096
rect 14516 33056 14522 33068
rect 14829 33065 14841 33068
rect 14875 33065 14887 33099
rect 14829 33059 14887 33065
rect 15381 33099 15439 33105
rect 15381 33065 15393 33099
rect 15427 33065 15439 33099
rect 15930 33096 15936 33108
rect 15381 33059 15439 33065
rect 15488 33068 15936 33096
rect 15396 33028 15424 33059
rect 14660 33000 15424 33028
rect 2317 32963 2375 32969
rect 2317 32929 2329 32963
rect 2363 32929 2375 32963
rect 2317 32923 2375 32929
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32892 1915 32895
rect 1946 32892 1952 32904
rect 1903 32864 1952 32892
rect 1903 32861 1915 32864
rect 1857 32855 1915 32861
rect 1946 32852 1952 32864
rect 2004 32852 2010 32904
rect 2332 32892 2360 32923
rect 2961 32895 3019 32901
rect 2961 32892 2973 32895
rect 2332 32864 2973 32892
rect 2961 32861 2973 32864
rect 3007 32861 3019 32895
rect 2961 32855 3019 32861
rect 14458 32852 14464 32904
rect 14516 32892 14522 32904
rect 14660 32901 14688 33000
rect 15488 32969 15516 33068
rect 15930 33056 15936 33068
rect 15988 33096 15994 33108
rect 17126 33096 17132 33108
rect 15988 33068 16436 33096
rect 17087 33068 17132 33096
rect 15988 33056 15994 33068
rect 16408 33040 16436 33068
rect 17126 33056 17132 33068
rect 17184 33056 17190 33108
rect 17310 33056 17316 33108
rect 17368 33096 17374 33108
rect 18049 33099 18107 33105
rect 18049 33096 18061 33099
rect 17368 33068 18061 33096
rect 17368 33056 17374 33068
rect 18049 33065 18061 33068
rect 18095 33065 18107 33099
rect 18049 33059 18107 33065
rect 20990 33056 20996 33108
rect 21048 33096 21054 33108
rect 21085 33099 21143 33105
rect 21085 33096 21097 33099
rect 21048 33068 21097 33096
rect 21048 33056 21054 33068
rect 21085 33065 21097 33068
rect 21131 33065 21143 33099
rect 21085 33059 21143 33065
rect 21634 33056 21640 33108
rect 21692 33096 21698 33108
rect 21913 33099 21971 33105
rect 21913 33096 21925 33099
rect 21692 33068 21925 33096
rect 21692 33056 21698 33068
rect 21913 33065 21925 33068
rect 21959 33065 21971 33099
rect 29362 33096 29368 33108
rect 21913 33059 21971 33065
rect 22066 33068 29368 33096
rect 15746 33028 15752 33040
rect 15659 33000 15752 33028
rect 15746 32988 15752 33000
rect 15804 33028 15810 33040
rect 16298 33028 16304 33040
rect 15804 33000 16304 33028
rect 15804 32988 15810 33000
rect 16298 32988 16304 33000
rect 16356 32988 16362 33040
rect 16390 32988 16396 33040
rect 16448 33028 16454 33040
rect 19613 33031 19671 33037
rect 19613 33028 19625 33031
rect 16448 33000 17540 33028
rect 16448 32988 16454 33000
rect 14921 32963 14979 32969
rect 14921 32929 14933 32963
rect 14967 32960 14979 32963
rect 15473 32963 15531 32969
rect 15473 32960 15485 32963
rect 14967 32932 15485 32960
rect 14967 32929 14979 32932
rect 14921 32923 14979 32929
rect 15473 32929 15485 32932
rect 15519 32929 15531 32963
rect 15473 32923 15531 32929
rect 17221 32963 17279 32969
rect 17221 32929 17233 32963
rect 17267 32929 17279 32963
rect 17221 32923 17279 32929
rect 14645 32895 14703 32901
rect 14645 32892 14657 32895
rect 14516 32864 14657 32892
rect 14516 32852 14522 32864
rect 14645 32861 14657 32864
rect 14691 32861 14703 32895
rect 14645 32855 14703 32861
rect 14737 32895 14795 32901
rect 14737 32861 14749 32895
rect 14783 32892 14795 32895
rect 15102 32892 15108 32904
rect 14783 32864 15108 32892
rect 14783 32861 14795 32864
rect 14737 32855 14795 32861
rect 15102 32852 15108 32864
rect 15160 32892 15166 32904
rect 15381 32895 15439 32901
rect 15381 32892 15393 32895
rect 15160 32864 15393 32892
rect 15160 32852 15166 32864
rect 15381 32861 15393 32864
rect 15427 32861 15439 32895
rect 17129 32895 17187 32901
rect 17129 32892 17141 32895
rect 15381 32855 15439 32861
rect 16224 32864 17141 32892
rect 16114 32784 16120 32836
rect 16172 32824 16178 32836
rect 16224 32833 16252 32864
rect 17129 32861 17141 32864
rect 17175 32861 17187 32895
rect 17129 32855 17187 32861
rect 16209 32827 16267 32833
rect 16209 32824 16221 32827
rect 16172 32796 16221 32824
rect 16172 32784 16178 32796
rect 16209 32793 16221 32796
rect 16255 32793 16267 32827
rect 16390 32824 16396 32836
rect 16351 32796 16396 32824
rect 16209 32787 16267 32793
rect 16390 32784 16396 32796
rect 16448 32824 16454 32836
rect 17236 32824 17264 32923
rect 17402 32892 17408 32904
rect 17363 32864 17408 32892
rect 17402 32852 17408 32864
rect 17460 32852 17466 32904
rect 17512 32892 17540 33000
rect 18248 33000 19625 33028
rect 18248 32969 18276 33000
rect 19613 32997 19625 33000
rect 19659 33028 19671 33031
rect 22066 33028 22094 33068
rect 29362 33056 29368 33068
rect 29420 33056 29426 33108
rect 30116 33068 31340 33096
rect 19659 33000 22094 33028
rect 19659 32997 19671 33000
rect 19613 32991 19671 32997
rect 22738 32988 22744 33040
rect 22796 33028 22802 33040
rect 23198 33028 23204 33040
rect 22796 33000 23204 33028
rect 22796 32988 22802 33000
rect 23198 32988 23204 33000
rect 23256 32988 23262 33040
rect 24854 33028 24860 33040
rect 24815 33000 24860 33028
rect 24854 32988 24860 33000
rect 24912 32988 24918 33040
rect 27154 33028 27160 33040
rect 27115 33000 27160 33028
rect 27154 32988 27160 33000
rect 27212 32988 27218 33040
rect 29914 32988 29920 33040
rect 29972 33028 29978 33040
rect 30009 33031 30067 33037
rect 30009 33028 30021 33031
rect 29972 33000 30021 33028
rect 29972 32988 29978 33000
rect 30009 32997 30021 33000
rect 30055 32997 30067 33031
rect 30009 32991 30067 32997
rect 18233 32963 18291 32969
rect 18233 32929 18245 32963
rect 18279 32929 18291 32963
rect 18233 32923 18291 32929
rect 25409 32963 25467 32969
rect 25409 32929 25421 32963
rect 25455 32960 25467 32963
rect 26970 32960 26976 32972
rect 25455 32932 26976 32960
rect 25455 32929 25467 32932
rect 25409 32923 25467 32929
rect 26970 32920 26976 32932
rect 27028 32960 27034 32972
rect 27430 32960 27436 32972
rect 27028 32932 27436 32960
rect 27028 32920 27034 32932
rect 27430 32920 27436 32932
rect 27488 32920 27494 32972
rect 29546 32920 29552 32972
rect 29604 32960 29610 32972
rect 30116 32960 30144 33068
rect 30282 32988 30288 33040
rect 30340 33028 30346 33040
rect 31205 33031 31263 33037
rect 31205 33028 31217 33031
rect 30340 33000 31217 33028
rect 30340 32988 30346 33000
rect 31205 32997 31217 33000
rect 31251 32997 31263 33031
rect 31312 33028 31340 33068
rect 31662 33056 31668 33108
rect 31720 33096 31726 33108
rect 31720 33068 35894 33096
rect 31720 33056 31726 33068
rect 32401 33031 32459 33037
rect 32401 33028 32413 33031
rect 31312 33000 32413 33028
rect 31205 32991 31263 32997
rect 32401 32997 32413 33000
rect 32447 32997 32459 33031
rect 35866 33028 35894 33068
rect 48038 33028 48044 33040
rect 35866 33000 48044 33028
rect 32401 32991 32459 32997
rect 48038 32988 48044 33000
rect 48096 32988 48102 33040
rect 30374 32960 30380 32972
rect 29604 32932 30144 32960
rect 30335 32932 30380 32960
rect 29604 32920 29610 32932
rect 18325 32895 18383 32901
rect 18325 32892 18337 32895
rect 17512 32864 18337 32892
rect 18325 32861 18337 32864
rect 18371 32861 18383 32895
rect 19242 32892 19248 32904
rect 19203 32864 19248 32892
rect 18325 32855 18383 32861
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 20993 32895 21051 32901
rect 20993 32861 21005 32895
rect 21039 32892 21051 32895
rect 21082 32892 21088 32904
rect 21039 32864 21088 32892
rect 21039 32861 21051 32864
rect 20993 32855 21051 32861
rect 21082 32852 21088 32864
rect 21140 32852 21146 32904
rect 23109 32895 23167 32901
rect 23109 32861 23121 32895
rect 23155 32892 23167 32895
rect 24394 32892 24400 32904
rect 23155 32864 24400 32892
rect 23155 32861 23167 32864
rect 23109 32855 23167 32861
rect 24394 32852 24400 32864
rect 24452 32852 24458 32904
rect 24762 32892 24768 32904
rect 24723 32864 24768 32892
rect 24762 32852 24768 32864
rect 24820 32852 24826 32904
rect 27338 32852 27344 32904
rect 27396 32892 27402 32904
rect 28166 32892 28172 32904
rect 27396 32864 28028 32892
rect 28127 32864 28172 32892
rect 27396 32852 27402 32864
rect 16448 32796 17264 32824
rect 18049 32827 18107 32833
rect 16448 32784 16454 32796
rect 18049 32793 18061 32827
rect 18095 32793 18107 32827
rect 18049 32787 18107 32793
rect 2406 32716 2412 32768
rect 2464 32756 2470 32768
rect 2777 32759 2835 32765
rect 2777 32756 2789 32759
rect 2464 32728 2789 32756
rect 2464 32716 2470 32728
rect 2777 32725 2789 32728
rect 2823 32725 2835 32759
rect 2777 32719 2835 32725
rect 15838 32716 15844 32768
rect 15896 32756 15902 32768
rect 16577 32759 16635 32765
rect 16577 32756 16589 32759
rect 15896 32728 16589 32756
rect 15896 32716 15902 32728
rect 16577 32725 16589 32728
rect 16623 32725 16635 32759
rect 16577 32719 16635 32725
rect 17589 32759 17647 32765
rect 17589 32725 17601 32759
rect 17635 32756 17647 32759
rect 18064 32756 18092 32787
rect 19058 32784 19064 32836
rect 19116 32824 19122 32836
rect 19429 32827 19487 32833
rect 19429 32824 19441 32827
rect 19116 32796 19441 32824
rect 19116 32784 19122 32796
rect 19429 32793 19441 32796
rect 19475 32793 19487 32827
rect 21821 32827 21879 32833
rect 19429 32787 19487 32793
rect 19536 32796 20300 32824
rect 17635 32728 18092 32756
rect 18509 32759 18567 32765
rect 17635 32725 17647 32728
rect 17589 32719 17647 32725
rect 18509 32725 18521 32759
rect 18555 32756 18567 32759
rect 19536 32756 19564 32796
rect 18555 32728 19564 32756
rect 20272 32756 20300 32796
rect 21821 32793 21833 32827
rect 21867 32824 21879 32827
rect 25590 32824 25596 32836
rect 21867 32796 25596 32824
rect 21867 32793 21879 32796
rect 21821 32787 21879 32793
rect 25590 32784 25596 32796
rect 25648 32784 25654 32836
rect 25682 32784 25688 32836
rect 25740 32824 25746 32836
rect 27430 32824 27436 32836
rect 25740 32796 25785 32824
rect 26910 32796 27436 32824
rect 25740 32784 25746 32796
rect 27430 32784 27436 32796
rect 27488 32784 27494 32836
rect 28000 32824 28028 32864
rect 28166 32852 28172 32864
rect 28224 32852 28230 32904
rect 29932 32901 29960 32932
rect 30374 32920 30380 32932
rect 30432 32920 30438 32972
rect 32214 32960 32220 32972
rect 31128 32932 32220 32960
rect 29917 32895 29975 32901
rect 29917 32861 29929 32895
rect 29963 32861 29975 32895
rect 30190 32892 30196 32904
rect 30151 32864 30196 32892
rect 29917 32855 29975 32861
rect 30190 32852 30196 32864
rect 30248 32852 30254 32904
rect 31128 32901 31156 32932
rect 32214 32920 32220 32932
rect 32272 32920 32278 32972
rect 31113 32895 31171 32901
rect 31113 32861 31125 32895
rect 31159 32861 31171 32895
rect 31386 32892 31392 32904
rect 31347 32864 31392 32892
rect 31113 32855 31171 32861
rect 31386 32852 31392 32864
rect 31444 32852 31450 32904
rect 31478 32852 31484 32904
rect 31536 32892 31542 32904
rect 32033 32895 32091 32901
rect 31536 32864 31581 32892
rect 31536 32852 31542 32864
rect 32033 32861 32045 32895
rect 32079 32892 32091 32895
rect 32582 32892 32588 32904
rect 32079 32864 32588 32892
rect 32079 32861 32091 32864
rect 32033 32855 32091 32861
rect 32582 32852 32588 32864
rect 32640 32852 32646 32904
rect 45833 32895 45891 32901
rect 45833 32861 45845 32895
rect 45879 32892 45891 32895
rect 46293 32895 46351 32901
rect 46293 32892 46305 32895
rect 45879 32864 46305 32892
rect 45879 32861 45891 32864
rect 45833 32855 45891 32861
rect 46293 32861 46305 32864
rect 46339 32861 46351 32895
rect 46293 32855 46351 32861
rect 31662 32824 31668 32836
rect 28000 32796 31668 32824
rect 31662 32784 31668 32796
rect 31720 32784 31726 32836
rect 32217 32827 32275 32833
rect 32217 32793 32229 32827
rect 32263 32824 32275 32827
rect 32306 32824 32312 32836
rect 32263 32796 32312 32824
rect 32263 32793 32275 32796
rect 32217 32787 32275 32793
rect 32306 32784 32312 32796
rect 32364 32824 32370 32836
rect 32766 32824 32772 32836
rect 32364 32796 32772 32824
rect 32364 32784 32370 32796
rect 32766 32784 32772 32796
rect 32824 32784 32830 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 46934 32824 46940 32836
rect 46523 32796 46940 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 46934 32784 46940 32796
rect 46992 32784 46998 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 22094 32756 22100 32768
rect 20272 32728 22100 32756
rect 18555 32725 18567 32728
rect 18509 32719 18567 32725
rect 22094 32716 22100 32728
rect 22152 32716 22158 32768
rect 22370 32716 22376 32768
rect 22428 32756 22434 32768
rect 22925 32759 22983 32765
rect 22925 32756 22937 32759
rect 22428 32728 22937 32756
rect 22428 32716 22434 32728
rect 22925 32725 22937 32728
rect 22971 32725 22983 32759
rect 22925 32719 22983 32725
rect 23198 32716 23204 32768
rect 23256 32756 23262 32768
rect 27890 32756 27896 32768
rect 23256 32728 27896 32756
rect 23256 32716 23262 32728
rect 27890 32716 27896 32728
rect 27948 32716 27954 32768
rect 28258 32756 28264 32768
rect 28219 32728 28264 32756
rect 28258 32716 28264 32728
rect 28316 32716 28322 32768
rect 28994 32716 29000 32768
rect 29052 32756 29058 32768
rect 29454 32756 29460 32768
rect 29052 32728 29460 32756
rect 29052 32716 29058 32728
rect 29454 32716 29460 32728
rect 29512 32716 29518 32768
rect 30374 32716 30380 32768
rect 30432 32756 30438 32768
rect 31478 32756 31484 32768
rect 30432 32728 31484 32756
rect 30432 32716 30438 32728
rect 31478 32716 31484 32728
rect 31536 32716 31542 32768
rect 31573 32759 31631 32765
rect 31573 32725 31585 32759
rect 31619 32756 31631 32759
rect 31754 32756 31760 32768
rect 31619 32728 31760 32756
rect 31619 32725 31631 32728
rect 31573 32719 31631 32725
rect 31754 32716 31760 32728
rect 31812 32716 31818 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 17402 32512 17408 32564
rect 17460 32552 17466 32564
rect 23382 32552 23388 32564
rect 17460 32524 23388 32552
rect 17460 32512 17466 32524
rect 23382 32512 23388 32524
rect 23440 32552 23446 32564
rect 23845 32555 23903 32561
rect 23845 32552 23857 32555
rect 23440 32524 23857 32552
rect 23440 32512 23446 32524
rect 23845 32521 23857 32524
rect 23891 32521 23903 32555
rect 25590 32552 25596 32564
rect 25551 32524 25596 32552
rect 23845 32515 23903 32521
rect 25590 32512 25596 32524
rect 25648 32512 25654 32564
rect 26142 32512 26148 32564
rect 26200 32552 26206 32564
rect 28353 32555 28411 32561
rect 28353 32552 28365 32555
rect 26200 32524 28365 32552
rect 26200 32512 26206 32524
rect 28353 32521 28365 32524
rect 28399 32521 28411 32555
rect 28353 32515 28411 32521
rect 29641 32555 29699 32561
rect 29641 32521 29653 32555
rect 29687 32552 29699 32555
rect 29914 32552 29920 32564
rect 29687 32524 29920 32552
rect 29687 32521 29699 32524
rect 29641 32515 29699 32521
rect 29914 32512 29920 32524
rect 29972 32512 29978 32564
rect 44174 32552 44180 32564
rect 31726 32524 44180 32552
rect 2406 32484 2412 32496
rect 2367 32456 2412 32484
rect 2406 32444 2412 32456
rect 2464 32444 2470 32496
rect 14734 32444 14740 32496
rect 14792 32484 14798 32496
rect 15102 32484 15108 32496
rect 14792 32456 15108 32484
rect 14792 32444 14798 32456
rect 15102 32444 15108 32456
rect 15160 32484 15166 32496
rect 15657 32487 15715 32493
rect 15657 32484 15669 32487
rect 15160 32456 15669 32484
rect 15160 32444 15166 32456
rect 15657 32453 15669 32456
rect 15703 32484 15715 32487
rect 17862 32484 17868 32496
rect 15703 32456 17868 32484
rect 15703 32453 15715 32456
rect 15657 32447 15715 32453
rect 17862 32444 17868 32456
rect 17920 32444 17926 32496
rect 20070 32444 20076 32496
rect 20128 32484 20134 32496
rect 20622 32484 20628 32496
rect 20128 32456 20628 32484
rect 20128 32444 20134 32456
rect 20622 32444 20628 32456
rect 20680 32484 20686 32496
rect 22370 32484 22376 32496
rect 20680 32456 22140 32484
rect 22331 32456 22376 32484
rect 20680 32444 20686 32456
rect 2222 32416 2228 32428
rect 2183 32388 2228 32416
rect 2222 32376 2228 32388
rect 2280 32376 2286 32428
rect 15838 32416 15844 32428
rect 15799 32388 15844 32416
rect 15838 32376 15844 32388
rect 15896 32376 15902 32428
rect 15930 32376 15936 32428
rect 15988 32416 15994 32428
rect 17218 32416 17224 32428
rect 15988 32388 16033 32416
rect 16132 32388 17224 32416
rect 15988 32376 15994 32388
rect 4065 32351 4123 32357
rect 4065 32317 4077 32351
rect 4111 32348 4123 32351
rect 4614 32348 4620 32360
rect 4111 32320 4620 32348
rect 4111 32317 4123 32320
rect 4065 32311 4123 32317
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 16132 32289 16160 32388
rect 17218 32376 17224 32388
rect 17276 32376 17282 32428
rect 22112 32425 22140 32456
rect 22370 32444 22376 32456
rect 22428 32444 22434 32496
rect 22646 32444 22652 32496
rect 22704 32484 22710 32496
rect 22704 32456 22862 32484
rect 22704 32444 22710 32456
rect 24762 32444 24768 32496
rect 24820 32484 24826 32496
rect 28261 32487 28319 32493
rect 28261 32484 28273 32487
rect 24820 32456 28273 32484
rect 24820 32444 24826 32456
rect 28261 32453 28273 32456
rect 28307 32484 28319 32487
rect 31726 32484 31754 32524
rect 44174 32512 44180 32524
rect 44232 32512 44238 32564
rect 46934 32552 46940 32564
rect 46895 32524 46940 32552
rect 46934 32512 46940 32524
rect 46992 32512 46998 32564
rect 48038 32552 48044 32564
rect 47999 32524 48044 32552
rect 48038 32512 48044 32524
rect 48096 32512 48102 32564
rect 28307 32456 31754 32484
rect 28307 32453 28319 32456
rect 28261 32447 28319 32453
rect 33042 32444 33048 32496
rect 33100 32444 33106 32496
rect 20809 32419 20867 32425
rect 20809 32385 20821 32419
rect 20855 32385 20867 32419
rect 20809 32379 20867 32385
rect 22097 32419 22155 32425
rect 22097 32385 22109 32419
rect 22143 32385 22155 32419
rect 24302 32416 24308 32428
rect 24263 32388 24308 32416
rect 22097 32379 22155 32385
rect 16206 32308 16212 32360
rect 16264 32348 16270 32360
rect 17497 32351 17555 32357
rect 17497 32348 17509 32351
rect 16264 32320 17509 32348
rect 16264 32308 16270 32320
rect 17497 32317 17509 32320
rect 17543 32317 17555 32351
rect 17497 32311 17555 32317
rect 16117 32283 16175 32289
rect 16117 32249 16129 32283
rect 16163 32249 16175 32283
rect 18230 32280 18236 32292
rect 16117 32243 16175 32249
rect 17512 32252 18236 32280
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1765 32215 1823 32221
rect 1765 32212 1777 32215
rect 1452 32184 1777 32212
rect 1452 32172 1458 32184
rect 1765 32181 1777 32184
rect 1811 32181 1823 32215
rect 1765 32175 1823 32181
rect 14458 32172 14464 32224
rect 14516 32212 14522 32224
rect 17512 32221 17540 32252
rect 18230 32240 18236 32252
rect 18288 32240 18294 32292
rect 20824 32280 20852 32379
rect 24302 32376 24308 32388
rect 24360 32376 24366 32428
rect 27341 32419 27399 32425
rect 27341 32385 27353 32419
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 27433 32419 27491 32425
rect 27433 32385 27445 32419
rect 27479 32416 27491 32419
rect 27709 32419 27767 32425
rect 27479 32388 27660 32416
rect 27479 32385 27491 32388
rect 27433 32379 27491 32385
rect 23658 32348 23664 32360
rect 22066 32320 23664 32348
rect 22066 32280 22094 32320
rect 23658 32308 23664 32320
rect 23716 32348 23722 32360
rect 24670 32348 24676 32360
rect 23716 32320 24676 32348
rect 23716 32308 23722 32320
rect 24670 32308 24676 32320
rect 24728 32308 24734 32360
rect 27356 32348 27384 32379
rect 27632 32348 27660 32388
rect 27709 32385 27721 32419
rect 27755 32416 27767 32419
rect 27798 32416 27804 32428
rect 27755 32388 27804 32416
rect 27755 32385 27767 32388
rect 27709 32379 27767 32385
rect 27798 32376 27804 32388
rect 27856 32376 27862 32428
rect 29273 32419 29331 32425
rect 29273 32385 29285 32419
rect 29319 32416 29331 32419
rect 29362 32416 29368 32428
rect 29319 32388 29368 32416
rect 29319 32385 29331 32388
rect 29273 32379 29331 32385
rect 29362 32376 29368 32388
rect 29420 32376 29426 32428
rect 29457 32419 29515 32425
rect 29457 32385 29469 32419
rect 29503 32385 29515 32419
rect 29457 32379 29515 32385
rect 27890 32348 27896 32360
rect 27356 32320 27476 32348
rect 27632 32320 27896 32348
rect 27338 32280 27344 32292
rect 20824 32252 22094 32280
rect 24136 32252 27344 32280
rect 15657 32215 15715 32221
rect 15657 32212 15669 32215
rect 14516 32184 15669 32212
rect 14516 32172 14522 32184
rect 15657 32181 15669 32184
rect 15703 32181 15715 32215
rect 15657 32175 15715 32181
rect 17497 32215 17555 32221
rect 17497 32181 17509 32215
rect 17543 32181 17555 32215
rect 17497 32175 17555 32181
rect 17586 32172 17592 32224
rect 17644 32212 17650 32224
rect 17773 32215 17831 32221
rect 17773 32212 17785 32215
rect 17644 32184 17785 32212
rect 17644 32172 17650 32184
rect 17773 32181 17785 32184
rect 17819 32181 17831 32215
rect 17773 32175 17831 32181
rect 18322 32172 18328 32224
rect 18380 32212 18386 32224
rect 20993 32215 21051 32221
rect 20993 32212 21005 32215
rect 18380 32184 21005 32212
rect 18380 32172 18386 32184
rect 20993 32181 21005 32184
rect 21039 32212 21051 32215
rect 24136 32212 24164 32252
rect 27338 32240 27344 32252
rect 27396 32240 27402 32292
rect 27448 32280 27476 32320
rect 27890 32308 27896 32320
rect 27948 32308 27954 32360
rect 28810 32308 28816 32360
rect 28868 32348 28874 32360
rect 29472 32348 29500 32379
rect 30006 32376 30012 32428
rect 30064 32416 30070 32428
rect 30377 32419 30435 32425
rect 30377 32416 30389 32419
rect 30064 32388 30389 32416
rect 30064 32376 30070 32388
rect 30377 32385 30389 32388
rect 30423 32385 30435 32419
rect 32122 32416 32128 32428
rect 32083 32388 32128 32416
rect 30377 32379 30435 32385
rect 32122 32376 32128 32388
rect 32180 32376 32186 32428
rect 45554 32376 45560 32428
rect 45612 32416 45618 32428
rect 46845 32419 46903 32425
rect 46845 32416 46857 32419
rect 45612 32388 46857 32416
rect 45612 32376 45618 32388
rect 46845 32385 46857 32388
rect 46891 32385 46903 32419
rect 47946 32416 47952 32428
rect 47907 32388 47952 32416
rect 46845 32379 46903 32385
rect 47946 32376 47952 32388
rect 48004 32376 48010 32428
rect 28868 32320 29500 32348
rect 28868 32308 28874 32320
rect 28902 32280 28908 32292
rect 27448 32252 28908 32280
rect 28902 32240 28908 32252
rect 28960 32240 28966 32292
rect 29472 32280 29500 32320
rect 30101 32351 30159 32357
rect 30101 32317 30113 32351
rect 30147 32348 30159 32351
rect 30190 32348 30196 32360
rect 30147 32320 30196 32348
rect 30147 32317 30159 32320
rect 30101 32311 30159 32317
rect 30190 32308 30196 32320
rect 30248 32308 30254 32360
rect 32401 32351 32459 32357
rect 32401 32317 32413 32351
rect 32447 32348 32459 32351
rect 32490 32348 32496 32360
rect 32447 32320 32496 32348
rect 32447 32317 32459 32320
rect 32401 32311 32459 32317
rect 32490 32308 32496 32320
rect 32548 32308 32554 32360
rect 32766 32308 32772 32360
rect 32824 32348 32830 32360
rect 33873 32351 33931 32357
rect 33873 32348 33885 32351
rect 32824 32320 33885 32348
rect 32824 32308 32830 32320
rect 33873 32317 33885 32320
rect 33919 32317 33931 32351
rect 33873 32311 33931 32317
rect 30926 32280 30932 32292
rect 29472 32252 30932 32280
rect 30926 32240 30932 32252
rect 30984 32240 30990 32292
rect 21039 32184 24164 32212
rect 27157 32215 27215 32221
rect 21039 32181 21051 32184
rect 20993 32175 21051 32181
rect 27157 32181 27169 32215
rect 27203 32212 27215 32215
rect 27246 32212 27252 32224
rect 27203 32184 27252 32212
rect 27203 32181 27215 32184
rect 27157 32175 27215 32181
rect 27246 32172 27252 32184
rect 27304 32172 27310 32224
rect 27617 32215 27675 32221
rect 27617 32181 27629 32215
rect 27663 32212 27675 32215
rect 27706 32212 27712 32224
rect 27663 32184 27712 32212
rect 27663 32181 27675 32184
rect 27617 32175 27675 32181
rect 27706 32172 27712 32184
rect 27764 32172 27770 32224
rect 28994 32172 29000 32224
rect 29052 32212 29058 32224
rect 29178 32212 29184 32224
rect 29052 32184 29184 32212
rect 29052 32172 29058 32184
rect 29178 32172 29184 32184
rect 29236 32212 29242 32224
rect 32214 32212 32220 32224
rect 29236 32184 32220 32212
rect 29236 32172 29242 32184
rect 32214 32172 32220 32184
rect 32272 32172 32278 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 16206 32008 16212 32020
rect 16167 31980 16212 32008
rect 16206 31968 16212 31980
rect 16264 31968 16270 32020
rect 16298 31968 16304 32020
rect 16356 32008 16362 32020
rect 16577 32011 16635 32017
rect 16577 32008 16589 32011
rect 16356 31980 16589 32008
rect 16356 31968 16362 31980
rect 16577 31977 16589 31980
rect 16623 31977 16635 32011
rect 16577 31971 16635 31977
rect 19242 31968 19248 32020
rect 19300 32008 19306 32020
rect 22646 32008 22652 32020
rect 19300 31980 22508 32008
rect 22607 31980 22652 32008
rect 19300 31968 19306 31980
rect 16390 31940 16396 31952
rect 16303 31912 16396 31940
rect 16390 31900 16396 31912
rect 16448 31940 16454 31952
rect 16448 31912 17908 31940
rect 16448 31900 16454 31912
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 1946 31832 1952 31884
rect 2004 31872 2010 31884
rect 3973 31875 4031 31881
rect 3973 31872 3985 31875
rect 2004 31844 3985 31872
rect 2004 31832 2010 31844
rect 3973 31841 3985 31844
rect 4019 31841 4031 31875
rect 4614 31872 4620 31884
rect 4575 31844 4620 31872
rect 3973 31835 4031 31841
rect 4614 31832 4620 31844
rect 4672 31872 4678 31884
rect 5442 31872 5448 31884
rect 4672 31844 5448 31872
rect 4672 31832 4678 31844
rect 5442 31832 5448 31844
rect 5500 31832 5506 31884
rect 16114 31832 16120 31884
rect 16172 31872 16178 31884
rect 16172 31844 16344 31872
rect 16172 31832 16178 31844
rect 3786 31804 3792 31816
rect 3747 31776 3792 31804
rect 3786 31764 3792 31776
rect 3844 31764 3850 31816
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 16316 31736 16344 31844
rect 16408 31813 16436 31900
rect 17880 31881 17908 31912
rect 16669 31875 16727 31881
rect 16669 31872 16681 31875
rect 16500 31844 16681 31872
rect 16393 31807 16451 31813
rect 16393 31773 16405 31807
rect 16439 31773 16451 31807
rect 16393 31767 16451 31773
rect 16500 31736 16528 31844
rect 16669 31841 16681 31844
rect 16715 31841 16727 31875
rect 16669 31835 16727 31841
rect 17865 31875 17923 31881
rect 17865 31841 17877 31875
rect 17911 31872 17923 31875
rect 19334 31872 19340 31884
rect 17911 31844 19340 31872
rect 17911 31841 17923 31844
rect 17865 31835 17923 31841
rect 19334 31832 19340 31844
rect 19392 31832 19398 31884
rect 20070 31872 20076 31884
rect 20031 31844 20076 31872
rect 20070 31832 20076 31844
rect 20128 31832 20134 31884
rect 20349 31875 20407 31881
rect 20349 31841 20361 31875
rect 20395 31872 20407 31875
rect 21082 31872 21088 31884
rect 20395 31844 21088 31872
rect 20395 31841 20407 31844
rect 20349 31835 20407 31841
rect 21082 31832 21088 31844
rect 21140 31832 21146 31884
rect 22480 31872 22508 31980
rect 22646 31968 22652 31980
rect 22704 31968 22710 32020
rect 24394 32008 24400 32020
rect 24355 31980 24400 32008
rect 24394 31968 24400 31980
rect 24452 31968 24458 32020
rect 25593 32011 25651 32017
rect 25593 31977 25605 32011
rect 25639 32008 25651 32011
rect 26326 32008 26332 32020
rect 25639 31980 26332 32008
rect 25639 31977 25651 31980
rect 25593 31971 25651 31977
rect 26326 31968 26332 31980
rect 26384 31968 26390 32020
rect 26436 31980 28994 32008
rect 26436 31940 26464 31980
rect 25700 31912 26464 31940
rect 28721 31943 28779 31949
rect 23474 31872 23480 31884
rect 22480 31844 22600 31872
rect 23435 31844 23480 31872
rect 17586 31804 17592 31816
rect 17547 31776 17592 31804
rect 17586 31764 17592 31776
rect 17644 31764 17650 31816
rect 17773 31807 17831 31813
rect 17773 31773 17785 31807
rect 17819 31804 17831 31807
rect 17957 31807 18015 31813
rect 17819 31776 17908 31804
rect 17819 31773 17831 31776
rect 17773 31767 17831 31773
rect 16316 31708 16528 31736
rect 17880 31736 17908 31776
rect 17957 31773 17969 31807
rect 18003 31804 18015 31807
rect 18141 31807 18199 31813
rect 18003 31776 18092 31804
rect 18003 31773 18015 31776
rect 17957 31767 18015 31773
rect 17880 31708 18000 31736
rect 17972 31680 18000 31708
rect 16942 31628 16948 31680
rect 17000 31668 17006 31680
rect 17126 31668 17132 31680
rect 17000 31640 17132 31668
rect 17000 31628 17006 31640
rect 17126 31628 17132 31640
rect 17184 31628 17190 31680
rect 17954 31628 17960 31680
rect 18012 31628 18018 31680
rect 18064 31668 18092 31776
rect 18141 31773 18153 31807
rect 18187 31804 18199 31807
rect 18322 31804 18328 31816
rect 18187 31776 18328 31804
rect 18187 31773 18199 31776
rect 18141 31767 18199 31773
rect 18322 31764 18328 31776
rect 18380 31764 18386 31816
rect 22462 31804 22468 31816
rect 21482 31776 22468 31804
rect 22462 31764 22468 31776
rect 22520 31764 22526 31816
rect 22572 31813 22600 31844
rect 23474 31832 23480 31844
rect 23532 31832 23538 31884
rect 23753 31875 23811 31881
rect 23753 31841 23765 31875
rect 23799 31872 23811 31875
rect 24857 31875 24915 31881
rect 24857 31872 24869 31875
rect 23799 31844 24869 31872
rect 23799 31841 23811 31844
rect 23753 31835 23811 31841
rect 24857 31841 24869 31844
rect 24903 31841 24915 31875
rect 25038 31872 25044 31884
rect 24999 31844 25044 31872
rect 24857 31835 24915 31841
rect 25038 31832 25044 31844
rect 25096 31832 25102 31884
rect 22557 31807 22615 31813
rect 22557 31773 22569 31807
rect 22603 31773 22615 31807
rect 23382 31804 23388 31816
rect 23343 31776 23388 31804
rect 22557 31767 22615 31773
rect 22572 31736 22600 31767
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31804 24823 31807
rect 25501 31807 25559 31813
rect 25501 31804 25513 31807
rect 24811 31776 25513 31804
rect 24811 31773 24823 31776
rect 24765 31767 24823 31773
rect 25501 31773 25513 31776
rect 25547 31804 25559 31807
rect 25700 31804 25728 31912
rect 28721 31909 28733 31943
rect 28767 31940 28779 31943
rect 28810 31940 28816 31952
rect 28767 31912 28816 31940
rect 28767 31909 28779 31912
rect 28721 31903 28779 31909
rect 28810 31900 28816 31912
rect 28868 31900 28874 31952
rect 28966 31940 28994 31980
rect 29822 31968 29828 32020
rect 29880 32008 29886 32020
rect 29917 32011 29975 32017
rect 29917 32008 29929 32011
rect 29880 31980 29929 32008
rect 29880 31968 29886 31980
rect 29917 31977 29929 31980
rect 29963 31977 29975 32011
rect 29917 31971 29975 31977
rect 30282 31968 30288 32020
rect 30340 32008 30346 32020
rect 30745 32011 30803 32017
rect 30745 32008 30757 32011
rect 30340 31980 30757 32008
rect 30340 31968 30346 31980
rect 30745 31977 30757 31980
rect 30791 31977 30803 32011
rect 32490 32008 32496 32020
rect 32451 31980 32496 32008
rect 30745 31971 30803 31977
rect 32490 31968 32496 31980
rect 32548 31968 32554 32020
rect 33042 32008 33048 32020
rect 33003 31980 33048 32008
rect 33042 31968 33048 31980
rect 33100 31968 33106 32020
rect 48222 32008 48228 32020
rect 38626 31980 48228 32008
rect 38626 31940 38654 31980
rect 48222 31968 48228 31980
rect 48280 31968 48286 32020
rect 28966 31912 38654 31940
rect 42702 31900 42708 31952
rect 42760 31940 42766 31952
rect 42760 31912 47440 31940
rect 42760 31900 42766 31912
rect 47412 31884 47440 31912
rect 26970 31872 26976 31884
rect 26931 31844 26976 31872
rect 26970 31832 26976 31844
rect 27028 31832 27034 31884
rect 27246 31872 27252 31884
rect 27207 31844 27252 31872
rect 27246 31832 27252 31844
rect 27304 31832 27310 31884
rect 27338 31832 27344 31884
rect 27396 31872 27402 31884
rect 28994 31872 29000 31884
rect 27396 31844 29000 31872
rect 27396 31832 27402 31844
rect 28994 31832 29000 31844
rect 29052 31832 29058 31884
rect 32033 31875 32091 31881
rect 29840 31844 31984 31872
rect 25547 31776 25728 31804
rect 25777 31807 25835 31813
rect 25547 31773 25559 31776
rect 25501 31767 25559 31773
rect 25777 31773 25789 31807
rect 25823 31804 25835 31807
rect 25958 31804 25964 31816
rect 25823 31776 25964 31804
rect 25823 31773 25835 31776
rect 25777 31767 25835 31773
rect 25958 31764 25964 31776
rect 26016 31764 26022 31816
rect 26053 31807 26111 31813
rect 26053 31773 26065 31807
rect 26099 31804 26111 31807
rect 26099 31776 26133 31804
rect 26099 31773 26111 31776
rect 26053 31767 26111 31773
rect 25682 31736 25688 31748
rect 22572 31708 25688 31736
rect 25682 31696 25688 31708
rect 25740 31696 25746 31748
rect 26068 31736 26096 31767
rect 28258 31764 28264 31816
rect 28316 31804 28322 31816
rect 28316 31776 28382 31804
rect 28316 31764 28322 31776
rect 28626 31764 28632 31816
rect 28684 31804 28690 31816
rect 29840 31804 29868 31844
rect 31956 31816 31984 31844
rect 32033 31841 32045 31875
rect 32079 31872 32091 31875
rect 32766 31872 32772 31884
rect 32079 31844 32772 31872
rect 32079 31841 32091 31844
rect 32033 31835 32091 31841
rect 32766 31832 32772 31844
rect 32824 31832 32830 31884
rect 46569 31875 46627 31881
rect 46569 31841 46581 31875
rect 46615 31872 46627 31875
rect 46750 31872 46756 31884
rect 46615 31844 46756 31872
rect 46615 31841 46627 31844
rect 46569 31835 46627 31841
rect 46750 31832 46756 31844
rect 46808 31832 46814 31884
rect 47394 31872 47400 31884
rect 47355 31844 47400 31872
rect 47394 31832 47400 31844
rect 47452 31832 47458 31884
rect 28684 31776 29868 31804
rect 29917 31807 29975 31813
rect 28684 31764 28690 31776
rect 29917 31773 29929 31807
rect 29963 31804 29975 31807
rect 30006 31804 30012 31816
rect 29963 31776 30012 31804
rect 29963 31773 29975 31776
rect 29917 31767 29975 31773
rect 30006 31764 30012 31776
rect 30064 31764 30070 31816
rect 30098 31764 30104 31816
rect 30156 31804 30162 31816
rect 30745 31807 30803 31813
rect 30745 31804 30757 31807
rect 30156 31776 30201 31804
rect 30300 31776 30757 31804
rect 30156 31764 30162 31776
rect 25884 31708 26096 31736
rect 18138 31668 18144 31680
rect 18064 31640 18144 31668
rect 18138 31628 18144 31640
rect 18196 31628 18202 31680
rect 18322 31668 18328 31680
rect 18283 31640 18328 31668
rect 18322 31628 18328 31640
rect 18380 31628 18386 31680
rect 21821 31671 21879 31677
rect 21821 31637 21833 31671
rect 21867 31668 21879 31671
rect 22002 31668 22008 31680
rect 21867 31640 22008 31668
rect 21867 31637 21879 31640
rect 21821 31631 21879 31637
rect 22002 31628 22008 31640
rect 22060 31628 22066 31680
rect 25222 31628 25228 31680
rect 25280 31668 25286 31680
rect 25884 31668 25912 31708
rect 29362 31696 29368 31748
rect 29420 31736 29426 31748
rect 30116 31736 30144 31764
rect 29420 31708 30144 31736
rect 29420 31696 29426 31708
rect 25280 31640 25912 31668
rect 25961 31671 26019 31677
rect 25280 31628 25286 31640
rect 25961 31637 25973 31671
rect 26007 31668 26019 31671
rect 26142 31668 26148 31680
rect 26007 31640 26148 31668
rect 26007 31637 26019 31640
rect 25961 31631 26019 31637
rect 26142 31628 26148 31640
rect 26200 31628 26206 31680
rect 28994 31628 29000 31680
rect 29052 31668 29058 31680
rect 30300 31677 30328 31776
rect 30745 31773 30757 31776
rect 30791 31773 30803 31807
rect 30926 31804 30932 31816
rect 30887 31776 30932 31804
rect 30745 31767 30803 31773
rect 30926 31764 30932 31776
rect 30984 31764 30990 31816
rect 31754 31804 31760 31816
rect 31715 31776 31760 31804
rect 31754 31764 31760 31776
rect 31812 31764 31818 31816
rect 31938 31764 31944 31816
rect 31996 31804 32002 31816
rect 31996 31776 32089 31804
rect 31996 31764 32002 31776
rect 32122 31764 32128 31816
rect 32180 31804 32186 31816
rect 32180 31776 32225 31804
rect 32180 31764 32186 31776
rect 32306 31764 32312 31816
rect 32364 31804 32370 31816
rect 32364 31776 32409 31804
rect 32364 31764 32370 31776
rect 32858 31764 32864 31816
rect 32916 31804 32922 31816
rect 32953 31807 33011 31813
rect 32953 31804 32965 31807
rect 32916 31776 32965 31804
rect 32916 31764 32922 31776
rect 32953 31773 32965 31776
rect 32999 31773 33011 31807
rect 32953 31767 33011 31773
rect 46658 31736 46664 31748
rect 46619 31708 46664 31736
rect 46658 31696 46664 31708
rect 46716 31696 46722 31748
rect 30285 31671 30343 31677
rect 30285 31668 30297 31671
rect 29052 31640 30297 31668
rect 29052 31628 29058 31640
rect 30285 31637 30297 31640
rect 30331 31637 30343 31671
rect 30285 31631 30343 31637
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 2225 31467 2283 31473
rect 2225 31464 2237 31467
rect 1636 31436 2237 31464
rect 1636 31424 1642 31436
rect 2225 31433 2237 31436
rect 2271 31433 2283 31467
rect 17310 31464 17316 31476
rect 2225 31427 2283 31433
rect 17144 31436 17316 31464
rect 17144 31340 17172 31436
rect 17310 31424 17316 31436
rect 17368 31424 17374 31476
rect 19334 31424 19340 31476
rect 19392 31464 19398 31476
rect 19521 31467 19579 31473
rect 19521 31464 19533 31467
rect 19392 31436 19533 31464
rect 19392 31424 19398 31436
rect 19521 31433 19533 31436
rect 19567 31433 19579 31467
rect 19521 31427 19579 31433
rect 21082 31424 21088 31476
rect 21140 31464 21146 31476
rect 21269 31467 21327 31473
rect 21269 31464 21281 31467
rect 21140 31436 21281 31464
rect 21140 31424 21146 31436
rect 21269 31433 21281 31436
rect 21315 31433 21327 31467
rect 21269 31427 21327 31433
rect 22462 31424 22468 31476
rect 22520 31464 22526 31476
rect 22649 31467 22707 31473
rect 22649 31464 22661 31467
rect 22520 31436 22661 31464
rect 22520 31424 22526 31436
rect 22649 31433 22661 31436
rect 22695 31433 22707 31467
rect 23585 31467 23643 31473
rect 23585 31464 23597 31467
rect 22649 31427 22707 31433
rect 22756 31436 23597 31464
rect 18049 31399 18107 31405
rect 18049 31365 18061 31399
rect 18095 31396 18107 31399
rect 18322 31396 18328 31408
rect 18095 31368 18328 31396
rect 18095 31365 18107 31368
rect 18049 31359 18107 31365
rect 18322 31356 18328 31368
rect 18380 31356 18386 31408
rect 20346 31356 20352 31408
rect 20404 31396 20410 31408
rect 20404 31368 20760 31396
rect 20404 31356 20410 31368
rect 20732 31340 20760 31368
rect 21634 31356 21640 31408
rect 21692 31396 21698 31408
rect 21913 31399 21971 31405
rect 21913 31396 21925 31399
rect 21692 31368 21925 31396
rect 21692 31356 21698 31368
rect 21913 31365 21925 31368
rect 21959 31365 21971 31399
rect 21913 31359 21971 31365
rect 2038 31288 2044 31340
rect 2096 31328 2102 31340
rect 2133 31331 2191 31337
rect 2133 31328 2145 31331
rect 2096 31300 2145 31328
rect 2096 31288 2102 31300
rect 2133 31297 2145 31300
rect 2179 31328 2191 31331
rect 2222 31328 2228 31340
rect 2179 31300 2228 31328
rect 2179 31297 2191 31300
rect 2133 31291 2191 31297
rect 2222 31288 2228 31300
rect 2280 31288 2286 31340
rect 14458 31328 14464 31340
rect 14371 31300 14464 31328
rect 14458 31288 14464 31300
rect 14516 31288 14522 31340
rect 15289 31331 15347 31337
rect 15289 31328 15301 31331
rect 14844 31300 15301 31328
rect 14476 31192 14504 31288
rect 14553 31263 14611 31269
rect 14553 31229 14565 31263
rect 14599 31260 14611 31263
rect 14734 31260 14740 31272
rect 14599 31232 14740 31260
rect 14599 31229 14611 31232
rect 14553 31223 14611 31229
rect 14734 31220 14740 31232
rect 14792 31220 14798 31272
rect 14844 31269 14872 31300
rect 15289 31297 15301 31300
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 15473 31331 15531 31337
rect 15473 31297 15485 31331
rect 15519 31328 15531 31331
rect 16850 31328 16856 31340
rect 15519 31300 16856 31328
rect 15519 31297 15531 31300
rect 15473 31291 15531 31297
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 17126 31328 17132 31340
rect 17087 31300 17132 31328
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 19334 31328 19340 31340
rect 19182 31300 19340 31328
rect 19334 31288 19340 31300
rect 19392 31288 19398 31340
rect 20530 31328 20536 31340
rect 20491 31300 20536 31328
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 20714 31328 20720 31340
rect 20675 31300 20720 31328
rect 20714 31288 20720 31300
rect 20772 31288 20778 31340
rect 21085 31331 21143 31337
rect 21085 31297 21097 31331
rect 21131 31328 21143 31331
rect 21818 31328 21824 31340
rect 21131 31300 21824 31328
rect 21131 31297 21143 31300
rect 21085 31291 21143 31297
rect 21818 31288 21824 31300
rect 21876 31288 21882 31340
rect 22554 31328 22560 31340
rect 21928 31300 22560 31328
rect 14829 31263 14887 31269
rect 14829 31229 14841 31263
rect 14875 31229 14887 31263
rect 14829 31223 14887 31229
rect 17218 31220 17224 31272
rect 17276 31260 17282 31272
rect 17773 31263 17831 31269
rect 17773 31260 17785 31263
rect 17276 31232 17785 31260
rect 17276 31220 17282 31232
rect 17773 31229 17785 31232
rect 17819 31229 17831 31263
rect 17773 31223 17831 31229
rect 18046 31220 18052 31272
rect 18104 31260 18110 31272
rect 20806 31260 20812 31272
rect 18104 31232 19104 31260
rect 20767 31232 20812 31260
rect 18104 31220 18110 31232
rect 14918 31192 14924 31204
rect 14476 31164 14924 31192
rect 14918 31152 14924 31164
rect 14976 31192 14982 31204
rect 17313 31195 17371 31201
rect 17313 31192 17325 31195
rect 14976 31164 17325 31192
rect 14976 31152 14982 31164
rect 17313 31161 17325 31164
rect 17359 31161 17371 31195
rect 19076 31192 19104 31232
rect 20806 31220 20812 31232
rect 20864 31220 20870 31272
rect 20901 31263 20959 31269
rect 20901 31229 20913 31263
rect 20947 31260 20959 31263
rect 21542 31260 21548 31272
rect 20947 31232 21548 31260
rect 20947 31229 20959 31232
rect 20901 31223 20959 31229
rect 20916 31192 20944 31223
rect 21542 31220 21548 31232
rect 21600 31220 21606 31272
rect 19076 31164 20944 31192
rect 17313 31155 17371 31161
rect 21174 31152 21180 31204
rect 21232 31192 21238 31204
rect 21928 31192 21956 31300
rect 22554 31288 22560 31300
rect 22612 31288 22618 31340
rect 21232 31164 21956 31192
rect 21232 31152 21238 31164
rect 22094 31152 22100 31204
rect 22152 31192 22158 31204
rect 22152 31164 22197 31192
rect 22152 31152 22158 31164
rect 15286 31124 15292 31136
rect 15247 31096 15292 31124
rect 15286 31084 15292 31096
rect 15344 31084 15350 31136
rect 17862 31084 17868 31136
rect 17920 31124 17926 31136
rect 22756 31124 22784 31436
rect 23585 31433 23597 31436
rect 23631 31433 23643 31467
rect 23750 31464 23756 31476
rect 23711 31436 23756 31464
rect 23585 31427 23643 31433
rect 23750 31424 23756 31436
rect 23808 31424 23814 31476
rect 24578 31464 24584 31476
rect 24539 31436 24584 31464
rect 24578 31424 24584 31436
rect 24636 31424 24642 31476
rect 25038 31424 25044 31476
rect 25096 31464 25102 31476
rect 25225 31467 25283 31473
rect 25225 31464 25237 31467
rect 25096 31436 25237 31464
rect 25096 31424 25102 31436
rect 25225 31433 25237 31436
rect 25271 31433 25283 31467
rect 27890 31464 27896 31476
rect 27851 31436 27896 31464
rect 25225 31427 25283 31433
rect 27890 31424 27896 31436
rect 27948 31424 27954 31476
rect 28442 31464 28448 31476
rect 28092 31436 28448 31464
rect 23385 31399 23443 31405
rect 23385 31365 23397 31399
rect 23431 31365 23443 31399
rect 24210 31396 24216 31408
rect 24171 31368 24216 31396
rect 23385 31359 23443 31365
rect 23400 31328 23428 31359
rect 24210 31356 24216 31368
rect 24268 31356 24274 31408
rect 24413 31399 24471 31405
rect 24413 31396 24425 31399
rect 24412 31365 24425 31396
rect 24459 31396 24471 31399
rect 24459 31368 25268 31396
rect 24459 31365 24471 31368
rect 24412 31359 24471 31365
rect 24228 31328 24256 31356
rect 23400 31300 24256 31328
rect 24412 31260 24440 31359
rect 25240 31340 25268 31368
rect 25590 31356 25596 31408
rect 25648 31396 25654 31408
rect 27065 31399 27123 31405
rect 27065 31396 27077 31399
rect 25648 31368 27077 31396
rect 25648 31356 25654 31368
rect 27065 31365 27077 31368
rect 27111 31365 27123 31399
rect 27065 31359 27123 31365
rect 27249 31399 27307 31405
rect 27249 31365 27261 31399
rect 27295 31396 27307 31399
rect 27522 31396 27528 31408
rect 27295 31368 27528 31396
rect 27295 31365 27307 31368
rect 27249 31359 27307 31365
rect 27522 31356 27528 31368
rect 27580 31356 27586 31408
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31297 25191 31331
rect 25133 31291 25191 31297
rect 25148 31260 25176 31291
rect 25222 31288 25228 31340
rect 25280 31288 25286 31340
rect 25777 31331 25835 31337
rect 25777 31297 25789 31331
rect 25823 31328 25835 31331
rect 25958 31328 25964 31340
rect 25823 31300 25964 31328
rect 25823 31297 25835 31300
rect 25777 31291 25835 31297
rect 25958 31288 25964 31300
rect 26016 31288 26022 31340
rect 27982 31288 27988 31340
rect 28040 31328 28046 31340
rect 28092 31337 28120 31436
rect 28442 31424 28448 31436
rect 28500 31424 28506 31476
rect 28902 31424 28908 31476
rect 28960 31464 28966 31476
rect 29273 31467 29331 31473
rect 29273 31464 29285 31467
rect 28960 31436 29285 31464
rect 28960 31424 28966 31436
rect 29273 31433 29285 31436
rect 29319 31433 29331 31467
rect 29273 31427 29331 31433
rect 32306 31424 32312 31476
rect 32364 31464 32370 31476
rect 32364 31436 32720 31464
rect 32364 31424 32370 31436
rect 30282 31396 30288 31408
rect 28184 31368 30288 31396
rect 28184 31337 28212 31368
rect 30282 31356 30288 31368
rect 30340 31356 30346 31408
rect 31938 31356 31944 31408
rect 31996 31396 32002 31408
rect 31996 31368 32352 31396
rect 31996 31356 32002 31368
rect 28077 31331 28135 31337
rect 28077 31328 28089 31331
rect 28040 31300 28089 31328
rect 28040 31288 28046 31300
rect 28077 31297 28089 31300
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 28169 31331 28227 31337
rect 28169 31297 28181 31331
rect 28215 31297 28227 31331
rect 28169 31291 28227 31297
rect 28445 31331 28503 31337
rect 28445 31297 28457 31331
rect 28491 31328 28503 31331
rect 28810 31328 28816 31340
rect 28491 31300 28816 31328
rect 28491 31297 28503 31300
rect 28445 31291 28503 31297
rect 28810 31288 28816 31300
rect 28868 31328 28874 31340
rect 28905 31331 28963 31337
rect 28905 31328 28917 31331
rect 28868 31300 28917 31328
rect 28868 31288 28874 31300
rect 28905 31297 28917 31300
rect 28951 31297 28963 31331
rect 28905 31291 28963 31297
rect 28994 31288 29000 31340
rect 29052 31328 29058 31340
rect 29089 31331 29147 31337
rect 29089 31328 29101 31331
rect 29052 31300 29101 31328
rect 29052 31288 29058 31300
rect 29089 31297 29101 31300
rect 29135 31297 29147 31331
rect 29089 31291 29147 31297
rect 29822 31288 29828 31340
rect 29880 31328 29886 31340
rect 29917 31331 29975 31337
rect 29917 31328 29929 31331
rect 29880 31300 29929 31328
rect 29880 31288 29886 31300
rect 29917 31297 29929 31300
rect 29963 31297 29975 31331
rect 29917 31291 29975 31297
rect 31110 31288 31116 31340
rect 31168 31328 31174 31340
rect 32324 31337 32352 31368
rect 32692 31337 32720 31436
rect 32125 31331 32183 31337
rect 32125 31328 32137 31331
rect 31168 31300 32137 31328
rect 31168 31288 31174 31300
rect 32125 31297 32137 31300
rect 32171 31297 32183 31331
rect 32125 31291 32183 31297
rect 32309 31331 32367 31337
rect 32309 31297 32321 31331
rect 32355 31297 32367 31331
rect 32309 31291 32367 31297
rect 32677 31331 32735 31337
rect 32677 31297 32689 31331
rect 32723 31297 32735 31331
rect 32677 31291 32735 31297
rect 25869 31263 25927 31269
rect 25869 31260 25881 31263
rect 23584 31232 24440 31260
rect 25056 31232 25881 31260
rect 23584 31136 23612 31232
rect 23566 31124 23572 31136
rect 17920 31096 22784 31124
rect 23527 31096 23572 31124
rect 17920 31084 17926 31096
rect 23566 31084 23572 31096
rect 23624 31084 23630 31136
rect 24397 31127 24455 31133
rect 24397 31093 24409 31127
rect 24443 31124 24455 31127
rect 25056 31124 25084 31232
rect 25869 31229 25881 31232
rect 25915 31229 25927 31263
rect 25869 31223 25927 31229
rect 26326 31220 26332 31272
rect 26384 31260 26390 31272
rect 28350 31260 28356 31272
rect 26384 31232 28356 31260
rect 26384 31220 26390 31232
rect 28350 31220 28356 31232
rect 28408 31220 28414 31272
rect 30098 31220 30104 31272
rect 30156 31260 30162 31272
rect 30193 31263 30251 31269
rect 30193 31260 30205 31263
rect 30156 31232 30205 31260
rect 30156 31220 30162 31232
rect 30193 31229 30205 31232
rect 30239 31260 30251 31263
rect 30282 31260 30288 31272
rect 30239 31232 30288 31260
rect 30239 31229 30251 31232
rect 30193 31223 30251 31229
rect 30282 31220 30288 31232
rect 30340 31220 30346 31272
rect 32398 31260 32404 31272
rect 32359 31232 32404 31260
rect 32398 31220 32404 31232
rect 32456 31220 32462 31272
rect 32493 31263 32551 31269
rect 32493 31229 32505 31263
rect 32539 31260 32551 31263
rect 40218 31260 40224 31272
rect 32539 31232 40224 31260
rect 32539 31229 32551 31232
rect 32493 31223 32551 31229
rect 40218 31220 40224 31232
rect 40276 31220 40282 31272
rect 25222 31152 25228 31204
rect 25280 31192 25286 31204
rect 30834 31192 30840 31204
rect 25280 31164 30840 31192
rect 25280 31152 25286 31164
rect 30834 31152 30840 31164
rect 30892 31152 30898 31204
rect 30006 31124 30012 31136
rect 24443 31096 25084 31124
rect 29967 31096 30012 31124
rect 24443 31093 24455 31096
rect 24397 31087 24455 31093
rect 30006 31084 30012 31096
rect 30064 31084 30070 31136
rect 30098 31084 30104 31136
rect 30156 31124 30162 31136
rect 30156 31096 30201 31124
rect 30156 31084 30162 31096
rect 32214 31084 32220 31136
rect 32272 31124 32278 31136
rect 32861 31127 32919 31133
rect 32861 31124 32873 31127
rect 32272 31096 32873 31124
rect 32272 31084 32278 31096
rect 32861 31093 32873 31096
rect 32907 31093 32919 31127
rect 32861 31087 32919 31093
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 16025 30923 16083 30929
rect 16025 30889 16037 30923
rect 16071 30920 16083 30923
rect 17126 30920 17132 30932
rect 16071 30892 17132 30920
rect 16071 30889 16083 30892
rect 16025 30883 16083 30889
rect 17126 30880 17132 30892
rect 17184 30880 17190 30932
rect 17862 30920 17868 30932
rect 17823 30892 17868 30920
rect 17862 30880 17868 30892
rect 17920 30880 17926 30932
rect 19334 30920 19340 30932
rect 19295 30892 19340 30920
rect 19334 30880 19340 30892
rect 19392 30880 19398 30932
rect 20806 30880 20812 30932
rect 20864 30920 20870 30932
rect 20993 30923 21051 30929
rect 20993 30920 21005 30923
rect 20864 30892 21005 30920
rect 20864 30880 20870 30892
rect 20993 30889 21005 30892
rect 21039 30889 21051 30923
rect 20993 30883 21051 30889
rect 23106 30880 23112 30932
rect 23164 30920 23170 30932
rect 25222 30920 25228 30932
rect 23164 30892 25228 30920
rect 23164 30880 23170 30892
rect 25222 30880 25228 30892
rect 25280 30880 25286 30932
rect 26234 30920 26240 30932
rect 25976 30892 26240 30920
rect 17218 30812 17224 30864
rect 17276 30812 17282 30864
rect 20714 30812 20720 30864
rect 20772 30852 20778 30864
rect 25130 30852 25136 30864
rect 20772 30824 25136 30852
rect 20772 30812 20778 30824
rect 25130 30812 25136 30824
rect 25188 30812 25194 30864
rect 14277 30787 14335 30793
rect 14277 30753 14289 30787
rect 14323 30784 14335 30787
rect 17236 30784 17264 30812
rect 14323 30756 17264 30784
rect 20809 30787 20867 30793
rect 14323 30753 14335 30756
rect 14277 30747 14335 30753
rect 20809 30753 20821 30787
rect 20855 30784 20867 30787
rect 20990 30784 20996 30796
rect 20855 30756 20996 30784
rect 20855 30753 20867 30756
rect 20809 30747 20867 30753
rect 20990 30744 20996 30756
rect 21048 30744 21054 30796
rect 23293 30787 23351 30793
rect 23293 30753 23305 30787
rect 23339 30784 23351 30787
rect 23566 30784 23572 30796
rect 23339 30756 23572 30784
rect 23339 30753 23351 30756
rect 23293 30747 23351 30753
rect 23566 30744 23572 30756
rect 23624 30744 23630 30796
rect 25976 30793 26004 30892
rect 26234 30880 26240 30892
rect 26292 30880 26298 30932
rect 27430 30920 27436 30932
rect 27391 30892 27436 30920
rect 27430 30880 27436 30892
rect 27488 30880 27494 30932
rect 29546 30880 29552 30932
rect 29604 30920 29610 30932
rect 29733 30923 29791 30929
rect 29733 30920 29745 30923
rect 29604 30892 29745 30920
rect 29604 30880 29610 30892
rect 29733 30889 29745 30892
rect 29779 30889 29791 30923
rect 30742 30920 30748 30932
rect 30703 30892 30748 30920
rect 29733 30883 29791 30889
rect 30742 30880 30748 30892
rect 30800 30880 30806 30932
rect 31110 30920 31116 30932
rect 31071 30892 31116 30920
rect 31110 30880 31116 30892
rect 31168 30880 31174 30932
rect 28721 30855 28779 30861
rect 28721 30821 28733 30855
rect 28767 30852 28779 30855
rect 29914 30852 29920 30864
rect 28767 30824 29920 30852
rect 28767 30821 28779 30824
rect 28721 30815 28779 30821
rect 29914 30812 29920 30824
rect 29972 30812 29978 30864
rect 25961 30787 26019 30793
rect 25961 30753 25973 30787
rect 26007 30753 26019 30787
rect 25961 30747 26019 30753
rect 26237 30787 26295 30793
rect 26237 30753 26249 30787
rect 26283 30753 26295 30787
rect 26237 30747 26295 30753
rect 16942 30676 16948 30728
rect 17000 30716 17006 30728
rect 17037 30719 17095 30725
rect 17037 30716 17049 30719
rect 17000 30688 17049 30716
rect 17000 30676 17006 30688
rect 17037 30685 17049 30688
rect 17083 30685 17095 30719
rect 17037 30679 17095 30685
rect 17221 30719 17279 30725
rect 17221 30685 17233 30719
rect 17267 30716 17279 30719
rect 17310 30716 17316 30728
rect 17267 30688 17316 30716
rect 17267 30685 17279 30688
rect 17221 30679 17279 30685
rect 14553 30651 14611 30657
rect 14553 30617 14565 30651
rect 14599 30617 14611 30651
rect 15838 30648 15844 30660
rect 15778 30620 15844 30648
rect 14553 30611 14611 30617
rect 14568 30580 14596 30611
rect 15838 30608 15844 30620
rect 15896 30608 15902 30660
rect 17052 30648 17080 30679
rect 17310 30676 17316 30688
rect 17368 30716 17374 30728
rect 17865 30719 17923 30725
rect 17865 30716 17877 30719
rect 17368 30688 17877 30716
rect 17368 30676 17374 30688
rect 17865 30685 17877 30688
rect 17911 30685 17923 30719
rect 17865 30679 17923 30685
rect 18049 30719 18107 30725
rect 18049 30685 18061 30719
rect 18095 30685 18107 30719
rect 19242 30716 19248 30728
rect 19203 30688 19248 30716
rect 18049 30679 18107 30685
rect 17770 30648 17776 30660
rect 17052 30620 17776 30648
rect 17770 30608 17776 30620
rect 17828 30648 17834 30660
rect 18064 30648 18092 30679
rect 19242 30676 19248 30688
rect 19300 30676 19306 30728
rect 20717 30719 20775 30725
rect 20717 30685 20729 30719
rect 20763 30716 20775 30719
rect 22002 30716 22008 30728
rect 20763 30688 22008 30716
rect 20763 30685 20775 30688
rect 20717 30679 20775 30685
rect 22002 30676 22008 30688
rect 22060 30676 22066 30728
rect 22278 30676 22284 30728
rect 22336 30716 22342 30728
rect 23017 30719 23075 30725
rect 23017 30716 23029 30719
rect 22336 30688 23029 30716
rect 22336 30676 22342 30688
rect 23017 30685 23029 30688
rect 23063 30685 23075 30719
rect 23017 30679 23075 30685
rect 25590 30676 25596 30728
rect 25648 30716 25654 30728
rect 25869 30719 25927 30725
rect 25869 30716 25881 30719
rect 25648 30688 25881 30716
rect 25648 30676 25654 30688
rect 25869 30685 25881 30688
rect 25915 30685 25927 30719
rect 26252 30716 26280 30747
rect 26602 30744 26608 30796
rect 26660 30784 26666 30796
rect 30098 30784 30104 30796
rect 26660 30756 26924 30784
rect 26660 30744 26666 30756
rect 26896 30725 26924 30756
rect 29012 30756 30104 30784
rect 29012 30725 29040 30756
rect 30098 30744 30104 30756
rect 30156 30744 30162 30796
rect 30834 30784 30840 30796
rect 30795 30756 30840 30784
rect 30834 30744 30840 30756
rect 30892 30744 30898 30796
rect 32214 30784 32220 30796
rect 32175 30756 32220 30784
rect 32214 30744 32220 30756
rect 32272 30744 32278 30796
rect 26697 30719 26755 30725
rect 26697 30716 26709 30719
rect 26252 30688 26709 30716
rect 25869 30679 25927 30685
rect 26697 30685 26709 30688
rect 26743 30685 26755 30719
rect 26697 30679 26755 30685
rect 26881 30719 26939 30725
rect 26881 30685 26893 30719
rect 26927 30685 26939 30719
rect 26881 30679 26939 30685
rect 27341 30719 27399 30725
rect 27341 30685 27353 30719
rect 27387 30685 27399 30719
rect 27341 30679 27399 30685
rect 28997 30719 29055 30725
rect 28997 30685 29009 30719
rect 29043 30685 29055 30719
rect 29549 30719 29607 30725
rect 29549 30716 29561 30719
rect 28997 30679 29055 30685
rect 29196 30688 29561 30716
rect 17828 30620 18092 30648
rect 17828 30608 17834 30620
rect 20070 30608 20076 30660
rect 20128 30648 20134 30660
rect 23290 30648 23296 30660
rect 20128 30620 23296 30648
rect 20128 30608 20134 30620
rect 23290 30608 23296 30620
rect 23348 30608 23354 30660
rect 25682 30608 25688 30660
rect 25740 30648 25746 30660
rect 26970 30648 26976 30660
rect 25740 30620 26976 30648
rect 25740 30608 25746 30620
rect 26970 30608 26976 30620
rect 27028 30648 27034 30660
rect 27356 30648 27384 30679
rect 29196 30660 29224 30688
rect 29549 30685 29561 30688
rect 29595 30685 29607 30719
rect 29549 30679 29607 30685
rect 30006 30676 30012 30728
rect 30064 30716 30070 30728
rect 30561 30719 30619 30725
rect 30561 30716 30573 30719
rect 30064 30688 30573 30716
rect 30064 30676 30070 30688
rect 30561 30685 30573 30688
rect 30607 30685 30619 30719
rect 30561 30679 30619 30685
rect 30926 30676 30932 30728
rect 30984 30716 30990 30728
rect 31941 30719 31999 30725
rect 31941 30716 31953 30719
rect 30984 30688 31953 30716
rect 30984 30676 30990 30688
rect 31941 30685 31953 30688
rect 31987 30685 31999 30719
rect 31941 30679 31999 30685
rect 27028 30620 27384 30648
rect 28721 30651 28779 30657
rect 27028 30608 27034 30620
rect 28721 30617 28733 30651
rect 28767 30648 28779 30651
rect 29178 30648 29184 30660
rect 28767 30620 29184 30648
rect 28767 30617 28779 30620
rect 28721 30611 28779 30617
rect 29178 30608 29184 30620
rect 29236 30608 29242 30660
rect 33226 30608 33232 30660
rect 33284 30608 33290 30660
rect 15470 30580 15476 30592
rect 14568 30552 15476 30580
rect 15470 30540 15476 30552
rect 15528 30540 15534 30592
rect 17402 30580 17408 30592
rect 17363 30552 17408 30580
rect 17402 30540 17408 30552
rect 17460 30540 17466 30592
rect 25130 30540 25136 30592
rect 25188 30580 25194 30592
rect 26050 30580 26056 30592
rect 25188 30552 26056 30580
rect 25188 30540 25194 30552
rect 26050 30540 26056 30552
rect 26108 30580 26114 30592
rect 26602 30580 26608 30592
rect 26108 30552 26608 30580
rect 26108 30540 26114 30552
rect 26602 30540 26608 30552
rect 26660 30540 26666 30592
rect 26786 30580 26792 30592
rect 26747 30552 26792 30580
rect 26786 30540 26792 30552
rect 26844 30540 26850 30592
rect 28905 30583 28963 30589
rect 28905 30549 28917 30583
rect 28951 30580 28963 30583
rect 28994 30580 29000 30592
rect 28951 30552 29000 30580
rect 28951 30549 28963 30552
rect 28905 30543 28963 30549
rect 28994 30540 29000 30552
rect 29052 30540 29058 30592
rect 32398 30540 32404 30592
rect 32456 30580 32462 30592
rect 33689 30583 33747 30589
rect 33689 30580 33701 30583
rect 32456 30552 33701 30580
rect 32456 30540 32462 30552
rect 33689 30549 33701 30552
rect 33735 30549 33747 30583
rect 33689 30543 33747 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 15286 30336 15292 30388
rect 15344 30336 15350 30388
rect 15470 30376 15476 30388
rect 15431 30348 15476 30376
rect 15470 30336 15476 30348
rect 15528 30336 15534 30388
rect 16850 30336 16856 30388
rect 16908 30376 16914 30388
rect 19334 30376 19340 30388
rect 16908 30348 19340 30376
rect 16908 30336 16914 30348
rect 19334 30336 19340 30348
rect 19392 30336 19398 30388
rect 25130 30376 25136 30388
rect 24228 30348 24992 30376
rect 25091 30348 25136 30376
rect 15304 30308 15332 30336
rect 14844 30280 15332 30308
rect 14844 30249 14872 30280
rect 15838 30268 15844 30320
rect 15896 30308 15902 30320
rect 16025 30311 16083 30317
rect 16025 30308 16037 30311
rect 15896 30280 16037 30308
rect 15896 30268 15902 30280
rect 16025 30277 16037 30280
rect 16071 30277 16083 30311
rect 23750 30308 23756 30320
rect 16025 30271 16083 30277
rect 17328 30280 23756 30308
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30209 14887 30243
rect 14829 30203 14887 30209
rect 14918 30200 14924 30252
rect 14976 30240 14982 30252
rect 15105 30243 15163 30249
rect 14976 30212 15021 30240
rect 14976 30200 14982 30212
rect 15105 30209 15117 30243
rect 15151 30209 15163 30243
rect 15105 30203 15163 30209
rect 15120 30104 15148 30203
rect 15194 30200 15200 30252
rect 15252 30240 15258 30252
rect 15335 30243 15393 30249
rect 15252 30212 15297 30240
rect 15252 30200 15258 30212
rect 15335 30209 15347 30243
rect 15381 30240 15393 30243
rect 15381 30212 15884 30240
rect 15381 30209 15393 30212
rect 15335 30203 15393 30209
rect 15856 30172 15884 30212
rect 15930 30200 15936 30252
rect 15988 30240 15994 30252
rect 17328 30249 17356 30280
rect 23750 30268 23756 30280
rect 23808 30268 23814 30320
rect 17313 30243 17371 30249
rect 15988 30212 16988 30240
rect 15988 30200 15994 30212
rect 16114 30172 16120 30184
rect 15856 30144 16120 30172
rect 16114 30132 16120 30144
rect 16172 30132 16178 30184
rect 16960 30172 16988 30212
rect 17313 30209 17325 30243
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 17402 30200 17408 30252
rect 17460 30240 17466 30252
rect 17497 30243 17555 30249
rect 17497 30240 17509 30243
rect 17460 30212 17509 30240
rect 17460 30200 17466 30212
rect 17497 30209 17509 30212
rect 17543 30209 17555 30243
rect 17497 30203 17555 30209
rect 17589 30243 17647 30249
rect 17589 30209 17601 30243
rect 17635 30240 17647 30243
rect 17862 30240 17868 30252
rect 17635 30212 17868 30240
rect 17635 30209 17647 30212
rect 17589 30203 17647 30209
rect 17862 30200 17868 30212
rect 17920 30200 17926 30252
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30240 18843 30243
rect 19426 30240 19432 30252
rect 18831 30212 19432 30240
rect 18831 30209 18843 30212
rect 18785 30203 18843 30209
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 20717 30243 20775 30249
rect 20717 30209 20729 30243
rect 20763 30240 20775 30243
rect 20806 30240 20812 30252
rect 20763 30212 20812 30240
rect 20763 30209 20775 30212
rect 20717 30203 20775 30209
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 20901 30243 20959 30249
rect 20901 30209 20913 30243
rect 20947 30240 20959 30243
rect 20990 30240 20996 30252
rect 20947 30212 20996 30240
rect 20947 30209 20959 30212
rect 20901 30203 20959 30209
rect 20990 30200 20996 30212
rect 21048 30200 21054 30252
rect 22278 30200 22284 30252
rect 22336 30240 22342 30252
rect 23937 30243 23995 30249
rect 23937 30240 23949 30243
rect 22336 30212 23949 30240
rect 22336 30200 22342 30212
rect 23937 30209 23949 30212
rect 23983 30209 23995 30243
rect 24228 30240 24256 30348
rect 24854 30308 24860 30320
rect 24320 30280 24860 30308
rect 24320 30249 24348 30280
rect 24854 30268 24860 30280
rect 24912 30268 24918 30320
rect 24964 30308 24992 30348
rect 25130 30336 25136 30348
rect 25188 30336 25194 30388
rect 25682 30336 25688 30388
rect 25740 30376 25746 30388
rect 25869 30379 25927 30385
rect 25869 30376 25881 30379
rect 25740 30348 25881 30376
rect 25740 30336 25746 30348
rect 25869 30345 25881 30348
rect 25915 30345 25927 30379
rect 25869 30339 25927 30345
rect 28994 30336 29000 30388
rect 29052 30376 29058 30388
rect 30282 30376 30288 30388
rect 29052 30348 30288 30376
rect 29052 30336 29058 30348
rect 30282 30336 30288 30348
rect 30340 30376 30346 30388
rect 31113 30379 31171 30385
rect 31113 30376 31125 30379
rect 30340 30348 31125 30376
rect 30340 30336 30346 30348
rect 31113 30345 31125 30348
rect 31159 30345 31171 30379
rect 31113 30339 31171 30345
rect 27065 30311 27123 30317
rect 24964 30280 25728 30308
rect 23937 30203 23995 30209
rect 24044 30212 24256 30240
rect 24305 30243 24363 30249
rect 19444 30172 19472 30200
rect 24044 30172 24072 30212
rect 24305 30209 24317 30243
rect 24351 30209 24363 30243
rect 24305 30203 24363 30209
rect 24394 30200 24400 30252
rect 24452 30240 24458 30252
rect 25700 30249 25728 30280
rect 27065 30277 27077 30311
rect 27111 30308 27123 30311
rect 27522 30308 27528 30320
rect 27111 30280 27528 30308
rect 27111 30277 27123 30280
rect 27065 30271 27123 30277
rect 27522 30268 27528 30280
rect 27580 30268 27586 30320
rect 28445 30311 28503 30317
rect 28445 30277 28457 30311
rect 28491 30308 28503 30311
rect 29641 30311 29699 30317
rect 29641 30308 29653 30311
rect 28491 30280 29653 30308
rect 28491 30277 28503 30280
rect 28445 30271 28503 30277
rect 29641 30277 29653 30280
rect 29687 30277 29699 30311
rect 29641 30271 29699 30277
rect 30650 30268 30656 30320
rect 30708 30268 30714 30320
rect 32953 30311 33011 30317
rect 32953 30277 32965 30311
rect 32999 30308 33011 30311
rect 33226 30308 33232 30320
rect 32999 30280 33232 30308
rect 32999 30277 33011 30280
rect 32953 30271 33011 30277
rect 33226 30268 33232 30280
rect 33284 30268 33290 30320
rect 24949 30243 25007 30249
rect 24949 30240 24961 30243
rect 24452 30212 24961 30240
rect 24452 30200 24458 30212
rect 24949 30209 24961 30212
rect 24995 30209 25007 30243
rect 24949 30203 25007 30209
rect 25685 30243 25743 30249
rect 25685 30209 25697 30243
rect 25731 30240 25743 30243
rect 25866 30240 25872 30252
rect 25731 30212 25872 30240
rect 25731 30209 25743 30212
rect 25685 30203 25743 30209
rect 25866 30200 25872 30212
rect 25924 30240 25930 30252
rect 27709 30243 27767 30249
rect 27709 30240 27721 30243
rect 25924 30212 27721 30240
rect 25924 30200 25930 30212
rect 27709 30209 27721 30212
rect 27755 30209 27767 30243
rect 28626 30240 28632 30252
rect 28587 30212 28632 30240
rect 27709 30203 27767 30209
rect 28626 30200 28632 30212
rect 28684 30200 28690 30252
rect 32858 30240 32864 30252
rect 32819 30212 32864 30240
rect 32858 30200 32864 30212
rect 32916 30200 32922 30252
rect 24486 30172 24492 30184
rect 16960 30144 19012 30172
rect 19444 30144 24072 30172
rect 24136 30144 24492 30172
rect 16850 30104 16856 30116
rect 15120 30076 16856 30104
rect 16850 30064 16856 30076
rect 16908 30104 16914 30116
rect 18230 30104 18236 30116
rect 16908 30076 18236 30104
rect 16908 30064 16914 30076
rect 18230 30064 18236 30076
rect 18288 30064 18294 30116
rect 18984 30113 19012 30144
rect 18969 30107 19027 30113
rect 18969 30073 18981 30107
rect 19015 30073 19027 30107
rect 18969 30067 19027 30073
rect 19334 30064 19340 30116
rect 19392 30104 19398 30116
rect 21634 30104 21640 30116
rect 19392 30076 21640 30104
rect 19392 30064 19398 30076
rect 21634 30064 21640 30076
rect 21692 30064 21698 30116
rect 23750 30064 23756 30116
rect 23808 30104 23814 30116
rect 24136 30104 24164 30144
rect 24486 30132 24492 30144
rect 24544 30132 24550 30184
rect 25130 30132 25136 30184
rect 25188 30172 25194 30184
rect 28534 30172 28540 30184
rect 25188 30144 28540 30172
rect 25188 30132 25194 30144
rect 28534 30132 28540 30144
rect 28592 30172 28598 30184
rect 28813 30175 28871 30181
rect 28813 30172 28825 30175
rect 28592 30144 28825 30172
rect 28592 30132 28598 30144
rect 28813 30141 28825 30144
rect 28859 30141 28871 30175
rect 28813 30135 28871 30141
rect 28905 30175 28963 30181
rect 28905 30141 28917 30175
rect 28951 30172 28963 30175
rect 28994 30172 29000 30184
rect 28951 30144 29000 30172
rect 28951 30141 28963 30144
rect 28905 30135 28963 30141
rect 28994 30132 29000 30144
rect 29052 30132 29058 30184
rect 29365 30175 29423 30181
rect 29365 30141 29377 30175
rect 29411 30172 29423 30175
rect 34330 30172 34336 30184
rect 29411 30144 29500 30172
rect 34291 30144 34336 30172
rect 29411 30141 29423 30144
rect 29365 30135 29423 30141
rect 25958 30104 25964 30116
rect 23808 30076 24164 30104
rect 24320 30076 25964 30104
rect 23808 30064 23814 30076
rect 16666 29996 16672 30048
rect 16724 30036 16730 30048
rect 17129 30039 17187 30045
rect 17129 30036 17141 30039
rect 16724 30008 17141 30036
rect 16724 29996 16730 30008
rect 17129 30005 17141 30008
rect 17175 30005 17187 30039
rect 17129 29999 17187 30005
rect 20714 29996 20720 30048
rect 20772 30036 20778 30048
rect 24320 30045 24348 30076
rect 25958 30064 25964 30076
rect 26016 30064 26022 30116
rect 27246 30104 27252 30116
rect 27159 30076 27252 30104
rect 27246 30064 27252 30076
rect 27304 30104 27310 30116
rect 29472 30104 29500 30144
rect 34330 30132 34336 30144
rect 34388 30132 34394 30184
rect 34517 30175 34575 30181
rect 34517 30141 34529 30175
rect 34563 30172 34575 30175
rect 34790 30172 34796 30184
rect 34563 30144 34796 30172
rect 34563 30141 34575 30144
rect 34517 30135 34575 30141
rect 34790 30132 34796 30144
rect 34848 30132 34854 30184
rect 34882 30132 34888 30184
rect 34940 30172 34946 30184
rect 34940 30144 34985 30172
rect 34940 30132 34946 30144
rect 27304 30076 29500 30104
rect 27304 30064 27310 30076
rect 20809 30039 20867 30045
rect 20809 30036 20821 30039
rect 20772 30008 20821 30036
rect 20772 29996 20778 30008
rect 20809 30005 20821 30008
rect 20855 30005 20867 30039
rect 20809 29999 20867 30005
rect 24305 30039 24363 30045
rect 24305 30005 24317 30039
rect 24351 30005 24363 30039
rect 24486 30036 24492 30048
rect 24447 30008 24492 30036
rect 24305 29999 24363 30005
rect 24486 29996 24492 30008
rect 24544 29996 24550 30048
rect 27893 30039 27951 30045
rect 27893 30005 27905 30039
rect 27939 30036 27951 30039
rect 28166 30036 28172 30048
rect 27939 30008 28172 30036
rect 27939 30005 27951 30008
rect 27893 29999 27951 30005
rect 28166 29996 28172 30008
rect 28224 29996 28230 30048
rect 29472 30036 29500 30076
rect 29822 30036 29828 30048
rect 29472 30008 29828 30036
rect 29822 29996 29828 30008
rect 29880 30036 29886 30048
rect 30926 30036 30932 30048
rect 29880 30008 30932 30036
rect 29880 29996 29886 30008
rect 30926 29996 30932 30008
rect 30984 29996 30990 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 17770 29792 17776 29844
rect 17828 29832 17834 29844
rect 17865 29835 17923 29841
rect 17865 29832 17877 29835
rect 17828 29804 17877 29832
rect 17828 29792 17834 29804
rect 17865 29801 17877 29804
rect 17911 29801 17923 29835
rect 17865 29795 17923 29801
rect 20806 29792 20812 29844
rect 20864 29832 20870 29844
rect 20901 29835 20959 29841
rect 20901 29832 20913 29835
rect 20864 29804 20913 29832
rect 20864 29792 20870 29804
rect 20901 29801 20913 29804
rect 20947 29801 20959 29835
rect 20901 29795 20959 29801
rect 20990 29792 20996 29844
rect 21048 29832 21054 29844
rect 21910 29832 21916 29844
rect 21048 29804 21916 29832
rect 21048 29792 21054 29804
rect 21910 29792 21916 29804
rect 21968 29792 21974 29844
rect 22646 29792 22652 29844
rect 22704 29832 22710 29844
rect 22830 29832 22836 29844
rect 22704 29804 22836 29832
rect 22704 29792 22710 29804
rect 22830 29792 22836 29804
rect 22888 29832 22894 29844
rect 25130 29832 25136 29844
rect 22888 29804 25136 29832
rect 22888 29792 22894 29804
rect 25130 29792 25136 29804
rect 25188 29792 25194 29844
rect 25884 29804 27108 29832
rect 21634 29724 21640 29776
rect 21692 29764 21698 29776
rect 25041 29767 25099 29773
rect 25041 29764 25053 29767
rect 21692 29736 25053 29764
rect 21692 29724 21698 29736
rect 25041 29733 25053 29736
rect 25087 29764 25099 29767
rect 25884 29764 25912 29804
rect 25087 29736 25912 29764
rect 27080 29764 27108 29804
rect 28626 29792 28632 29844
rect 28684 29832 28690 29844
rect 29549 29835 29607 29841
rect 29549 29832 29561 29835
rect 28684 29804 29561 29832
rect 28684 29792 28690 29804
rect 29549 29801 29561 29804
rect 29595 29801 29607 29835
rect 30650 29832 30656 29844
rect 30611 29804 30656 29832
rect 29549 29795 29607 29801
rect 30650 29792 30656 29804
rect 30708 29792 30714 29844
rect 34790 29832 34796 29844
rect 34751 29804 34796 29832
rect 34790 29792 34796 29804
rect 34848 29792 34854 29844
rect 27982 29764 27988 29776
rect 27080 29736 27988 29764
rect 25087 29733 25099 29736
rect 25041 29727 25099 29733
rect 27982 29724 27988 29736
rect 28040 29724 28046 29776
rect 28994 29724 29000 29776
rect 29052 29764 29058 29776
rect 29454 29764 29460 29776
rect 29052 29736 29460 29764
rect 29052 29724 29058 29736
rect 29454 29724 29460 29736
rect 29512 29764 29518 29776
rect 30006 29764 30012 29776
rect 29512 29736 30012 29764
rect 29512 29724 29518 29736
rect 30006 29724 30012 29736
rect 30064 29724 30070 29776
rect 16117 29699 16175 29705
rect 16117 29665 16129 29699
rect 16163 29696 16175 29699
rect 17126 29696 17132 29708
rect 16163 29668 17132 29696
rect 16163 29665 16175 29668
rect 16117 29659 16175 29665
rect 17126 29656 17132 29668
rect 17184 29656 17190 29708
rect 21174 29696 21180 29708
rect 20180 29668 21180 29696
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29628 18383 29631
rect 19242 29628 19248 29640
rect 18371 29600 19248 29628
rect 18371 29597 18383 29600
rect 18325 29591 18383 29597
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 20180 29637 20208 29668
rect 21174 29656 21180 29668
rect 21232 29656 21238 29708
rect 22646 29656 22652 29708
rect 22704 29696 22710 29708
rect 25777 29699 25835 29705
rect 25777 29696 25789 29699
rect 22704 29668 25789 29696
rect 22704 29656 22710 29668
rect 25777 29665 25789 29668
rect 25823 29696 25835 29699
rect 27246 29696 27252 29708
rect 25823 29668 27252 29696
rect 25823 29665 25835 29668
rect 25777 29659 25835 29665
rect 27246 29656 27252 29668
rect 27304 29656 27310 29708
rect 29546 29656 29552 29708
rect 29604 29696 29610 29708
rect 29604 29668 29868 29696
rect 29604 29656 29610 29668
rect 20165 29631 20223 29637
rect 20165 29597 20177 29631
rect 20211 29597 20223 29631
rect 20165 29591 20223 29597
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29597 20867 29631
rect 20809 29591 20867 29597
rect 20993 29631 21051 29637
rect 20993 29597 21005 29631
rect 21039 29628 21051 29631
rect 21266 29628 21272 29640
rect 21039 29600 21272 29628
rect 21039 29597 21051 29600
rect 20993 29591 21051 29597
rect 16390 29560 16396 29572
rect 16351 29532 16396 29560
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 18417 29563 18475 29569
rect 18417 29560 18429 29563
rect 17618 29532 18429 29560
rect 18417 29529 18429 29532
rect 18463 29529 18475 29563
rect 20824 29560 20852 29591
rect 21266 29588 21272 29600
rect 21324 29588 21330 29640
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29628 21787 29631
rect 21818 29628 21824 29640
rect 21775 29600 21824 29628
rect 21775 29597 21787 29600
rect 21729 29591 21787 29597
rect 21818 29588 21824 29600
rect 21876 29588 21882 29640
rect 22002 29628 22008 29640
rect 21963 29600 22008 29628
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 22554 29588 22560 29640
rect 22612 29628 22618 29640
rect 22925 29631 22983 29637
rect 22925 29628 22937 29631
rect 22612 29600 22937 29628
rect 22612 29588 22618 29600
rect 22925 29597 22937 29600
rect 22971 29597 22983 29631
rect 22925 29591 22983 29597
rect 23661 29631 23719 29637
rect 23661 29597 23673 29631
rect 23707 29628 23719 29631
rect 24486 29628 24492 29640
rect 23707 29600 24492 29628
rect 23707 29597 23719 29600
rect 23661 29591 23719 29597
rect 24486 29588 24492 29600
rect 24544 29628 24550 29640
rect 29840 29637 29868 29668
rect 29914 29656 29920 29708
rect 29972 29696 29978 29708
rect 29972 29668 30144 29696
rect 29972 29656 29978 29668
rect 24857 29631 24915 29637
rect 24857 29628 24869 29631
rect 24544 29600 24869 29628
rect 24544 29588 24550 29600
rect 24857 29597 24869 29600
rect 24903 29597 24915 29631
rect 24857 29591 24915 29597
rect 29733 29631 29791 29637
rect 29733 29597 29745 29631
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29825 29631 29883 29637
rect 29825 29597 29837 29631
rect 29871 29597 29883 29631
rect 30006 29628 30012 29640
rect 29967 29600 30012 29628
rect 29825 29591 29883 29597
rect 21634 29560 21640 29572
rect 20824 29532 21640 29560
rect 18417 29523 18475 29529
rect 21634 29520 21640 29532
rect 21692 29520 21698 29572
rect 26053 29563 26111 29569
rect 26053 29529 26065 29563
rect 26099 29560 26111 29563
rect 26326 29560 26332 29572
rect 26099 29532 26332 29560
rect 26099 29529 26111 29532
rect 26053 29523 26111 29529
rect 26326 29520 26332 29532
rect 26384 29520 26390 29572
rect 27062 29520 27068 29572
rect 27120 29520 27126 29572
rect 29748 29560 29776 29591
rect 30006 29588 30012 29600
rect 30064 29588 30070 29640
rect 30116 29637 30144 29668
rect 30392 29668 38654 29696
rect 30101 29631 30159 29637
rect 30101 29597 30113 29631
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 30392 29560 30420 29668
rect 30558 29628 30564 29640
rect 30519 29600 30564 29628
rect 30558 29588 30564 29600
rect 30616 29628 30622 29640
rect 32858 29628 32864 29640
rect 30616 29600 32864 29628
rect 30616 29588 30622 29600
rect 32858 29588 32864 29600
rect 32916 29588 32922 29640
rect 34701 29631 34759 29637
rect 34701 29597 34713 29631
rect 34747 29628 34759 29631
rect 35342 29628 35348 29640
rect 34747 29600 35348 29628
rect 34747 29597 34759 29600
rect 34701 29591 34759 29597
rect 35342 29588 35348 29600
rect 35400 29588 35406 29640
rect 29748 29532 30420 29560
rect 38626 29560 38654 29668
rect 47210 29656 47216 29708
rect 47268 29696 47274 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 47268 29668 47593 29696
rect 47268 29656 47274 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 47305 29631 47363 29637
rect 47305 29597 47317 29631
rect 47351 29628 47363 29631
rect 47394 29628 47400 29640
rect 47351 29600 47400 29628
rect 47351 29597 47363 29600
rect 47305 29591 47363 29597
rect 47394 29588 47400 29600
rect 47452 29588 47458 29640
rect 43898 29560 43904 29572
rect 38626 29532 43904 29560
rect 43898 29520 43904 29532
rect 43956 29520 43962 29572
rect 15194 29452 15200 29504
rect 15252 29492 15258 29504
rect 17126 29492 17132 29504
rect 15252 29464 17132 29492
rect 15252 29452 15258 29464
rect 17126 29452 17132 29464
rect 17184 29492 17190 29504
rect 20070 29492 20076 29504
rect 17184 29464 20076 29492
rect 17184 29452 17190 29464
rect 20070 29452 20076 29464
rect 20128 29452 20134 29504
rect 20254 29492 20260 29504
rect 20215 29464 20260 29492
rect 20254 29452 20260 29464
rect 20312 29452 20318 29504
rect 21545 29495 21603 29501
rect 21545 29461 21557 29495
rect 21591 29492 21603 29495
rect 21726 29492 21732 29504
rect 21591 29464 21732 29492
rect 21591 29461 21603 29464
rect 21545 29455 21603 29461
rect 21726 29452 21732 29464
rect 21784 29452 21790 29504
rect 23014 29492 23020 29504
rect 22975 29464 23020 29492
rect 23014 29452 23020 29464
rect 23072 29452 23078 29504
rect 23106 29452 23112 29504
rect 23164 29492 23170 29504
rect 23753 29495 23811 29501
rect 23753 29492 23765 29495
rect 23164 29464 23765 29492
rect 23164 29452 23170 29464
rect 23753 29461 23765 29464
rect 23799 29492 23811 29495
rect 23842 29492 23848 29504
rect 23799 29464 23848 29492
rect 23799 29461 23811 29464
rect 23753 29455 23811 29461
rect 23842 29452 23848 29464
rect 23900 29452 23906 29504
rect 25682 29452 25688 29504
rect 25740 29492 25746 29504
rect 26786 29492 26792 29504
rect 25740 29464 26792 29492
rect 25740 29452 25746 29464
rect 26786 29452 26792 29464
rect 26844 29452 26850 29504
rect 26878 29452 26884 29504
rect 26936 29492 26942 29504
rect 27525 29495 27583 29501
rect 27525 29492 27537 29495
rect 26936 29464 27537 29492
rect 26936 29452 26942 29464
rect 27525 29461 27537 29464
rect 27571 29461 27583 29495
rect 27525 29455 27583 29461
rect 28166 29452 28172 29504
rect 28224 29492 28230 29504
rect 30558 29492 30564 29504
rect 28224 29464 30564 29492
rect 28224 29452 28230 29464
rect 30558 29452 30564 29464
rect 30616 29452 30622 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 16390 29248 16396 29300
rect 16448 29288 16454 29300
rect 17313 29291 17371 29297
rect 17313 29288 17325 29291
rect 16448 29260 17325 29288
rect 16448 29248 16454 29260
rect 17313 29257 17325 29260
rect 17359 29257 17371 29291
rect 21266 29288 21272 29300
rect 21179 29260 21272 29288
rect 17313 29251 17371 29257
rect 21266 29248 21272 29260
rect 21324 29248 21330 29300
rect 21910 29248 21916 29300
rect 21968 29288 21974 29300
rect 22189 29291 22247 29297
rect 22189 29288 22201 29291
rect 21968 29260 22201 29288
rect 21968 29248 21974 29260
rect 22189 29257 22201 29260
rect 22235 29257 22247 29291
rect 22189 29251 22247 29257
rect 22922 29248 22928 29300
rect 22980 29288 22986 29300
rect 25225 29291 25283 29297
rect 25225 29288 25237 29291
rect 22980 29260 25237 29288
rect 22980 29248 22986 29260
rect 25225 29257 25237 29260
rect 25271 29257 25283 29291
rect 25225 29251 25283 29257
rect 17770 29220 17776 29232
rect 16776 29192 17776 29220
rect 16666 29152 16672 29164
rect 16627 29124 16672 29152
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 16776 29161 16804 29192
rect 17770 29180 17776 29192
rect 17828 29180 17834 29232
rect 20254 29180 20260 29232
rect 20312 29180 20318 29232
rect 21284 29220 21312 29248
rect 21634 29220 21640 29232
rect 21284 29192 21640 29220
rect 21634 29180 21640 29192
rect 21692 29220 21698 29232
rect 22005 29223 22063 29229
rect 22005 29220 22017 29223
rect 21692 29192 22017 29220
rect 21692 29180 21698 29192
rect 22005 29189 22017 29192
rect 22051 29189 22063 29223
rect 22005 29183 22063 29189
rect 23014 29180 23020 29232
rect 23072 29220 23078 29232
rect 25240 29220 25268 29251
rect 26326 29248 26332 29300
rect 26384 29288 26390 29300
rect 26421 29291 26479 29297
rect 26421 29288 26433 29291
rect 26384 29260 26433 29288
rect 26384 29248 26390 29260
rect 26421 29257 26433 29260
rect 26467 29257 26479 29291
rect 27062 29288 27068 29300
rect 27023 29260 27068 29288
rect 26421 29251 26479 29257
rect 27062 29248 27068 29260
rect 27120 29248 27126 29300
rect 26145 29223 26203 29229
rect 26145 29220 26157 29223
rect 23072 29192 23414 29220
rect 25240 29192 26157 29220
rect 23072 29180 23078 29192
rect 26145 29189 26157 29192
rect 26191 29220 26203 29223
rect 26510 29220 26516 29232
rect 26191 29192 26516 29220
rect 26191 29189 26203 29192
rect 26145 29183 26203 29189
rect 26510 29180 26516 29192
rect 26568 29180 26574 29232
rect 16762 29155 16820 29161
rect 16762 29121 16774 29155
rect 16808 29121 16820 29155
rect 16762 29115 16820 29121
rect 16850 29112 16856 29164
rect 16908 29152 16914 29164
rect 16945 29155 17003 29161
rect 16945 29152 16957 29155
rect 16908 29124 16957 29152
rect 16908 29112 16914 29124
rect 16945 29121 16957 29124
rect 16991 29121 17003 29155
rect 16945 29115 17003 29121
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17175 29155 17233 29161
rect 17175 29121 17187 29155
rect 17221 29152 17233 29155
rect 17494 29152 17500 29164
rect 17221 29124 17500 29152
rect 17221 29121 17233 29124
rect 17175 29115 17233 29121
rect 17052 29084 17080 29115
rect 17494 29112 17500 29124
rect 17552 29112 17558 29164
rect 21542 29112 21548 29164
rect 21600 29152 21606 29164
rect 21821 29155 21879 29161
rect 21821 29152 21833 29155
rect 21600 29124 21833 29152
rect 21600 29112 21606 29124
rect 21821 29121 21833 29124
rect 21867 29121 21879 29155
rect 22646 29152 22652 29164
rect 22607 29124 22652 29152
rect 21821 29115 21879 29121
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 25041 29155 25099 29161
rect 25041 29121 25053 29155
rect 25087 29152 25099 29155
rect 25130 29152 25136 29164
rect 25087 29124 25136 29152
rect 25087 29121 25099 29124
rect 25041 29115 25099 29121
rect 25130 29112 25136 29124
rect 25188 29112 25194 29164
rect 25682 29112 25688 29164
rect 25740 29152 25746 29164
rect 25777 29155 25835 29161
rect 25777 29152 25789 29155
rect 25740 29124 25789 29152
rect 25740 29112 25746 29124
rect 25777 29121 25789 29124
rect 25823 29121 25835 29155
rect 25777 29115 25835 29121
rect 25870 29155 25928 29161
rect 25870 29121 25882 29155
rect 25916 29121 25928 29155
rect 25870 29115 25928 29121
rect 19521 29087 19579 29093
rect 17052 29056 17172 29084
rect 17144 29028 17172 29056
rect 19521 29053 19533 29087
rect 19567 29053 19579 29087
rect 19794 29084 19800 29096
rect 19755 29056 19800 29084
rect 19521 29047 19579 29053
rect 17126 28976 17132 29028
rect 17184 28976 17190 29028
rect 17218 28976 17224 29028
rect 17276 29016 17282 29028
rect 19536 29016 19564 29047
rect 19794 29044 19800 29056
rect 19852 29044 19858 29096
rect 22922 29084 22928 29096
rect 22883 29056 22928 29084
rect 22922 29044 22928 29056
rect 22980 29044 22986 29096
rect 23290 29044 23296 29096
rect 23348 29084 23354 29096
rect 24397 29087 24455 29093
rect 24397 29084 24409 29087
rect 23348 29056 24409 29084
rect 23348 29044 23354 29056
rect 24397 29053 24409 29056
rect 24443 29053 24455 29087
rect 24397 29047 24455 29053
rect 25590 29044 25596 29096
rect 25648 29084 25654 29096
rect 25884 29084 25912 29115
rect 26050 29112 26056 29164
rect 26108 29152 26114 29164
rect 26283 29155 26341 29161
rect 26108 29124 26153 29152
rect 26108 29112 26114 29124
rect 26283 29121 26295 29155
rect 26329 29152 26341 29155
rect 26418 29152 26424 29164
rect 26329 29124 26424 29152
rect 26329 29121 26341 29124
rect 26283 29115 26341 29121
rect 26418 29112 26424 29124
rect 26476 29112 26482 29164
rect 26970 29152 26976 29164
rect 26931 29124 26976 29152
rect 26970 29112 26976 29124
rect 27028 29112 27034 29164
rect 28813 29155 28871 29161
rect 28813 29121 28825 29155
rect 28859 29152 28871 29155
rect 29178 29152 29184 29164
rect 28859 29124 29184 29152
rect 28859 29121 28871 29124
rect 28813 29115 28871 29121
rect 29178 29112 29184 29124
rect 29236 29112 29242 29164
rect 26878 29084 26884 29096
rect 25648 29056 26884 29084
rect 25648 29044 25654 29056
rect 26878 29044 26884 29056
rect 26936 29044 26942 29096
rect 32674 29084 32680 29096
rect 32635 29056 32680 29084
rect 32674 29044 32680 29056
rect 32732 29044 32738 29096
rect 32858 29084 32864 29096
rect 32819 29056 32864 29084
rect 32858 29044 32864 29056
rect 32916 29044 32922 29096
rect 33134 29084 33140 29096
rect 33095 29056 33140 29084
rect 33134 29044 33140 29056
rect 33192 29044 33198 29096
rect 17276 28988 19564 29016
rect 17276 28976 17282 28988
rect 25130 28908 25136 28960
rect 25188 28948 25194 28960
rect 28905 28951 28963 28957
rect 28905 28948 28917 28951
rect 25188 28920 28917 28948
rect 25188 28908 25194 28920
rect 28905 28917 28917 28920
rect 28951 28948 28963 28951
rect 29546 28948 29552 28960
rect 28951 28920 29552 28948
rect 28951 28917 28963 28920
rect 28905 28911 28963 28917
rect 29546 28908 29552 28920
rect 29604 28908 29610 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 19794 28704 19800 28756
rect 19852 28744 19858 28756
rect 20993 28747 21051 28753
rect 20993 28744 21005 28747
rect 19852 28716 21005 28744
rect 19852 28704 19858 28716
rect 20993 28713 21005 28716
rect 21039 28713 21051 28747
rect 21726 28744 21732 28756
rect 21687 28716 21732 28744
rect 20993 28707 21051 28713
rect 21726 28704 21732 28716
rect 21784 28704 21790 28756
rect 22189 28747 22247 28753
rect 22189 28713 22201 28747
rect 22235 28744 22247 28747
rect 22646 28744 22652 28756
rect 22235 28716 22652 28744
rect 22235 28713 22247 28716
rect 22189 28707 22247 28713
rect 22646 28704 22652 28716
rect 22704 28704 22710 28756
rect 22922 28704 22928 28756
rect 22980 28744 22986 28756
rect 23385 28747 23443 28753
rect 23385 28744 23397 28747
rect 22980 28716 23397 28744
rect 22980 28704 22986 28716
rect 23385 28713 23397 28716
rect 23431 28713 23443 28747
rect 23385 28707 23443 28713
rect 30009 28747 30067 28753
rect 30009 28713 30021 28747
rect 30055 28713 30067 28747
rect 30190 28744 30196 28756
rect 30151 28716 30196 28744
rect 30009 28707 30067 28713
rect 21266 28676 21272 28688
rect 17512 28648 21272 28676
rect 15010 28568 15016 28620
rect 15068 28608 15074 28620
rect 17512 28617 17540 28648
rect 21266 28636 21272 28648
rect 21324 28676 21330 28688
rect 26050 28676 26056 28688
rect 21324 28648 21680 28676
rect 21324 28636 21330 28648
rect 17497 28611 17555 28617
rect 15068 28580 16620 28608
rect 15068 28568 15074 28580
rect 16592 28549 16620 28580
rect 17497 28577 17509 28611
rect 17543 28577 17555 28611
rect 17497 28571 17555 28577
rect 18230 28568 18236 28620
rect 18288 28608 18294 28620
rect 18288 28580 20668 28608
rect 18288 28568 18294 28580
rect 16485 28543 16543 28549
rect 16485 28509 16497 28543
rect 16531 28509 16543 28543
rect 16485 28503 16543 28509
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28509 16635 28543
rect 16577 28503 16635 28509
rect 17405 28543 17463 28549
rect 17405 28509 17417 28543
rect 17451 28540 17463 28543
rect 17954 28540 17960 28552
rect 17451 28512 17960 28540
rect 17451 28509 17463 28512
rect 17405 28503 17463 28509
rect 16500 28472 16528 28503
rect 17954 28500 17960 28512
rect 18012 28500 18018 28552
rect 20346 28540 20352 28552
rect 20307 28512 20352 28540
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 20530 28549 20536 28552
rect 20497 28543 20536 28549
rect 20497 28509 20509 28543
rect 20497 28503 20536 28509
rect 20530 28500 20536 28503
rect 20588 28500 20594 28552
rect 20640 28540 20668 28580
rect 21652 28549 21680 28648
rect 21744 28648 26056 28676
rect 20814 28543 20872 28549
rect 20814 28540 20826 28543
rect 20640 28512 20826 28540
rect 20814 28509 20826 28512
rect 20860 28540 20872 28543
rect 21637 28543 21695 28549
rect 20860 28512 21588 28540
rect 20860 28509 20872 28512
rect 20814 28503 20872 28509
rect 20070 28472 20076 28484
rect 16500 28444 20076 28472
rect 20070 28432 20076 28444
rect 20128 28432 20134 28484
rect 20625 28475 20683 28481
rect 20625 28441 20637 28475
rect 20671 28441 20683 28475
rect 20625 28435 20683 28441
rect 20717 28475 20775 28481
rect 20717 28441 20729 28475
rect 20763 28441 20775 28475
rect 21560 28472 21588 28512
rect 21637 28509 21649 28543
rect 21683 28509 21695 28543
rect 21637 28503 21695 28509
rect 21744 28472 21772 28648
rect 26050 28636 26056 28648
rect 26108 28636 26114 28688
rect 29546 28636 29552 28688
rect 29604 28676 29610 28688
rect 30024 28676 30052 28707
rect 30190 28704 30196 28716
rect 30248 28704 30254 28756
rect 30653 28747 30711 28753
rect 30653 28713 30665 28747
rect 30699 28744 30711 28747
rect 30742 28744 30748 28756
rect 30699 28716 30748 28744
rect 30699 28713 30711 28716
rect 30653 28707 30711 28713
rect 30742 28704 30748 28716
rect 30800 28704 30806 28756
rect 32858 28744 32864 28756
rect 32819 28716 32864 28744
rect 32858 28704 32864 28716
rect 32916 28704 32922 28756
rect 34330 28704 34336 28756
rect 34388 28744 34394 28756
rect 36449 28747 36507 28753
rect 36449 28744 36461 28747
rect 34388 28716 36461 28744
rect 34388 28704 34394 28716
rect 36449 28713 36461 28716
rect 36495 28713 36507 28747
rect 36449 28707 36507 28713
rect 29604 28648 31156 28676
rect 29604 28636 29610 28648
rect 21818 28568 21824 28620
rect 21876 28608 21882 28620
rect 22925 28611 22983 28617
rect 22925 28608 22937 28611
rect 21876 28580 22937 28608
rect 21876 28568 21882 28580
rect 22925 28577 22937 28580
rect 22971 28608 22983 28611
rect 23290 28608 23296 28620
rect 22971 28580 23296 28608
rect 22971 28577 22983 28580
rect 22925 28571 22983 28577
rect 23290 28568 23296 28580
rect 23348 28568 23354 28620
rect 29454 28568 29460 28620
rect 29512 28608 29518 28620
rect 29825 28611 29883 28617
rect 29825 28608 29837 28611
rect 29512 28580 29837 28608
rect 29512 28568 29518 28580
rect 29825 28577 29837 28580
rect 29871 28577 29883 28611
rect 29825 28571 29883 28577
rect 30282 28568 30288 28620
rect 30340 28608 30346 28620
rect 31021 28611 31079 28617
rect 31021 28608 31033 28611
rect 30340 28580 31033 28608
rect 30340 28568 30346 28580
rect 31021 28577 31033 28580
rect 31067 28577 31079 28611
rect 31021 28571 31079 28577
rect 21913 28543 21971 28549
rect 21913 28509 21925 28543
rect 21959 28509 21971 28543
rect 22646 28540 22652 28552
rect 22607 28512 22652 28540
rect 21913 28503 21971 28509
rect 21560 28444 21772 28472
rect 20717 28435 20775 28441
rect 16761 28407 16819 28413
rect 16761 28373 16773 28407
rect 16807 28404 16819 28407
rect 17586 28404 17592 28416
rect 16807 28376 17592 28404
rect 16807 28373 16819 28376
rect 16761 28367 16819 28373
rect 17586 28364 17592 28376
rect 17644 28364 17650 28416
rect 17770 28404 17776 28416
rect 17731 28376 17776 28404
rect 17770 28364 17776 28376
rect 17828 28364 17834 28416
rect 19978 28364 19984 28416
rect 20036 28404 20042 28416
rect 20640 28404 20668 28435
rect 20036 28376 20668 28404
rect 20732 28404 20760 28435
rect 21634 28404 21640 28416
rect 20732 28376 21640 28404
rect 20036 28364 20042 28376
rect 21634 28364 21640 28376
rect 21692 28364 21698 28416
rect 21928 28404 21956 28503
rect 22646 28500 22652 28512
rect 22704 28500 22710 28552
rect 22830 28540 22836 28552
rect 22791 28512 22836 28540
rect 22830 28500 22836 28512
rect 22888 28500 22894 28552
rect 23014 28500 23020 28552
rect 23072 28540 23078 28552
rect 23072 28512 23117 28540
rect 23072 28500 23078 28512
rect 23198 28500 23204 28552
rect 23256 28540 23262 28552
rect 31128 28549 31156 28648
rect 36170 28608 36176 28620
rect 32784 28580 36176 28608
rect 30009 28543 30067 28549
rect 23256 28512 23301 28540
rect 23256 28500 23262 28512
rect 30009 28509 30021 28543
rect 30055 28540 30067 28543
rect 30837 28543 30895 28549
rect 30837 28540 30849 28543
rect 30055 28512 30849 28540
rect 30055 28509 30067 28512
rect 30009 28503 30067 28509
rect 30837 28509 30849 28512
rect 30883 28509 30895 28543
rect 30837 28503 30895 28509
rect 31113 28543 31171 28549
rect 31113 28509 31125 28543
rect 31159 28540 31171 28543
rect 31662 28540 31668 28552
rect 31159 28512 31668 28540
rect 31159 28509 31171 28512
rect 31113 28503 31171 28509
rect 29730 28472 29736 28484
rect 29691 28444 29736 28472
rect 29730 28432 29736 28444
rect 29788 28432 29794 28484
rect 30852 28472 30880 28503
rect 31662 28500 31668 28512
rect 31720 28500 31726 28552
rect 32784 28549 32812 28580
rect 36170 28568 36176 28580
rect 36228 28568 36234 28620
rect 32769 28543 32827 28549
rect 32769 28509 32781 28543
rect 32815 28509 32827 28543
rect 32769 28503 32827 28509
rect 33686 28500 33692 28552
rect 33744 28540 33750 28552
rect 34701 28543 34759 28549
rect 34701 28540 34713 28543
rect 33744 28512 34713 28540
rect 33744 28500 33750 28512
rect 34701 28509 34713 28512
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 46934 28500 46940 28552
rect 46992 28540 46998 28552
rect 47673 28543 47731 28549
rect 47673 28540 47685 28543
rect 46992 28512 47685 28540
rect 46992 28500 46998 28512
rect 47673 28509 47685 28512
rect 47719 28509 47731 28543
rect 47673 28503 47731 28509
rect 32398 28472 32404 28484
rect 30852 28444 32404 28472
rect 32398 28432 32404 28444
rect 32456 28432 32462 28484
rect 34974 28472 34980 28484
rect 34935 28444 34980 28472
rect 34974 28432 34980 28444
rect 35032 28432 35038 28484
rect 35434 28432 35440 28484
rect 35492 28432 35498 28484
rect 23842 28404 23848 28416
rect 21928 28376 23848 28404
rect 23842 28364 23848 28376
rect 23900 28364 23906 28416
rect 28994 28364 29000 28416
rect 29052 28404 29058 28416
rect 29362 28404 29368 28416
rect 29052 28376 29368 28404
rect 29052 28364 29058 28376
rect 29362 28364 29368 28376
rect 29420 28364 29426 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1486 28160 1492 28212
rect 1544 28200 1550 28212
rect 1544 28172 6914 28200
rect 1544 28160 1550 28172
rect 6886 28132 6914 28172
rect 20346 28160 20352 28212
rect 20404 28200 20410 28212
rect 20441 28203 20499 28209
rect 20441 28200 20453 28203
rect 20404 28172 20453 28200
rect 20404 28160 20410 28172
rect 20441 28169 20453 28172
rect 20487 28169 20499 28203
rect 24489 28203 24547 28209
rect 24489 28200 24501 28203
rect 20441 28163 20499 28169
rect 23584 28172 24501 28200
rect 6886 28104 22094 28132
rect 17586 28064 17592 28076
rect 17547 28036 17592 28064
rect 17586 28024 17592 28036
rect 17644 28024 17650 28076
rect 17770 28073 17776 28076
rect 17737 28067 17776 28073
rect 17737 28033 17749 28067
rect 17737 28027 17776 28033
rect 17770 28024 17776 28027
rect 17828 28024 17834 28076
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28033 17923 28067
rect 17865 28027 17923 28033
rect 17880 27996 17908 28027
rect 17954 28024 17960 28076
rect 18012 28064 18018 28076
rect 18095 28067 18153 28073
rect 18012 28036 18057 28064
rect 18012 28024 18018 28036
rect 18095 28033 18107 28067
rect 18141 28064 18153 28067
rect 18230 28064 18236 28076
rect 18141 28036 18236 28064
rect 18141 28033 18153 28036
rect 18095 28027 18153 28033
rect 18230 28024 18236 28036
rect 18288 28024 18294 28076
rect 20070 28064 20076 28076
rect 20031 28036 20076 28064
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28064 20315 28067
rect 20438 28064 20444 28076
rect 20303 28036 20444 28064
rect 20303 28033 20315 28036
rect 20257 28027 20315 28033
rect 20438 28024 20444 28036
rect 20496 28024 20502 28076
rect 21634 28024 21640 28076
rect 21692 28064 21698 28076
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21692 28036 21833 28064
rect 21692 28024 21698 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 21910 28024 21916 28076
rect 21968 28064 21974 28076
rect 21968 28036 22013 28064
rect 21968 28024 21974 28036
rect 19978 27996 19984 28008
rect 17880 27968 19984 27996
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 20088 27928 20116 28024
rect 22066 27996 22094 28104
rect 23584 28073 23612 28172
rect 24489 28169 24501 28172
rect 24535 28200 24547 28203
rect 24670 28200 24676 28212
rect 24535 28172 24676 28200
rect 24535 28169 24547 28172
rect 24489 28163 24547 28169
rect 24670 28160 24676 28172
rect 24728 28160 24734 28212
rect 26329 28203 26387 28209
rect 26329 28169 26341 28203
rect 26375 28200 26387 28203
rect 26510 28200 26516 28212
rect 26375 28172 26516 28200
rect 26375 28169 26387 28172
rect 26329 28163 26387 28169
rect 26510 28160 26516 28172
rect 26568 28160 26574 28212
rect 26973 28203 27031 28209
rect 26973 28169 26985 28203
rect 27019 28169 27031 28203
rect 26973 28163 27031 28169
rect 28353 28203 28411 28209
rect 28353 28169 28365 28203
rect 28399 28200 28411 28203
rect 28994 28200 29000 28212
rect 28399 28172 29000 28200
rect 28399 28169 28411 28172
rect 28353 28163 28411 28169
rect 24397 28135 24455 28141
rect 24397 28101 24409 28135
rect 24443 28132 24455 28135
rect 25038 28132 25044 28144
rect 24443 28104 25044 28132
rect 24443 28101 24455 28104
rect 24397 28095 24455 28101
rect 25038 28092 25044 28104
rect 25096 28092 25102 28144
rect 26988 28132 27016 28163
rect 28994 28160 29000 28172
rect 29052 28160 29058 28212
rect 29362 28160 29368 28212
rect 29420 28200 29426 28212
rect 29420 28172 29500 28200
rect 29420 28160 29426 28172
rect 29472 28141 29500 28172
rect 29638 28160 29644 28212
rect 29696 28160 29702 28212
rect 33686 28200 33692 28212
rect 33647 28172 33692 28200
rect 33686 28160 33692 28172
rect 33744 28160 33750 28212
rect 35345 28203 35403 28209
rect 35345 28169 35357 28203
rect 35391 28200 35403 28203
rect 35434 28200 35440 28212
rect 35391 28172 35440 28200
rect 35391 28169 35403 28172
rect 35345 28163 35403 28169
rect 35434 28160 35440 28172
rect 35492 28160 35498 28212
rect 42794 28160 42800 28212
rect 42852 28200 42858 28212
rect 46842 28200 46848 28212
rect 42852 28172 46848 28200
rect 42852 28160 42858 28172
rect 46842 28160 46848 28172
rect 46900 28160 46906 28212
rect 26160 28104 27016 28132
rect 29457 28135 29515 28141
rect 23569 28067 23627 28073
rect 23569 28033 23581 28067
rect 23615 28064 23627 28067
rect 23658 28064 23664 28076
rect 23615 28036 23664 28064
rect 23615 28033 23627 28036
rect 23569 28027 23627 28033
rect 23658 28024 23664 28036
rect 23716 28024 23722 28076
rect 26160 28073 26188 28104
rect 29457 28101 29469 28135
rect 29503 28101 29515 28135
rect 29457 28095 29515 28101
rect 29549 28135 29607 28141
rect 29549 28101 29561 28135
rect 29595 28132 29607 28135
rect 29656 28132 29684 28160
rect 29595 28104 29684 28132
rect 29595 28101 29607 28104
rect 29549 28095 29607 28101
rect 26145 28067 26203 28073
rect 26145 28033 26157 28067
rect 26191 28033 26203 28067
rect 26145 28027 26203 28033
rect 26421 28067 26479 28073
rect 26421 28033 26433 28067
rect 26467 28033 26479 28067
rect 27341 28067 27399 28073
rect 27341 28064 27353 28067
rect 26421 28027 26479 28033
rect 26528 28036 27353 28064
rect 26436 27996 26464 28027
rect 22066 27968 26464 27996
rect 20088 27900 23152 27928
rect 18230 27860 18236 27872
rect 18191 27832 18236 27860
rect 18230 27820 18236 27832
rect 18288 27820 18294 27872
rect 21818 27860 21824 27872
rect 21779 27832 21824 27860
rect 21818 27820 21824 27832
rect 21876 27820 21882 27872
rect 21910 27820 21916 27872
rect 21968 27860 21974 27872
rect 22189 27863 22247 27869
rect 22189 27860 22201 27863
rect 21968 27832 22201 27860
rect 21968 27820 21974 27832
rect 22189 27829 22201 27832
rect 22235 27829 22247 27863
rect 23124 27860 23152 27900
rect 23198 27888 23204 27940
rect 23256 27928 23262 27940
rect 23753 27931 23811 27937
rect 23753 27928 23765 27931
rect 23256 27900 23765 27928
rect 23256 27888 23262 27900
rect 23753 27897 23765 27900
rect 23799 27897 23811 27931
rect 23753 27891 23811 27897
rect 24578 27888 24584 27940
rect 24636 27928 24642 27940
rect 26528 27928 26556 28036
rect 27341 28033 27353 28036
rect 27387 28033 27399 28067
rect 28169 28067 28227 28073
rect 28169 28064 28181 28067
rect 27341 28027 27399 28033
rect 27448 28036 28181 28064
rect 26602 27956 26608 28008
rect 26660 27996 26666 28008
rect 27448 28005 27476 28036
rect 28169 28033 28181 28036
rect 28215 28033 28227 28067
rect 28169 28027 28227 28033
rect 29273 28067 29331 28073
rect 29273 28033 29285 28067
rect 29319 28033 29331 28067
rect 29273 28027 29331 28033
rect 29641 28070 29699 28073
rect 29641 28067 29708 28070
rect 29641 28033 29653 28067
rect 29687 28064 29708 28067
rect 30469 28067 30527 28073
rect 29687 28036 29776 28064
rect 29687 28033 29699 28036
rect 29641 28027 29699 28033
rect 27433 27999 27491 28005
rect 27433 27996 27445 27999
rect 26660 27968 27445 27996
rect 26660 27956 26666 27968
rect 27433 27965 27445 27968
rect 27479 27965 27491 27999
rect 27433 27959 27491 27965
rect 27525 27999 27583 28005
rect 27525 27965 27537 27999
rect 27571 27996 27583 27999
rect 28074 27996 28080 28008
rect 27571 27968 28080 27996
rect 27571 27965 27583 27968
rect 27525 27959 27583 27965
rect 28074 27956 28080 27968
rect 28132 27956 28138 28008
rect 29288 27996 29316 28027
rect 29546 27996 29552 28008
rect 29288 27968 29552 27996
rect 29546 27956 29552 27968
rect 29604 27956 29610 28008
rect 24636 27900 26556 27928
rect 24636 27888 24642 27900
rect 29362 27888 29368 27940
rect 29420 27928 29426 27940
rect 29748 27928 29776 28036
rect 30469 28033 30481 28067
rect 30515 28064 30527 28067
rect 31662 28064 31668 28076
rect 30515 28036 31668 28064
rect 30515 28033 30527 28036
rect 30469 28027 30527 28033
rect 31662 28024 31668 28036
rect 31720 28024 31726 28076
rect 32490 28024 32496 28076
rect 32548 28064 32554 28076
rect 33597 28067 33655 28073
rect 33597 28064 33609 28067
rect 32548 28036 33609 28064
rect 32548 28024 32554 28036
rect 33597 28033 33609 28036
rect 33643 28033 33655 28067
rect 33597 28027 33655 28033
rect 34330 28024 34336 28076
rect 34388 28064 34394 28076
rect 34425 28067 34483 28073
rect 34425 28064 34437 28067
rect 34388 28036 34437 28064
rect 34388 28024 34394 28036
rect 34425 28033 34437 28036
rect 34471 28033 34483 28067
rect 34425 28027 34483 28033
rect 35253 28067 35311 28073
rect 35253 28033 35265 28067
rect 35299 28064 35311 28067
rect 35526 28064 35532 28076
rect 35299 28036 35532 28064
rect 35299 28033 35311 28036
rect 35253 28027 35311 28033
rect 35526 28024 35532 28036
rect 35584 28024 35590 28076
rect 47026 28024 47032 28076
rect 47084 28064 47090 28076
rect 47394 28064 47400 28076
rect 47084 28036 47400 28064
rect 47084 28024 47090 28036
rect 47394 28024 47400 28036
rect 47452 28064 47458 28076
rect 47581 28067 47639 28073
rect 47581 28064 47593 28067
rect 47452 28036 47593 28064
rect 47452 28024 47458 28036
rect 47581 28033 47593 28036
rect 47627 28033 47639 28067
rect 47581 28027 47639 28033
rect 30282 27956 30288 28008
rect 30340 27996 30346 28008
rect 30377 27999 30435 28005
rect 30377 27996 30389 27999
rect 30340 27968 30389 27996
rect 30340 27956 30346 27968
rect 30377 27965 30389 27968
rect 30423 27965 30435 27999
rect 30377 27959 30435 27965
rect 34517 27999 34575 28005
rect 34517 27965 34529 27999
rect 34563 27996 34575 27999
rect 34698 27996 34704 28008
rect 34563 27968 34704 27996
rect 34563 27965 34575 27968
rect 34517 27959 34575 27965
rect 34698 27956 34704 27968
rect 34756 27956 34762 28008
rect 34793 27999 34851 28005
rect 34793 27965 34805 27999
rect 34839 27996 34851 27999
rect 34974 27996 34980 28008
rect 34839 27968 34980 27996
rect 34839 27965 34851 27968
rect 34793 27959 34851 27965
rect 34974 27956 34980 27968
rect 35032 27956 35038 28008
rect 29420 27900 29776 27928
rect 29420 27888 29426 27900
rect 25130 27860 25136 27872
rect 23124 27832 25136 27860
rect 22189 27823 22247 27829
rect 25130 27820 25136 27832
rect 25188 27820 25194 27872
rect 25961 27863 26019 27869
rect 25961 27829 25973 27863
rect 26007 27860 26019 27863
rect 26878 27860 26884 27872
rect 26007 27832 26884 27860
rect 26007 27829 26019 27832
rect 25961 27823 26019 27829
rect 26878 27820 26884 27832
rect 26936 27820 26942 27872
rect 29825 27863 29883 27869
rect 29825 27829 29837 27863
rect 29871 27860 29883 27863
rect 30374 27860 30380 27872
rect 29871 27832 30380 27860
rect 29871 27829 29883 27832
rect 29825 27823 29883 27829
rect 30374 27820 30380 27832
rect 30432 27820 30438 27872
rect 30742 27860 30748 27872
rect 30703 27832 30748 27860
rect 30742 27820 30748 27832
rect 30800 27820 30806 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 3510 27616 3516 27668
rect 3568 27656 3574 27668
rect 31662 27656 31668 27668
rect 3568 27628 14688 27656
rect 31623 27628 31668 27656
rect 3568 27616 3574 27628
rect 7466 27480 7472 27532
rect 7524 27520 7530 27532
rect 14660 27520 14688 27628
rect 31662 27616 31668 27628
rect 31720 27616 31726 27668
rect 15102 27548 15108 27600
rect 15160 27588 15166 27600
rect 17862 27588 17868 27600
rect 15160 27560 17868 27588
rect 15160 27548 15166 27560
rect 17862 27548 17868 27560
rect 17920 27548 17926 27600
rect 22830 27588 22836 27600
rect 20088 27560 22836 27588
rect 15565 27523 15623 27529
rect 15565 27520 15577 27523
rect 7524 27492 12434 27520
rect 14660 27492 15577 27520
rect 7524 27480 7530 27492
rect 12406 27316 12434 27492
rect 15565 27489 15577 27492
rect 15611 27489 15623 27523
rect 15565 27483 15623 27489
rect 15102 27452 15108 27464
rect 15063 27424 15108 27452
rect 15102 27412 15108 27424
rect 15160 27412 15166 27464
rect 19889 27455 19947 27461
rect 19889 27421 19901 27455
rect 19935 27452 19947 27455
rect 19978 27452 19984 27464
rect 19935 27424 19984 27452
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 19978 27412 19984 27424
rect 20036 27412 20042 27464
rect 20088 27461 20116 27560
rect 22830 27548 22836 27560
rect 22888 27548 22894 27600
rect 26050 27548 26056 27600
rect 26108 27588 26114 27600
rect 26605 27591 26663 27597
rect 26605 27588 26617 27591
rect 26108 27560 26617 27588
rect 26108 27548 26114 27560
rect 26605 27557 26617 27560
rect 26651 27557 26663 27591
rect 29454 27588 29460 27600
rect 26605 27551 26663 27557
rect 28276 27560 29460 27588
rect 20165 27523 20223 27529
rect 20165 27489 20177 27523
rect 20211 27520 20223 27523
rect 23198 27520 23204 27532
rect 20211 27492 20392 27520
rect 20211 27489 20223 27492
rect 20165 27483 20223 27489
rect 20073 27455 20131 27461
rect 20073 27421 20085 27455
rect 20119 27421 20131 27455
rect 20073 27415 20131 27421
rect 20257 27455 20315 27461
rect 20257 27421 20269 27455
rect 20303 27421 20315 27455
rect 20257 27415 20315 27421
rect 15289 27387 15347 27393
rect 15289 27353 15301 27387
rect 15335 27384 15347 27387
rect 15378 27384 15384 27396
rect 15335 27356 15384 27384
rect 15335 27353 15347 27356
rect 15289 27347 15347 27353
rect 15378 27344 15384 27356
rect 15436 27344 15442 27396
rect 20272 27316 20300 27415
rect 20364 27384 20392 27492
rect 20456 27492 23204 27520
rect 20456 27461 20484 27492
rect 23198 27480 23204 27492
rect 23256 27480 23262 27532
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27421 20499 27455
rect 21082 27452 21088 27464
rect 21043 27424 21088 27452
rect 20441 27415 20499 27421
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 21266 27452 21272 27464
rect 21227 27424 21272 27452
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 24489 27455 24547 27461
rect 24489 27421 24501 27455
rect 24535 27421 24547 27455
rect 24489 27415 24547 27421
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27452 24639 27455
rect 25038 27452 25044 27464
rect 24627 27424 25044 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 20806 27384 20812 27396
rect 20364 27356 20812 27384
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 23842 27344 23848 27396
rect 23900 27384 23906 27396
rect 24504 27384 24532 27415
rect 25038 27412 25044 27424
rect 25096 27412 25102 27464
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27452 27491 27455
rect 27890 27452 27896 27464
rect 27479 27424 27896 27452
rect 27479 27421 27491 27424
rect 27433 27415 27491 27421
rect 27890 27412 27896 27424
rect 27948 27412 27954 27464
rect 28074 27452 28080 27464
rect 28035 27424 28080 27452
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28276 27461 28304 27560
rect 29454 27548 29460 27560
rect 29512 27548 29518 27600
rect 46934 27588 46940 27600
rect 46308 27560 46940 27588
rect 29822 27480 29828 27532
rect 29880 27520 29886 27532
rect 46308 27529 46336 27560
rect 46934 27548 46940 27560
rect 46992 27548 46998 27600
rect 29917 27523 29975 27529
rect 29917 27520 29929 27523
rect 29880 27492 29929 27520
rect 29880 27480 29886 27492
rect 29917 27489 29929 27492
rect 29963 27489 29975 27523
rect 29917 27483 29975 27489
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46293 27483 46351 27489
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 47670 27520 47676 27532
rect 46523 27492 47676 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 47670 27480 47676 27492
rect 47728 27480 47734 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 28261 27455 28319 27461
rect 28261 27421 28273 27455
rect 28307 27421 28319 27455
rect 28997 27455 29055 27461
rect 28997 27452 29009 27455
rect 28261 27415 28319 27421
rect 28552 27424 29009 27452
rect 25222 27384 25228 27396
rect 23900 27356 25228 27384
rect 23900 27344 23906 27356
rect 25222 27344 25228 27356
rect 25280 27344 25286 27396
rect 26421 27387 26479 27393
rect 26421 27353 26433 27387
rect 26467 27384 26479 27387
rect 26602 27384 26608 27396
rect 26467 27356 26608 27384
rect 26467 27353 26479 27356
rect 26421 27347 26479 27353
rect 26602 27344 26608 27356
rect 26660 27344 26666 27396
rect 28169 27387 28227 27393
rect 28169 27353 28181 27387
rect 28215 27384 28227 27387
rect 28552 27384 28580 27424
rect 28997 27421 29009 27424
rect 29043 27421 29055 27455
rect 32490 27452 32496 27464
rect 32451 27424 32496 27452
rect 28997 27415 29055 27421
rect 32490 27412 32496 27424
rect 32548 27412 32554 27464
rect 33321 27455 33379 27461
rect 33321 27421 33333 27455
rect 33367 27452 33379 27455
rect 35526 27452 35532 27464
rect 33367 27424 35532 27452
rect 33367 27421 33379 27424
rect 33321 27415 33379 27421
rect 35526 27412 35532 27424
rect 35584 27412 35590 27464
rect 28721 27387 28779 27393
rect 28721 27384 28733 27387
rect 28215 27356 28580 27384
rect 28644 27356 28733 27384
rect 28215 27353 28227 27356
rect 28169 27347 28227 27353
rect 20622 27316 20628 27328
rect 12406 27288 20300 27316
rect 20583 27288 20628 27316
rect 20622 27276 20628 27288
rect 20680 27276 20686 27328
rect 21174 27316 21180 27328
rect 21135 27288 21180 27316
rect 21174 27276 21180 27288
rect 21232 27276 21238 27328
rect 24762 27316 24768 27328
rect 24723 27288 24768 27316
rect 24762 27276 24768 27288
rect 24820 27276 24826 27328
rect 27522 27316 27528 27328
rect 27483 27288 27528 27316
rect 27522 27276 27528 27288
rect 27580 27276 27586 27328
rect 27982 27276 27988 27328
rect 28040 27316 28046 27328
rect 28644 27316 28672 27356
rect 28721 27353 28733 27356
rect 28767 27353 28779 27387
rect 30190 27384 30196 27396
rect 30151 27356 30196 27384
rect 28721 27347 28779 27353
rect 30190 27344 30196 27356
rect 30248 27344 30254 27396
rect 31202 27344 31208 27396
rect 31260 27344 31266 27396
rect 28810 27316 28816 27328
rect 28868 27325 28874 27328
rect 28040 27288 28672 27316
rect 28777 27288 28816 27316
rect 28040 27276 28046 27288
rect 28810 27276 28816 27288
rect 28868 27279 28877 27325
rect 28905 27319 28963 27325
rect 28905 27285 28917 27319
rect 28951 27316 28963 27319
rect 30282 27316 30288 27328
rect 28951 27288 30288 27316
rect 28951 27285 28963 27288
rect 28905 27279 28963 27285
rect 28868 27276 28874 27279
rect 30282 27276 30288 27288
rect 30340 27276 30346 27328
rect 32306 27276 32312 27328
rect 32364 27316 32370 27328
rect 32493 27319 32551 27325
rect 32493 27316 32505 27319
rect 32364 27288 32505 27316
rect 32364 27276 32370 27288
rect 32493 27285 32505 27288
rect 32539 27285 32551 27319
rect 32493 27279 32551 27285
rect 33318 27276 33324 27328
rect 33376 27316 33382 27328
rect 33413 27319 33471 27325
rect 33413 27316 33425 27319
rect 33376 27288 33425 27316
rect 33376 27276 33382 27288
rect 33413 27285 33425 27288
rect 33459 27285 33471 27319
rect 33413 27279 33471 27285
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 15378 27112 15384 27124
rect 15339 27084 15384 27112
rect 15378 27072 15384 27084
rect 15436 27072 15442 27124
rect 22002 27072 22008 27124
rect 22060 27112 22066 27124
rect 22060 27072 22094 27112
rect 28074 27072 28080 27124
rect 28132 27112 28138 27124
rect 28721 27115 28779 27121
rect 28721 27112 28733 27115
rect 28132 27084 28733 27112
rect 28132 27072 28138 27084
rect 28721 27081 28733 27084
rect 28767 27081 28779 27115
rect 30190 27112 30196 27124
rect 30151 27084 30196 27112
rect 28721 27075 28779 27081
rect 21821 27047 21879 27053
rect 19904 27016 20852 27044
rect 15289 26979 15347 26985
rect 15289 26945 15301 26979
rect 15335 26976 15347 26979
rect 15470 26976 15476 26988
rect 15335 26948 15476 26976
rect 15335 26945 15347 26948
rect 15289 26939 15347 26945
rect 15470 26936 15476 26948
rect 15528 26976 15534 26988
rect 15933 26979 15991 26985
rect 15933 26976 15945 26979
rect 15528 26948 15945 26976
rect 15528 26936 15534 26948
rect 15933 26945 15945 26948
rect 15979 26945 15991 26979
rect 15933 26939 15991 26945
rect 18598 26936 18604 26988
rect 18656 26936 18662 26988
rect 19904 26985 19932 27016
rect 20824 26988 20852 27016
rect 21821 27013 21833 27047
rect 21867 27044 21879 27047
rect 21910 27044 21916 27056
rect 21867 27016 21916 27044
rect 21867 27013 21879 27016
rect 21821 27007 21879 27013
rect 21910 27004 21916 27016
rect 21968 27004 21974 27056
rect 22066 27044 22094 27072
rect 22833 27047 22891 27053
rect 22833 27044 22845 27047
rect 22066 27016 22845 27044
rect 22833 27013 22845 27016
rect 22879 27013 22891 27047
rect 27246 27044 27252 27056
rect 22833 27007 22891 27013
rect 23768 27016 24624 27044
rect 23768 26988 23796 27016
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26945 19947 26979
rect 20625 26979 20683 26985
rect 20625 26976 20637 26979
rect 19889 26939 19947 26945
rect 20180 26948 20637 26976
rect 17218 26908 17224 26920
rect 17179 26880 17224 26908
rect 17218 26868 17224 26880
rect 17276 26868 17282 26920
rect 17497 26911 17555 26917
rect 17497 26877 17509 26911
rect 17543 26908 17555 26911
rect 18230 26908 18236 26920
rect 17543 26880 18236 26908
rect 17543 26877 17555 26880
rect 17497 26871 17555 26877
rect 18230 26868 18236 26880
rect 18288 26868 18294 26920
rect 19705 26911 19763 26917
rect 19705 26877 19717 26911
rect 19751 26908 19763 26911
rect 20070 26908 20076 26920
rect 19751 26880 20076 26908
rect 19751 26877 19763 26880
rect 19705 26871 19763 26877
rect 20070 26868 20076 26880
rect 20128 26868 20134 26920
rect 20180 26917 20208 26948
rect 20625 26945 20637 26948
rect 20671 26945 20683 26979
rect 20806 26976 20812 26988
rect 20767 26948 20812 26976
rect 20625 26939 20683 26945
rect 20806 26936 20812 26948
rect 20864 26936 20870 26988
rect 21542 26936 21548 26988
rect 21600 26976 21606 26988
rect 21726 26976 21732 26988
rect 21600 26948 21732 26976
rect 21600 26936 21606 26948
rect 21726 26936 21732 26948
rect 21784 26976 21790 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21784 26948 22017 26976
rect 21784 26936 21790 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 22649 26979 22707 26985
rect 22649 26945 22661 26979
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 23661 26979 23719 26985
rect 23661 26945 23673 26979
rect 23707 26976 23719 26979
rect 23750 26976 23756 26988
rect 23707 26948 23756 26976
rect 23707 26945 23719 26948
rect 23661 26939 23719 26945
rect 20165 26911 20223 26917
rect 20165 26877 20177 26911
rect 20211 26877 20223 26911
rect 20165 26871 20223 26877
rect 20993 26911 21051 26917
rect 20993 26877 21005 26911
rect 21039 26908 21051 26911
rect 21082 26908 21088 26920
rect 21039 26880 21088 26908
rect 21039 26877 21051 26880
rect 20993 26871 21051 26877
rect 20180 26840 20208 26871
rect 21082 26868 21088 26880
rect 21140 26908 21146 26920
rect 21634 26908 21640 26920
rect 21140 26880 21640 26908
rect 21140 26868 21146 26880
rect 21634 26868 21640 26880
rect 21692 26908 21698 26920
rect 22664 26908 22692 26939
rect 23750 26936 23756 26948
rect 23808 26936 23814 26988
rect 23842 26936 23848 26988
rect 23900 26976 23906 26988
rect 24596 26985 24624 27016
rect 26988 27016 27252 27044
rect 26988 26985 27016 27016
rect 27246 27004 27252 27016
rect 27304 27004 27310 27056
rect 27522 27004 27528 27056
rect 27580 27044 27586 27056
rect 28736 27044 28764 27075
rect 30190 27072 30196 27084
rect 30248 27072 30254 27124
rect 31202 27112 31208 27124
rect 31163 27084 31208 27112
rect 31202 27072 31208 27084
rect 31260 27072 31266 27124
rect 32674 27072 32680 27124
rect 32732 27112 32738 27124
rect 34057 27115 34115 27121
rect 34057 27112 34069 27115
rect 32732 27084 34069 27112
rect 32732 27072 32738 27084
rect 34057 27081 34069 27084
rect 34103 27112 34115 27115
rect 34330 27112 34336 27124
rect 34103 27084 34336 27112
rect 34103 27081 34115 27084
rect 34057 27075 34115 27081
rect 34330 27072 34336 27084
rect 34388 27072 34394 27124
rect 35802 27112 35808 27124
rect 34532 27084 35808 27112
rect 29273 27047 29331 27053
rect 29273 27044 29285 27047
rect 27580 27016 27738 27044
rect 28736 27016 29285 27044
rect 27580 27004 27586 27016
rect 29273 27013 29285 27016
rect 29319 27044 29331 27047
rect 29730 27044 29736 27056
rect 29319 27016 29736 27044
rect 29319 27013 29331 27016
rect 29273 27007 29331 27013
rect 29730 27004 29736 27016
rect 29788 27004 29794 27056
rect 30561 27047 30619 27053
rect 30561 27013 30573 27047
rect 30607 27044 30619 27047
rect 31386 27044 31392 27056
rect 30607 27016 31392 27044
rect 30607 27013 30619 27016
rect 30561 27007 30619 27013
rect 31386 27004 31392 27016
rect 31444 27004 31450 27056
rect 33318 27004 33324 27056
rect 33376 27004 33382 27056
rect 33962 27004 33968 27056
rect 34020 27044 34026 27056
rect 34532 27053 34560 27084
rect 35802 27072 35808 27084
rect 35860 27072 35866 27124
rect 34517 27047 34575 27053
rect 34517 27044 34529 27047
rect 34020 27016 34529 27044
rect 34020 27004 34026 27016
rect 34517 27013 34529 27016
rect 34563 27013 34575 27047
rect 34517 27007 34575 27013
rect 34606 27004 34612 27056
rect 34664 27044 34670 27056
rect 34717 27047 34775 27053
rect 34717 27044 34729 27047
rect 34664 27016 34729 27044
rect 34664 27004 34670 27016
rect 34717 27013 34729 27016
rect 34763 27013 34775 27047
rect 34717 27007 34775 27013
rect 24489 26979 24547 26985
rect 23900 26948 23945 26976
rect 23900 26936 23906 26948
rect 24489 26945 24501 26979
rect 24535 26945 24547 26979
rect 24489 26939 24547 26945
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26945 24639 26979
rect 24581 26939 24639 26945
rect 26973 26979 27031 26985
rect 26973 26945 26985 26979
rect 27019 26945 27031 26979
rect 29454 26976 29460 26988
rect 29415 26948 29460 26976
rect 26973 26939 27031 26945
rect 21692 26880 22692 26908
rect 23017 26911 23075 26917
rect 21692 26868 21698 26880
rect 23017 26877 23029 26911
rect 23063 26908 23075 26911
rect 23382 26908 23388 26920
rect 23063 26880 23388 26908
rect 23063 26877 23075 26880
rect 23017 26871 23075 26877
rect 23382 26868 23388 26880
rect 23440 26908 23446 26920
rect 24504 26908 24532 26939
rect 29454 26936 29460 26948
rect 29512 26936 29518 26988
rect 30374 26976 30380 26988
rect 30335 26948 30380 26976
rect 30374 26936 30380 26948
rect 30432 26936 30438 26988
rect 30653 26979 30711 26985
rect 30653 26945 30665 26979
rect 30699 26976 30711 26979
rect 30742 26976 30748 26988
rect 30699 26948 30748 26976
rect 30699 26945 30711 26948
rect 30653 26939 30711 26945
rect 30742 26936 30748 26948
rect 30800 26936 30806 26988
rect 31113 26979 31171 26985
rect 31113 26945 31125 26979
rect 31159 26945 31171 26979
rect 32306 26976 32312 26988
rect 32267 26948 32312 26976
rect 31113 26939 31171 26945
rect 23440 26880 24532 26908
rect 23440 26868 23446 26880
rect 24854 26868 24860 26920
rect 24912 26868 24918 26920
rect 26878 26868 26884 26920
rect 26936 26908 26942 26920
rect 27249 26911 27307 26917
rect 27249 26908 27261 26911
rect 26936 26880 27261 26908
rect 26936 26868 26942 26880
rect 27249 26877 27261 26880
rect 27295 26877 27307 26911
rect 27249 26871 27307 26877
rect 29641 26911 29699 26917
rect 29641 26877 29653 26911
rect 29687 26908 29699 26911
rect 30282 26908 30288 26920
rect 29687 26880 30288 26908
rect 29687 26877 29699 26880
rect 29641 26871 29699 26877
rect 30282 26868 30288 26880
rect 30340 26868 30346 26920
rect 18984 26812 20208 26840
rect 15010 26732 15016 26784
rect 15068 26772 15074 26784
rect 16025 26775 16083 26781
rect 16025 26772 16037 26775
rect 15068 26744 16037 26772
rect 15068 26732 15074 26744
rect 16025 26741 16037 26744
rect 16071 26741 16083 26775
rect 16025 26735 16083 26741
rect 17954 26732 17960 26784
rect 18012 26772 18018 26784
rect 18984 26781 19012 26812
rect 21542 26800 21548 26852
rect 21600 26840 21606 26852
rect 24029 26843 24087 26849
rect 24029 26840 24041 26843
rect 21600 26812 24041 26840
rect 21600 26800 21606 26812
rect 24029 26809 24041 26812
rect 24075 26809 24087 26843
rect 24872 26840 24900 26868
rect 24029 26803 24087 26809
rect 24688 26812 24900 26840
rect 18969 26775 19027 26781
rect 18969 26772 18981 26775
rect 18012 26744 18981 26772
rect 18012 26732 18018 26744
rect 18969 26741 18981 26744
rect 19015 26741 19027 26775
rect 18969 26735 19027 26741
rect 20073 26775 20131 26781
rect 20073 26741 20085 26775
rect 20119 26772 20131 26775
rect 21266 26772 21272 26784
rect 20119 26744 21272 26772
rect 20119 26741 20131 26744
rect 20073 26735 20131 26741
rect 21266 26732 21272 26744
rect 21324 26772 21330 26784
rect 22002 26772 22008 26784
rect 21324 26744 22008 26772
rect 21324 26732 21330 26744
rect 22002 26732 22008 26744
rect 22060 26772 22066 26784
rect 22097 26775 22155 26781
rect 22097 26772 22109 26775
rect 22060 26744 22109 26772
rect 22060 26732 22066 26744
rect 22097 26741 22109 26744
rect 22143 26741 22155 26775
rect 22097 26735 22155 26741
rect 23474 26732 23480 26784
rect 23532 26772 23538 26784
rect 24688 26781 24716 26812
rect 24673 26775 24731 26781
rect 24673 26772 24685 26775
rect 23532 26744 24685 26772
rect 23532 26732 23538 26744
rect 24673 26741 24685 26744
rect 24719 26741 24731 26775
rect 24854 26772 24860 26784
rect 24815 26744 24860 26772
rect 24673 26735 24731 26741
rect 24854 26732 24860 26744
rect 24912 26732 24918 26784
rect 27890 26732 27896 26784
rect 27948 26772 27954 26784
rect 31128 26772 31156 26939
rect 32306 26936 32312 26948
rect 32364 26936 32370 26988
rect 33870 26936 33876 26988
rect 33928 26976 33934 26988
rect 35345 26979 35403 26985
rect 35345 26976 35357 26979
rect 33928 26948 35357 26976
rect 33928 26936 33934 26948
rect 35345 26945 35357 26948
rect 35391 26945 35403 26979
rect 35345 26939 35403 26945
rect 35529 26979 35587 26985
rect 35529 26945 35541 26979
rect 35575 26945 35587 26979
rect 35529 26939 35587 26945
rect 32585 26911 32643 26917
rect 32585 26877 32597 26911
rect 32631 26908 32643 26911
rect 33134 26908 33140 26920
rect 32631 26880 33140 26908
rect 32631 26877 32643 26880
rect 32585 26871 32643 26877
rect 33134 26868 33140 26880
rect 33192 26868 33198 26920
rect 35544 26908 35572 26939
rect 34900 26880 35572 26908
rect 34606 26800 34612 26852
rect 34664 26840 34670 26852
rect 34900 26849 34928 26880
rect 34885 26843 34943 26849
rect 34885 26840 34897 26843
rect 34664 26812 34897 26840
rect 34664 26800 34670 26812
rect 34885 26809 34897 26812
rect 34931 26809 34943 26843
rect 34885 26803 34943 26809
rect 27948 26744 31156 26772
rect 34701 26775 34759 26781
rect 27948 26732 27954 26744
rect 34701 26741 34713 26775
rect 34747 26772 34759 26775
rect 34790 26772 34796 26784
rect 34747 26744 34796 26772
rect 34747 26741 34759 26744
rect 34701 26735 34759 26741
rect 34790 26732 34796 26744
rect 34848 26732 34854 26784
rect 35342 26772 35348 26784
rect 35303 26744 35348 26772
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 18598 26568 18604 26580
rect 18559 26540 18604 26568
rect 18598 26528 18604 26540
rect 18656 26528 18662 26580
rect 19508 26571 19566 26577
rect 19508 26537 19520 26571
rect 19554 26568 19566 26571
rect 20622 26568 20628 26580
rect 19554 26540 20628 26568
rect 19554 26537 19566 26540
rect 19508 26531 19566 26537
rect 20622 26528 20628 26540
rect 20680 26528 20686 26580
rect 20806 26528 20812 26580
rect 20864 26568 20870 26580
rect 20993 26571 21051 26577
rect 20993 26568 21005 26571
rect 20864 26540 21005 26568
rect 20864 26528 20870 26540
rect 20993 26537 21005 26540
rect 21039 26537 21051 26571
rect 20993 26531 21051 26537
rect 21821 26571 21879 26577
rect 21821 26537 21833 26571
rect 21867 26568 21879 26571
rect 21910 26568 21916 26580
rect 21867 26540 21916 26568
rect 21867 26537 21879 26540
rect 21821 26531 21879 26537
rect 21910 26528 21916 26540
rect 21968 26528 21974 26580
rect 23308 26540 24532 26568
rect 21174 26460 21180 26512
rect 21232 26500 21238 26512
rect 22005 26503 22063 26509
rect 21232 26472 21772 26500
rect 21232 26460 21238 26472
rect 15010 26432 15016 26444
rect 14971 26404 15016 26432
rect 15010 26392 15016 26404
rect 15068 26392 15074 26444
rect 16482 26432 16488 26444
rect 16443 26404 16488 26432
rect 16482 26392 16488 26404
rect 16540 26392 16546 26444
rect 17218 26392 17224 26444
rect 17276 26432 17282 26444
rect 19245 26435 19303 26441
rect 19245 26432 19257 26435
rect 17276 26404 19257 26432
rect 17276 26392 17282 26404
rect 19245 26401 19257 26404
rect 19291 26432 19303 26435
rect 21634 26432 21640 26444
rect 19291 26404 20944 26432
rect 21595 26404 21640 26432
rect 19291 26401 19303 26404
rect 19245 26395 19303 26401
rect 13722 26324 13728 26376
rect 13780 26364 13786 26376
rect 14829 26367 14887 26373
rect 14829 26364 14841 26367
rect 13780 26336 14841 26364
rect 13780 26324 13786 26336
rect 14829 26333 14841 26336
rect 14875 26333 14887 26367
rect 14829 26327 14887 26333
rect 18509 26367 18567 26373
rect 18509 26333 18521 26367
rect 18555 26364 18567 26367
rect 20916 26364 20944 26404
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 21744 26432 21772 26472
rect 22005 26469 22017 26503
rect 22051 26500 22063 26503
rect 22278 26500 22284 26512
rect 22051 26472 22284 26500
rect 22051 26469 22063 26472
rect 22005 26463 22063 26469
rect 22278 26460 22284 26472
rect 22336 26460 22342 26512
rect 23308 26432 23336 26540
rect 23382 26460 23388 26512
rect 23440 26500 23446 26512
rect 23440 26472 23612 26500
rect 23440 26460 23446 26472
rect 21744 26404 23336 26432
rect 21821 26367 21879 26373
rect 18555 26336 19288 26364
rect 20916 26336 21772 26364
rect 18555 26333 18567 26336
rect 18509 26327 18567 26333
rect 19260 26308 19288 26336
rect 19242 26256 19248 26308
rect 19300 26256 19306 26308
rect 19978 26256 19984 26308
rect 20036 26256 20042 26308
rect 21542 26296 21548 26308
rect 21503 26268 21548 26296
rect 21542 26256 21548 26268
rect 21600 26256 21606 26308
rect 21744 26296 21772 26336
rect 21821 26333 21833 26367
rect 21867 26364 21879 26367
rect 22186 26364 22192 26376
rect 21867 26336 22192 26364
rect 21867 26333 21879 26336
rect 21821 26327 21879 26333
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 23474 26364 23480 26376
rect 23435 26336 23480 26364
rect 23474 26324 23480 26336
rect 23532 26324 23538 26376
rect 23584 26373 23612 26472
rect 23658 26460 23664 26512
rect 23716 26460 23722 26512
rect 23750 26460 23756 26512
rect 23808 26500 23814 26512
rect 23808 26472 24440 26500
rect 23808 26460 23814 26472
rect 23676 26373 23704 26460
rect 24412 26444 24440 26472
rect 24394 26432 24400 26444
rect 24307 26404 24400 26432
rect 24394 26392 24400 26404
rect 24452 26392 24458 26444
rect 23569 26367 23627 26373
rect 23569 26333 23581 26367
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 23661 26367 23719 26373
rect 23661 26333 23673 26367
rect 23707 26333 23719 26367
rect 23661 26327 23719 26333
rect 23750 26324 23756 26376
rect 23808 26364 23814 26376
rect 23845 26367 23903 26373
rect 23845 26364 23857 26367
rect 23808 26336 23857 26364
rect 23808 26324 23814 26336
rect 23845 26333 23857 26336
rect 23891 26333 23903 26367
rect 23845 26327 23903 26333
rect 23201 26299 23259 26305
rect 21744 26268 22094 26296
rect 22066 26240 22094 26268
rect 23201 26265 23213 26299
rect 23247 26296 23259 26299
rect 24504 26296 24532 26540
rect 28626 26528 28632 26580
rect 28684 26568 28690 26580
rect 33134 26568 33140 26580
rect 28684 26540 30144 26568
rect 33095 26540 33140 26568
rect 28684 26528 28690 26540
rect 26602 26500 26608 26512
rect 24688 26472 26372 26500
rect 26515 26472 26608 26500
rect 24688 26444 24716 26472
rect 24670 26432 24676 26444
rect 24631 26404 24676 26432
rect 24670 26392 24676 26404
rect 24728 26392 24734 26444
rect 24762 26392 24768 26444
rect 24820 26432 24826 26444
rect 24882 26435 24940 26441
rect 24882 26432 24894 26435
rect 24820 26404 24894 26432
rect 24820 26392 24826 26404
rect 24882 26401 24894 26404
rect 24928 26401 24940 26435
rect 24882 26395 24940 26401
rect 26145 26367 26203 26373
rect 26145 26333 26157 26367
rect 26191 26364 26203 26367
rect 26234 26364 26240 26376
rect 26191 26336 26240 26364
rect 26191 26333 26203 26336
rect 26145 26327 26203 26333
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 26344 26373 26372 26472
rect 26602 26460 26608 26472
rect 26660 26500 26666 26512
rect 30116 26509 30144 26540
rect 33134 26528 33140 26540
rect 33192 26528 33198 26580
rect 33870 26568 33876 26580
rect 33831 26540 33876 26568
rect 33870 26528 33876 26540
rect 33928 26528 33934 26580
rect 30101 26503 30159 26509
rect 26660 26472 29776 26500
rect 26660 26460 26666 26472
rect 26697 26435 26755 26441
rect 26697 26401 26709 26435
rect 26743 26432 26755 26435
rect 27525 26435 27583 26441
rect 27525 26432 27537 26435
rect 26743 26404 27537 26432
rect 26743 26401 26755 26404
rect 26697 26395 26755 26401
rect 27525 26401 27537 26404
rect 27571 26432 27583 26435
rect 27571 26404 29132 26432
rect 27571 26401 27583 26404
rect 27525 26395 27583 26401
rect 26329 26367 26387 26373
rect 26329 26333 26341 26367
rect 26375 26333 26387 26367
rect 26329 26327 26387 26333
rect 28169 26367 28227 26373
rect 28169 26333 28181 26367
rect 28215 26364 28227 26367
rect 28997 26367 29055 26373
rect 28997 26364 29009 26367
rect 28215 26336 29009 26364
rect 28215 26333 28227 26336
rect 28169 26327 28227 26333
rect 28997 26333 29009 26336
rect 29043 26333 29055 26367
rect 29104 26364 29132 26404
rect 29178 26364 29184 26376
rect 29104 26336 29184 26364
rect 28997 26327 29055 26333
rect 29178 26324 29184 26336
rect 29236 26364 29242 26376
rect 29236 26336 29329 26364
rect 29236 26324 29242 26336
rect 24765 26299 24823 26305
rect 24765 26296 24777 26299
rect 23247 26268 23888 26296
rect 24504 26268 24777 26296
rect 23247 26265 23259 26268
rect 23201 26259 23259 26265
rect 23860 26240 23888 26268
rect 24765 26265 24777 26268
rect 24811 26265 24823 26299
rect 24765 26259 24823 26265
rect 25958 26256 25964 26308
rect 26016 26296 26022 26308
rect 27341 26299 27399 26305
rect 27341 26296 27353 26299
rect 26016 26268 27353 26296
rect 26016 26256 26022 26268
rect 27341 26265 27353 26268
rect 27387 26296 27399 26299
rect 27430 26296 27436 26308
rect 27387 26268 27436 26296
rect 27387 26265 27399 26268
rect 27341 26259 27399 26265
rect 27430 26256 27436 26268
rect 27488 26256 27494 26308
rect 28626 26296 28632 26308
rect 28587 26268 28632 26296
rect 28626 26256 28632 26268
rect 28684 26256 28690 26308
rect 28810 26296 28816 26308
rect 28771 26268 28816 26296
rect 28810 26256 28816 26268
rect 28868 26256 28874 26308
rect 22066 26200 22100 26240
rect 22094 26188 22100 26200
rect 22152 26188 22158 26240
rect 23842 26188 23848 26240
rect 23900 26188 23906 26240
rect 25041 26231 25099 26237
rect 25041 26197 25053 26231
rect 25087 26228 25099 26231
rect 25130 26228 25136 26240
rect 25087 26200 25136 26228
rect 25087 26197 25099 26200
rect 25041 26191 25099 26197
rect 25130 26188 25136 26200
rect 25188 26188 25194 26240
rect 27982 26228 27988 26240
rect 27943 26200 27988 26228
rect 27982 26188 27988 26200
rect 28040 26188 28046 26240
rect 29288 26228 29316 26336
rect 29454 26324 29460 26376
rect 29512 26364 29518 26376
rect 29748 26373 29776 26472
rect 30101 26469 30113 26503
rect 30147 26469 30159 26503
rect 30101 26463 30159 26469
rect 32861 26435 32919 26441
rect 32861 26401 32873 26435
rect 32907 26432 32919 26435
rect 34606 26432 34612 26444
rect 32907 26404 34612 26432
rect 32907 26401 32919 26404
rect 32861 26395 32919 26401
rect 34606 26392 34612 26404
rect 34664 26392 34670 26444
rect 34977 26435 35035 26441
rect 34977 26401 34989 26435
rect 35023 26432 35035 26435
rect 35342 26432 35348 26444
rect 35023 26404 35348 26432
rect 35023 26401 35035 26404
rect 34977 26395 35035 26401
rect 35342 26392 35348 26404
rect 35400 26392 35406 26444
rect 35986 26392 35992 26444
rect 36044 26432 36050 26444
rect 36449 26435 36507 26441
rect 36449 26432 36461 26435
rect 36044 26404 36461 26432
rect 36044 26392 36050 26404
rect 36449 26401 36461 26404
rect 36495 26401 36507 26435
rect 36449 26395 36507 26401
rect 39301 26435 39359 26441
rect 39301 26401 39313 26435
rect 39347 26432 39359 26435
rect 42794 26432 42800 26444
rect 39347 26404 42800 26432
rect 39347 26401 39359 26404
rect 39301 26395 39359 26401
rect 42794 26392 42800 26404
rect 42852 26392 42858 26444
rect 29549 26367 29607 26373
rect 29549 26364 29561 26367
rect 29512 26336 29561 26364
rect 29512 26324 29518 26336
rect 29549 26333 29561 26336
rect 29595 26333 29607 26367
rect 29549 26327 29607 26333
rect 29733 26367 29791 26373
rect 29733 26333 29745 26367
rect 29779 26333 29791 26367
rect 29914 26364 29920 26376
rect 29875 26336 29920 26364
rect 29733 26327 29791 26333
rect 29914 26324 29920 26336
rect 29972 26324 29978 26376
rect 32674 26324 32680 26376
rect 32732 26364 32738 26376
rect 32769 26367 32827 26373
rect 32769 26364 32781 26367
rect 32732 26336 32781 26364
rect 32732 26324 32738 26336
rect 32769 26333 32781 26336
rect 32815 26333 32827 26367
rect 32769 26327 32827 26333
rect 33873 26367 33931 26373
rect 33873 26333 33885 26367
rect 33919 26364 33931 26367
rect 33962 26364 33968 26376
rect 33919 26336 33968 26364
rect 33919 26333 33931 26336
rect 33873 26327 33931 26333
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34149 26367 34207 26373
rect 34149 26333 34161 26367
rect 34195 26333 34207 26367
rect 34149 26327 34207 26333
rect 29825 26299 29883 26305
rect 29825 26296 29837 26299
rect 29472 26268 29837 26296
rect 29472 26228 29500 26268
rect 29825 26265 29837 26268
rect 29871 26265 29883 26299
rect 29825 26259 29883 26265
rect 34057 26299 34115 26305
rect 34057 26265 34069 26299
rect 34103 26265 34115 26299
rect 34164 26296 34192 26327
rect 34422 26324 34428 26376
rect 34480 26364 34486 26376
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 34480 26336 34713 26364
rect 34480 26324 34486 26336
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34701 26327 34759 26333
rect 36906 26324 36912 26376
rect 36964 26364 36970 26376
rect 37461 26367 37519 26373
rect 37461 26364 37473 26367
rect 36964 26336 37473 26364
rect 36964 26324 36970 26336
rect 37461 26333 37473 26336
rect 37507 26333 37519 26367
rect 37461 26327 37519 26333
rect 34606 26296 34612 26308
rect 34164 26268 34612 26296
rect 34057 26259 34115 26265
rect 29288 26200 29500 26228
rect 34072 26228 34100 26259
rect 34606 26256 34612 26268
rect 34664 26256 34670 26308
rect 35986 26256 35992 26308
rect 36044 26256 36050 26308
rect 37642 26296 37648 26308
rect 37603 26268 37648 26296
rect 37642 26256 37648 26268
rect 37700 26256 37706 26308
rect 34882 26228 34888 26240
rect 34072 26200 34888 26228
rect 34882 26188 34888 26200
rect 34940 26188 34946 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 19337 26027 19395 26033
rect 19337 25993 19349 26027
rect 19383 26024 19395 26027
rect 19978 26024 19984 26036
rect 19383 25996 19984 26024
rect 19383 25993 19395 25996
rect 19337 25987 19395 25993
rect 19978 25984 19984 25996
rect 20036 25984 20042 26036
rect 20162 25984 20168 26036
rect 20220 26024 20226 26036
rect 20257 26027 20315 26033
rect 20257 26024 20269 26027
rect 20220 25996 20269 26024
rect 20220 25984 20226 25996
rect 20257 25993 20269 25996
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 24305 26027 24363 26033
rect 24305 25993 24317 26027
rect 24351 26024 24363 26027
rect 24394 26024 24400 26036
rect 24351 25996 24400 26024
rect 24351 25993 24363 25996
rect 24305 25987 24363 25993
rect 24394 25984 24400 25996
rect 24452 25984 24458 26036
rect 29454 25984 29460 26036
rect 29512 26024 29518 26036
rect 30101 26027 30159 26033
rect 30101 26024 30113 26027
rect 29512 25996 30113 26024
rect 29512 25984 29518 25996
rect 30101 25993 30113 25996
rect 30147 25993 30159 26027
rect 30101 25987 30159 25993
rect 33781 26027 33839 26033
rect 33781 25993 33793 26027
rect 33827 26024 33839 26027
rect 34422 26024 34428 26036
rect 33827 25996 34428 26024
rect 33827 25993 33839 25996
rect 33781 25987 33839 25993
rect 34422 25984 34428 25996
rect 34480 25984 34486 26036
rect 34790 25984 34796 26036
rect 34848 26024 34854 26036
rect 34885 26027 34943 26033
rect 34885 26024 34897 26027
rect 34848 25996 34897 26024
rect 34848 25984 34854 25996
rect 34885 25993 34897 25996
rect 34931 25993 34943 26027
rect 34885 25987 34943 25993
rect 35713 26027 35771 26033
rect 35713 25993 35725 26027
rect 35759 26024 35771 26027
rect 35986 26024 35992 26036
rect 35759 25996 35992 26024
rect 35759 25993 35771 25996
rect 35713 25987 35771 25993
rect 35986 25984 35992 25996
rect 36044 25984 36050 26036
rect 23566 25916 23572 25968
rect 23624 25916 23630 25968
rect 24854 25916 24860 25968
rect 24912 25956 24918 25968
rect 24949 25959 25007 25965
rect 24949 25956 24961 25959
rect 24912 25928 24961 25956
rect 24912 25916 24918 25928
rect 24949 25925 24961 25928
rect 24995 25925 25007 25959
rect 24949 25919 25007 25925
rect 25041 25959 25099 25965
rect 25041 25925 25053 25959
rect 25087 25956 25099 25959
rect 26510 25956 26516 25968
rect 25087 25928 26516 25956
rect 25087 25925 25099 25928
rect 25041 25919 25099 25925
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25888 12311 25891
rect 19242 25888 19248 25900
rect 12299 25860 14320 25888
rect 19203 25860 19248 25888
rect 12299 25857 12311 25860
rect 12253 25851 12311 25857
rect 14292 25832 14320 25860
rect 19242 25848 19248 25860
rect 19300 25848 19306 25900
rect 19334 25848 19340 25900
rect 19392 25888 19398 25900
rect 19889 25891 19947 25897
rect 19889 25888 19901 25891
rect 19392 25860 19901 25888
rect 19392 25848 19398 25860
rect 19889 25857 19901 25860
rect 19935 25857 19947 25891
rect 19889 25851 19947 25857
rect 20073 25891 20131 25897
rect 20073 25857 20085 25891
rect 20119 25888 20131 25891
rect 21174 25888 21180 25900
rect 20119 25860 21180 25888
rect 20119 25857 20131 25860
rect 20073 25851 20131 25857
rect 21174 25848 21180 25860
rect 21232 25848 21238 25900
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22557 25891 22615 25897
rect 22557 25888 22569 25891
rect 22152 25860 22569 25888
rect 22152 25848 22158 25860
rect 22557 25857 22569 25860
rect 22603 25857 22615 25891
rect 24762 25888 24768 25900
rect 24723 25860 24768 25888
rect 22557 25851 22615 25857
rect 24762 25848 24768 25860
rect 24820 25848 24826 25900
rect 12342 25820 12348 25832
rect 12303 25792 12348 25820
rect 12342 25780 12348 25792
rect 12400 25780 12406 25832
rect 14274 25780 14280 25832
rect 14332 25820 14338 25832
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 14332 25792 16681 25820
rect 14332 25780 14338 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 16850 25820 16856 25832
rect 16811 25792 16856 25820
rect 16669 25783 16727 25789
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 17129 25823 17187 25829
rect 17129 25789 17141 25823
rect 17175 25789 17187 25823
rect 17129 25783 17187 25789
rect 22833 25823 22891 25829
rect 22833 25789 22845 25823
rect 22879 25820 22891 25823
rect 23290 25820 23296 25832
rect 22879 25792 23296 25820
rect 22879 25789 22891 25792
rect 22833 25783 22891 25789
rect 12621 25755 12679 25761
rect 12621 25721 12633 25755
rect 12667 25752 12679 25755
rect 12802 25752 12808 25764
rect 12667 25724 12808 25752
rect 12667 25721 12679 25724
rect 12621 25715 12679 25721
rect 12802 25712 12808 25724
rect 12860 25712 12866 25764
rect 16758 25712 16764 25764
rect 16816 25752 16822 25764
rect 17144 25752 17172 25783
rect 23290 25780 23296 25792
rect 23348 25780 23354 25832
rect 24118 25780 24124 25832
rect 24176 25820 24182 25832
rect 25056 25820 25084 25919
rect 26510 25916 26516 25928
rect 26568 25916 26574 25968
rect 27982 25916 27988 25968
rect 28040 25956 28046 25968
rect 28629 25959 28687 25965
rect 28629 25956 28641 25959
rect 28040 25928 28641 25956
rect 28040 25916 28046 25928
rect 28629 25925 28641 25928
rect 28675 25925 28687 25959
rect 28629 25919 28687 25925
rect 29638 25916 29644 25968
rect 29696 25916 29702 25968
rect 34330 25956 34336 25968
rect 34291 25928 34336 25956
rect 34330 25916 34336 25928
rect 34388 25916 34394 25968
rect 34517 25959 34575 25965
rect 34517 25925 34529 25959
rect 34563 25956 34575 25959
rect 35802 25956 35808 25968
rect 34563 25928 35808 25956
rect 34563 25925 34575 25928
rect 34517 25919 34575 25925
rect 35802 25916 35808 25928
rect 35860 25916 35866 25968
rect 25133 25891 25191 25897
rect 25133 25857 25145 25891
rect 25179 25888 25191 25891
rect 25314 25888 25320 25900
rect 25179 25860 25320 25888
rect 25179 25857 25191 25860
rect 25133 25851 25191 25857
rect 25314 25848 25320 25860
rect 25372 25848 25378 25900
rect 27246 25848 27252 25900
rect 27304 25888 27310 25900
rect 28353 25891 28411 25897
rect 28353 25888 28365 25891
rect 27304 25860 28365 25888
rect 27304 25848 27310 25860
rect 28353 25857 28365 25860
rect 28399 25857 28411 25891
rect 28353 25851 28411 25857
rect 33597 25891 33655 25897
rect 33597 25857 33609 25891
rect 33643 25857 33655 25891
rect 33597 25851 33655 25857
rect 34609 25891 34667 25897
rect 34609 25857 34621 25891
rect 34655 25857 34667 25891
rect 34609 25851 34667 25857
rect 24176 25792 25084 25820
rect 24176 25780 24182 25792
rect 27338 25780 27344 25832
rect 27396 25820 27402 25832
rect 32490 25820 32496 25832
rect 27396 25792 32496 25820
rect 27396 25780 27402 25792
rect 32490 25780 32496 25792
rect 32548 25820 32554 25832
rect 33612 25820 33640 25851
rect 32548 25792 33640 25820
rect 34624 25820 34652 25851
rect 34698 25848 34704 25900
rect 34756 25888 34762 25900
rect 34756 25860 34801 25888
rect 34756 25848 34762 25860
rect 35526 25848 35532 25900
rect 35584 25888 35590 25900
rect 35621 25891 35679 25897
rect 35621 25888 35633 25891
rect 35584 25860 35633 25888
rect 35584 25848 35590 25860
rect 35621 25857 35633 25860
rect 35667 25857 35679 25891
rect 44910 25888 44916 25900
rect 44871 25860 44916 25888
rect 35621 25851 35679 25857
rect 34790 25820 34796 25832
rect 34624 25792 34796 25820
rect 32548 25780 32554 25792
rect 34790 25780 34796 25792
rect 34848 25780 34854 25832
rect 16816 25724 17172 25752
rect 16816 25712 16822 25724
rect 34514 25712 34520 25764
rect 34572 25752 34578 25764
rect 35636 25752 35664 25851
rect 44910 25848 44916 25860
rect 44968 25848 44974 25900
rect 34572 25724 35664 25752
rect 34572 25712 34578 25724
rect 20070 25684 20076 25696
rect 20031 25656 20076 25684
rect 20070 25644 20076 25656
rect 20128 25644 20134 25696
rect 25038 25644 25044 25696
rect 25096 25684 25102 25696
rect 25317 25687 25375 25693
rect 25317 25684 25329 25687
rect 25096 25656 25329 25684
rect 25096 25644 25102 25656
rect 25317 25653 25329 25656
rect 25363 25653 25375 25687
rect 25317 25647 25375 25653
rect 45005 25687 45063 25693
rect 45005 25653 45017 25687
rect 45051 25684 45063 25687
rect 45462 25684 45468 25696
rect 45051 25656 45468 25684
rect 45051 25653 45063 25656
rect 45005 25647 45063 25653
rect 45462 25644 45468 25656
rect 45520 25644 45526 25696
rect 46198 25644 46204 25696
rect 46256 25684 46262 25696
rect 47765 25687 47823 25693
rect 47765 25684 47777 25687
rect 46256 25656 47777 25684
rect 46256 25644 46262 25656
rect 47765 25653 47777 25656
rect 47811 25653 47823 25687
rect 47765 25647 47823 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 12342 25440 12348 25492
rect 12400 25480 12406 25492
rect 12713 25483 12771 25489
rect 12713 25480 12725 25483
rect 12400 25452 12725 25480
rect 12400 25440 12406 25452
rect 12713 25449 12725 25452
rect 12759 25449 12771 25483
rect 19426 25480 19432 25492
rect 19387 25452 19432 25480
rect 12713 25443 12771 25449
rect 19426 25440 19432 25452
rect 19484 25440 19490 25492
rect 21453 25483 21511 25489
rect 21453 25449 21465 25483
rect 21499 25480 21511 25483
rect 21542 25480 21548 25492
rect 21499 25452 21548 25480
rect 21499 25449 21511 25452
rect 21453 25443 21511 25449
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 21637 25483 21695 25489
rect 21637 25449 21649 25483
rect 21683 25480 21695 25483
rect 21910 25480 21916 25492
rect 21683 25452 21916 25480
rect 21683 25449 21695 25452
rect 21637 25443 21695 25449
rect 21910 25440 21916 25452
rect 21968 25440 21974 25492
rect 23290 25480 23296 25492
rect 23251 25452 23296 25480
rect 23290 25440 23296 25452
rect 23348 25440 23354 25492
rect 25130 25480 25136 25492
rect 23860 25452 25136 25480
rect 19242 25372 19248 25424
rect 19300 25412 19306 25424
rect 20165 25415 20223 25421
rect 20165 25412 20177 25415
rect 19300 25384 20177 25412
rect 19300 25372 19306 25384
rect 20165 25381 20177 25384
rect 20211 25412 20223 25415
rect 23658 25412 23664 25424
rect 20211 25384 23664 25412
rect 20211 25381 20223 25384
rect 20165 25375 20223 25381
rect 23658 25372 23664 25384
rect 23716 25372 23722 25424
rect 8294 25304 8300 25356
rect 8352 25344 8358 25356
rect 16669 25347 16727 25353
rect 16669 25344 16681 25347
rect 8352 25316 16681 25344
rect 8352 25304 8358 25316
rect 16669 25313 16681 25316
rect 16715 25313 16727 25347
rect 16669 25307 16727 25313
rect 21545 25347 21603 25353
rect 21545 25313 21557 25347
rect 21591 25344 21603 25347
rect 21634 25344 21640 25356
rect 21591 25316 21640 25344
rect 21591 25313 21603 25316
rect 21545 25307 21603 25313
rect 21634 25304 21640 25316
rect 21692 25304 21698 25356
rect 23860 25344 23888 25452
rect 25130 25440 25136 25452
rect 25188 25440 25194 25492
rect 25222 25440 25228 25492
rect 25280 25480 25286 25492
rect 26513 25483 26571 25489
rect 26513 25480 26525 25483
rect 25280 25452 26525 25480
rect 25280 25440 25286 25452
rect 26513 25449 26525 25452
rect 26559 25449 26571 25483
rect 29638 25480 29644 25492
rect 29599 25452 29644 25480
rect 26513 25443 26571 25449
rect 29638 25440 29644 25452
rect 29696 25440 29702 25492
rect 32769 25483 32827 25489
rect 32769 25449 32781 25483
rect 32815 25480 32827 25483
rect 34514 25480 34520 25492
rect 32815 25452 34520 25480
rect 32815 25449 32827 25452
rect 32769 25443 32827 25449
rect 34514 25440 34520 25452
rect 34572 25440 34578 25492
rect 37642 25440 37648 25492
rect 37700 25480 37706 25492
rect 37921 25483 37979 25489
rect 37921 25480 37933 25483
rect 37700 25452 37933 25480
rect 37700 25440 37706 25452
rect 37921 25449 37933 25452
rect 37967 25449 37979 25483
rect 37921 25443 37979 25449
rect 37182 25372 37188 25424
rect 37240 25412 37246 25424
rect 45830 25412 45836 25424
rect 37240 25384 45836 25412
rect 37240 25372 37246 25384
rect 45830 25372 45836 25384
rect 45888 25372 45894 25424
rect 23768 25316 23888 25344
rect 24765 25347 24823 25353
rect 11977 25279 12035 25285
rect 11977 25245 11989 25279
rect 12023 25276 12035 25279
rect 12250 25276 12256 25288
rect 12023 25248 12256 25276
rect 12023 25245 12035 25248
rect 11977 25239 12035 25245
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25245 12679 25279
rect 12621 25239 12679 25245
rect 12805 25279 12863 25285
rect 12805 25245 12817 25279
rect 12851 25276 12863 25279
rect 13722 25276 13728 25288
rect 12851 25248 13728 25276
rect 12851 25245 12863 25248
rect 12805 25239 12863 25245
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 12636 25208 12664 25239
rect 13722 25236 13728 25248
rect 13780 25236 13786 25288
rect 13906 25236 13912 25288
rect 13964 25276 13970 25288
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 13964 25248 14105 25276
rect 13964 25236 13970 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 15286 25236 15292 25288
rect 15344 25276 15350 25288
rect 16022 25276 16028 25288
rect 15344 25248 16028 25276
rect 15344 25236 15350 25248
rect 16022 25236 16028 25248
rect 16080 25276 16086 25288
rect 16209 25279 16267 25285
rect 16209 25276 16221 25279
rect 16080 25248 16221 25276
rect 16080 25236 16086 25248
rect 16209 25245 16221 25248
rect 16255 25245 16267 25279
rect 16209 25239 16267 25245
rect 18138 25236 18144 25288
rect 18196 25276 18202 25288
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 18196 25248 19257 25276
rect 18196 25236 18202 25248
rect 19245 25245 19257 25248
rect 19291 25276 19303 25279
rect 19981 25279 20039 25285
rect 19981 25276 19993 25279
rect 19291 25248 19993 25276
rect 19291 25245 19303 25248
rect 19245 25239 19303 25245
rect 19981 25245 19993 25248
rect 20027 25276 20039 25279
rect 20530 25276 20536 25288
rect 20027 25248 20536 25276
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 21358 25276 21364 25288
rect 21319 25248 21364 25276
rect 21358 25236 21364 25248
rect 21416 25236 21422 25288
rect 21726 25276 21732 25288
rect 21687 25248 21732 25276
rect 21726 25236 21732 25248
rect 21784 25236 21790 25288
rect 23474 25276 23480 25288
rect 23435 25248 23480 25276
rect 23474 25236 23480 25248
rect 23532 25236 23538 25288
rect 23768 25285 23796 25316
rect 24765 25313 24777 25347
rect 24811 25344 24823 25347
rect 27246 25344 27252 25356
rect 24811 25316 27252 25344
rect 24811 25313 24823 25316
rect 24765 25307 24823 25313
rect 27246 25304 27252 25316
rect 27304 25304 27310 25356
rect 36078 25304 36084 25356
rect 36136 25344 36142 25356
rect 39945 25347 40003 25353
rect 39945 25344 39957 25347
rect 36136 25316 39957 25344
rect 36136 25304 36142 25316
rect 39945 25313 39957 25316
rect 39991 25313 40003 25347
rect 41782 25344 41788 25356
rect 41743 25316 41788 25344
rect 39945 25307 40003 25313
rect 41782 25304 41788 25316
rect 41840 25304 41846 25356
rect 45462 25344 45468 25356
rect 45423 25316 45468 25344
rect 45462 25304 45468 25316
rect 45520 25304 45526 25356
rect 46842 25344 46848 25356
rect 46803 25316 46848 25344
rect 46842 25304 46848 25316
rect 46900 25304 46906 25356
rect 23569 25279 23627 25285
rect 23569 25245 23581 25279
rect 23615 25245 23627 25279
rect 23569 25239 23627 25245
rect 23753 25279 23811 25285
rect 23753 25245 23765 25279
rect 23799 25245 23811 25279
rect 23753 25239 23811 25245
rect 13354 25208 13360 25220
rect 12636 25180 13360 25208
rect 13354 25168 13360 25180
rect 13412 25168 13418 25220
rect 16393 25211 16451 25217
rect 16393 25177 16405 25211
rect 16439 25208 16451 25211
rect 17402 25208 17408 25220
rect 16439 25180 17408 25208
rect 16439 25177 16451 25180
rect 16393 25171 16451 25177
rect 17402 25168 17408 25180
rect 17460 25168 17466 25220
rect 23584 25208 23612 25239
rect 23842 25236 23848 25288
rect 23900 25276 23906 25288
rect 23900 25248 23945 25276
rect 23900 25236 23906 25248
rect 27890 25236 27896 25288
rect 27948 25276 27954 25288
rect 28902 25276 28908 25288
rect 27948 25248 28908 25276
rect 27948 25236 27954 25248
rect 28902 25236 28908 25248
rect 28960 25276 28966 25288
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 28960 25248 29561 25276
rect 28960 25236 28966 25248
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 29730 25236 29736 25288
rect 29788 25276 29794 25288
rect 32585 25279 32643 25285
rect 32585 25276 32597 25279
rect 29788 25248 32597 25276
rect 29788 25236 29794 25248
rect 32585 25245 32597 25248
rect 32631 25245 32643 25279
rect 32585 25239 32643 25245
rect 35894 25236 35900 25288
rect 35952 25276 35958 25288
rect 36170 25276 36176 25288
rect 35952 25248 36176 25276
rect 35952 25236 35958 25248
rect 36170 25236 36176 25248
rect 36228 25276 36234 25288
rect 37182 25276 37188 25288
rect 36228 25248 37188 25276
rect 36228 25236 36234 25248
rect 37182 25236 37188 25248
rect 37240 25236 37246 25288
rect 37826 25276 37832 25288
rect 37787 25248 37832 25276
rect 37826 25236 37832 25248
rect 37884 25236 37890 25288
rect 45002 25236 45008 25288
rect 45060 25276 45066 25288
rect 45281 25279 45339 25285
rect 45281 25276 45293 25279
rect 45060 25248 45293 25276
rect 45060 25236 45066 25248
rect 45281 25245 45293 25248
rect 45327 25245 45339 25279
rect 47762 25276 47768 25288
rect 47723 25248 47768 25276
rect 45281 25239 45339 25245
rect 47762 25236 47768 25248
rect 47820 25236 47826 25288
rect 24118 25208 24124 25220
rect 23584 25180 24124 25208
rect 24118 25168 24124 25180
rect 24176 25168 24182 25220
rect 25038 25208 25044 25220
rect 24999 25180 25044 25208
rect 25038 25168 25044 25180
rect 25096 25168 25102 25220
rect 25590 25168 25596 25220
rect 25648 25168 25654 25220
rect 40126 25208 40132 25220
rect 40087 25180 40132 25208
rect 40126 25168 40132 25180
rect 40184 25168 40190 25220
rect 2130 25140 2136 25152
rect 2091 25112 2136 25140
rect 2130 25100 2136 25112
rect 2188 25100 2194 25152
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 12526 25140 12532 25152
rect 12115 25112 12532 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 12526 25100 12532 25112
rect 12584 25100 12590 25152
rect 14182 25140 14188 25152
rect 14143 25112 14188 25140
rect 14182 25100 14188 25112
rect 14240 25100 14246 25152
rect 21085 25143 21143 25149
rect 21085 25109 21097 25143
rect 21131 25140 21143 25143
rect 22370 25140 22376 25152
rect 21131 25112 22376 25140
rect 21131 25109 21143 25112
rect 21085 25103 21143 25109
rect 22370 25100 22376 25112
rect 22428 25140 22434 25152
rect 27522 25140 27528 25152
rect 22428 25112 27528 25140
rect 22428 25100 22434 25112
rect 27522 25100 27528 25112
rect 27580 25100 27586 25152
rect 37277 25143 37335 25149
rect 37277 25109 37289 25143
rect 37323 25140 37335 25143
rect 37458 25140 37464 25152
rect 37323 25112 37464 25140
rect 37323 25109 37335 25112
rect 37277 25103 37335 25109
rect 37458 25100 37464 25112
rect 37516 25100 37522 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 2130 24896 2136 24948
rect 2188 24936 2194 24948
rect 2188 24908 22094 24936
rect 2188 24896 2194 24908
rect 12802 24868 12808 24880
rect 12763 24840 12808 24868
rect 12802 24828 12808 24840
rect 12860 24828 12866 24880
rect 14182 24868 14188 24880
rect 14030 24840 14188 24868
rect 14182 24828 14188 24840
rect 14240 24828 14246 24880
rect 22066 24868 22094 24908
rect 25866 24896 25872 24948
rect 25924 24936 25930 24948
rect 27798 24936 27804 24948
rect 25924 24908 27804 24936
rect 25924 24896 25930 24908
rect 27798 24896 27804 24908
rect 27856 24896 27862 24948
rect 27890 24896 27896 24948
rect 27948 24936 27954 24948
rect 28445 24939 28503 24945
rect 28445 24936 28457 24939
rect 27948 24908 28457 24936
rect 27948 24896 27954 24908
rect 28445 24905 28457 24908
rect 28491 24905 28503 24939
rect 40126 24936 40132 24948
rect 40087 24908 40132 24936
rect 28445 24899 28503 24905
rect 40126 24896 40132 24908
rect 40184 24896 40190 24948
rect 44818 24868 44824 24880
rect 14936 24840 15976 24868
rect 22066 24840 38700 24868
rect 11977 24803 12035 24809
rect 11977 24769 11989 24803
rect 12023 24800 12035 24803
rect 12250 24800 12256 24812
rect 12023 24772 12256 24800
rect 12023 24769 12035 24772
rect 11977 24763 12035 24769
rect 12250 24760 12256 24772
rect 12308 24760 12314 24812
rect 12526 24800 12532 24812
rect 12487 24772 12532 24800
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 14090 24760 14096 24812
rect 14148 24800 14154 24812
rect 14936 24800 14964 24840
rect 14148 24772 14964 24800
rect 15013 24803 15071 24809
rect 14148 24760 14154 24772
rect 15013 24769 15025 24803
rect 15059 24800 15071 24803
rect 15654 24800 15660 24812
rect 15059 24772 15660 24800
rect 15059 24769 15071 24772
rect 15013 24763 15071 24769
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 15746 24760 15752 24812
rect 15804 24800 15810 24812
rect 15948 24800 15976 24840
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 15804 24772 15849 24800
rect 15948 24772 16681 24800
rect 15804 24760 15810 24772
rect 16669 24769 16681 24772
rect 16715 24800 16727 24803
rect 17126 24800 17132 24812
rect 16715 24772 17132 24800
rect 16715 24769 16727 24772
rect 16669 24763 16727 24769
rect 17126 24760 17132 24772
rect 17184 24760 17190 24812
rect 17310 24800 17316 24812
rect 17271 24772 17316 24800
rect 17310 24760 17316 24772
rect 17368 24760 17374 24812
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 18138 24800 18144 24812
rect 17460 24772 17505 24800
rect 18099 24772 18144 24800
rect 17460 24760 17466 24772
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 19334 24800 19340 24812
rect 19295 24772 19340 24800
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 23477 24803 23535 24809
rect 23477 24769 23489 24803
rect 23523 24769 23535 24803
rect 23477 24763 23535 24769
rect 14274 24732 14280 24744
rect 14235 24704 14280 24732
rect 14274 24692 14280 24704
rect 14332 24692 14338 24744
rect 14826 24732 14832 24744
rect 14787 24704 14832 24732
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 15197 24735 15255 24741
rect 15197 24732 15209 24735
rect 15120 24704 15209 24732
rect 15120 24664 15148 24704
rect 15197 24701 15209 24704
rect 15243 24701 15255 24735
rect 15197 24695 15255 24701
rect 15286 24692 15292 24744
rect 15344 24732 15350 24744
rect 15344 24704 15389 24732
rect 15344 24692 15350 24704
rect 15930 24692 15936 24744
rect 15988 24732 15994 24744
rect 19521 24735 19579 24741
rect 19521 24732 19533 24735
rect 15988 24704 19533 24732
rect 15988 24692 15994 24704
rect 19521 24701 19533 24704
rect 19567 24732 19579 24735
rect 20990 24732 20996 24744
rect 19567 24704 20996 24732
rect 19567 24701 19579 24704
rect 19521 24695 19579 24701
rect 20990 24692 20996 24704
rect 21048 24692 21054 24744
rect 23492 24732 23520 24763
rect 23566 24760 23572 24812
rect 23624 24800 23630 24812
rect 25501 24803 25559 24809
rect 23624 24772 23669 24800
rect 23624 24760 23630 24772
rect 25501 24769 25513 24803
rect 25547 24769 25559 24803
rect 25501 24763 25559 24769
rect 23658 24732 23664 24744
rect 23492 24704 23664 24732
rect 23658 24692 23664 24704
rect 23716 24732 23722 24744
rect 24762 24732 24768 24744
rect 23716 24704 24768 24732
rect 23716 24692 23722 24704
rect 24762 24692 24768 24704
rect 24820 24732 24826 24744
rect 25516 24732 25544 24763
rect 25590 24760 25596 24812
rect 25648 24800 25654 24812
rect 25648 24772 25693 24800
rect 25648 24760 25654 24772
rect 26786 24760 26792 24812
rect 26844 24800 26850 24812
rect 27433 24803 27491 24809
rect 26844 24798 27384 24800
rect 27433 24798 27445 24803
rect 26844 24772 27445 24798
rect 26844 24760 26850 24772
rect 27356 24770 27445 24772
rect 27433 24769 27445 24770
rect 27479 24769 27491 24803
rect 27433 24763 27491 24769
rect 27540 24772 27752 24800
rect 27540 24744 27568 24772
rect 27522 24732 27528 24744
rect 24820 24704 25544 24732
rect 27483 24704 27528 24732
rect 24820 24692 24826 24704
rect 27522 24692 27528 24704
rect 27580 24692 27586 24744
rect 27724 24732 27752 24772
rect 27798 24760 27804 24812
rect 27856 24800 27862 24812
rect 28261 24803 28319 24809
rect 28261 24800 28273 24803
rect 27856 24772 28273 24800
rect 27856 24760 27862 24772
rect 28261 24769 28273 24772
rect 28307 24769 28319 24803
rect 28261 24763 28319 24769
rect 31205 24803 31263 24809
rect 31205 24769 31217 24803
rect 31251 24800 31263 24803
rect 31294 24800 31300 24812
rect 31251 24772 31300 24800
rect 31251 24769 31263 24772
rect 31205 24763 31263 24769
rect 31294 24760 31300 24772
rect 31352 24760 31358 24812
rect 31389 24803 31447 24809
rect 31389 24769 31401 24803
rect 31435 24800 31447 24803
rect 31478 24800 31484 24812
rect 31435 24772 31484 24800
rect 31435 24769 31447 24772
rect 31389 24763 31447 24769
rect 31478 24760 31484 24772
rect 31536 24760 31542 24812
rect 32861 24803 32919 24809
rect 32861 24800 32873 24803
rect 32324 24772 32873 24800
rect 31570 24732 31576 24744
rect 27724 24704 31576 24732
rect 31570 24692 31576 24704
rect 31628 24732 31634 24744
rect 32324 24732 32352 24772
rect 32861 24769 32873 24772
rect 32907 24769 32919 24803
rect 32861 24763 32919 24769
rect 33045 24803 33103 24809
rect 33045 24769 33057 24803
rect 33091 24800 33103 24803
rect 33502 24800 33508 24812
rect 33091 24772 33364 24800
rect 33463 24772 33508 24800
rect 33091 24769 33103 24772
rect 33045 24763 33103 24769
rect 31628 24704 32352 24732
rect 32677 24735 32735 24741
rect 31628 24692 31634 24704
rect 32677 24701 32689 24735
rect 32723 24732 32735 24735
rect 33226 24732 33232 24744
rect 32723 24704 33232 24732
rect 32723 24701 32735 24704
rect 32677 24695 32735 24701
rect 33226 24692 33232 24704
rect 33284 24692 33290 24744
rect 33336 24732 33364 24772
rect 33502 24760 33508 24772
rect 33560 24760 33566 24812
rect 33689 24803 33747 24809
rect 33689 24769 33701 24803
rect 33735 24769 33747 24803
rect 33689 24763 33747 24769
rect 34701 24803 34759 24809
rect 34701 24769 34713 24803
rect 34747 24800 34759 24803
rect 34790 24800 34796 24812
rect 34747 24772 34796 24800
rect 34747 24769 34759 24772
rect 34701 24763 34759 24769
rect 33704 24732 33732 24763
rect 34790 24760 34796 24772
rect 34848 24800 34854 24812
rect 36906 24800 36912 24812
rect 34848 24772 36912 24800
rect 34848 24760 34854 24772
rect 36906 24760 36912 24772
rect 36964 24760 36970 24812
rect 34606 24732 34612 24744
rect 33336 24704 34612 24732
rect 34606 24692 34612 24704
rect 34664 24692 34670 24744
rect 35526 24692 35532 24744
rect 35584 24732 35590 24744
rect 37277 24735 37335 24741
rect 37277 24732 37289 24735
rect 35584 24704 37289 24732
rect 35584 24692 35590 24704
rect 37277 24701 37289 24704
rect 37323 24701 37335 24735
rect 37458 24732 37464 24744
rect 37419 24704 37464 24732
rect 37277 24695 37335 24701
rect 37458 24692 37464 24704
rect 37516 24692 37522 24744
rect 38470 24732 38476 24744
rect 38431 24704 38476 24732
rect 38470 24692 38476 24704
rect 38528 24692 38534 24744
rect 38672 24732 38700 24840
rect 38856 24840 44824 24868
rect 38856 24732 38884 24840
rect 44818 24828 44824 24840
rect 44876 24828 44882 24880
rect 46198 24868 46204 24880
rect 45204 24840 46204 24868
rect 40034 24800 40040 24812
rect 39995 24772 40040 24800
rect 40034 24760 40040 24772
rect 40092 24760 40098 24812
rect 45204 24809 45232 24840
rect 46198 24828 46204 24840
rect 46256 24828 46262 24880
rect 46566 24828 46572 24880
rect 46624 24868 46630 24880
rect 46750 24868 46756 24880
rect 46624 24840 46756 24868
rect 46624 24828 46630 24840
rect 46750 24828 46756 24840
rect 46808 24828 46814 24880
rect 47026 24868 47032 24880
rect 46987 24840 47032 24868
rect 47026 24828 47032 24840
rect 47084 24828 47090 24880
rect 45189 24803 45247 24809
rect 45189 24769 45201 24803
rect 45235 24769 45247 24803
rect 45189 24763 45247 24769
rect 47486 24760 47492 24812
rect 47544 24800 47550 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47544 24772 47593 24800
rect 47544 24760 47550 24772
rect 47581 24769 47593 24772
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 38672 24704 38884 24732
rect 45373 24735 45431 24741
rect 45373 24701 45385 24735
rect 45419 24732 45431 24735
rect 46566 24732 46572 24744
rect 45419 24704 46572 24732
rect 45419 24701 45431 24704
rect 45373 24695 45431 24701
rect 46566 24692 46572 24704
rect 46624 24692 46630 24744
rect 19334 24664 19340 24676
rect 13832 24636 15148 24664
rect 15488 24636 19340 24664
rect 11790 24596 11796 24608
rect 11751 24568 11796 24596
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 13446 24556 13452 24608
rect 13504 24596 13510 24608
rect 13832 24596 13860 24636
rect 13504 24568 13860 24596
rect 13504 24556 13510 24568
rect 14366 24556 14372 24608
rect 14424 24596 14430 24608
rect 15488 24596 15516 24636
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 23290 24664 23296 24676
rect 22066 24636 23296 24664
rect 15838 24596 15844 24608
rect 14424 24568 15516 24596
rect 15799 24568 15844 24596
rect 14424 24556 14430 24568
rect 15838 24556 15844 24568
rect 15896 24556 15902 24608
rect 16758 24596 16764 24608
rect 16719 24568 16764 24596
rect 16758 24556 16764 24568
rect 16816 24556 16822 24608
rect 18322 24596 18328 24608
rect 18235 24568 18328 24596
rect 18322 24556 18328 24568
rect 18380 24596 18386 24608
rect 22066 24596 22094 24636
rect 23290 24624 23296 24636
rect 23348 24624 23354 24676
rect 27890 24624 27896 24676
rect 27948 24664 27954 24676
rect 46382 24664 46388 24676
rect 27948 24636 46388 24664
rect 27948 24624 27954 24636
rect 46382 24624 46388 24636
rect 46440 24624 46446 24676
rect 18380 24568 22094 24596
rect 27801 24599 27859 24605
rect 18380 24556 18386 24568
rect 27801 24565 27813 24599
rect 27847 24596 27859 24599
rect 28258 24596 28264 24608
rect 27847 24568 28264 24596
rect 27847 24565 27859 24568
rect 27801 24559 27859 24565
rect 28258 24556 28264 24568
rect 28316 24556 28322 24608
rect 30742 24556 30748 24608
rect 30800 24596 30806 24608
rect 31205 24599 31263 24605
rect 31205 24596 31217 24599
rect 30800 24568 31217 24596
rect 30800 24556 30806 24568
rect 31205 24565 31217 24568
rect 31251 24565 31263 24599
rect 31205 24559 31263 24565
rect 33505 24599 33563 24605
rect 33505 24565 33517 24599
rect 33551 24596 33563 24599
rect 33962 24596 33968 24608
rect 33551 24568 33968 24596
rect 33551 24565 33563 24568
rect 33505 24559 33563 24565
rect 33962 24556 33968 24568
rect 34020 24556 34026 24608
rect 35069 24599 35127 24605
rect 35069 24565 35081 24599
rect 35115 24596 35127 24599
rect 35434 24596 35440 24608
rect 35115 24568 35440 24596
rect 35115 24565 35127 24568
rect 35069 24559 35127 24565
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 37826 24556 37832 24608
rect 37884 24596 37890 24608
rect 40034 24596 40040 24608
rect 37884 24568 40040 24596
rect 37884 24556 37890 24568
rect 40034 24556 40040 24568
rect 40092 24556 40098 24608
rect 46474 24556 46480 24608
rect 46532 24596 46538 24608
rect 47673 24599 47731 24605
rect 47673 24596 47685 24599
rect 46532 24568 47685 24596
rect 46532 24556 46538 24568
rect 47673 24565 47685 24568
rect 47719 24565 47731 24599
rect 47673 24559 47731 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 12066 24352 12072 24404
rect 12124 24392 12130 24404
rect 15930 24392 15936 24404
rect 12124 24364 15936 24392
rect 12124 24352 12130 24364
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 16022 24352 16028 24404
rect 16080 24392 16086 24404
rect 16761 24395 16819 24401
rect 16761 24392 16773 24395
rect 16080 24364 16773 24392
rect 16080 24352 16086 24364
rect 16761 24361 16773 24364
rect 16807 24361 16819 24395
rect 16761 24355 16819 24361
rect 17310 24352 17316 24404
rect 17368 24392 17374 24404
rect 22462 24392 22468 24404
rect 17368 24364 22468 24392
rect 17368 24352 17374 24364
rect 22462 24352 22468 24364
rect 22520 24392 22526 24404
rect 46014 24392 46020 24404
rect 22520 24364 23612 24392
rect 22520 24352 22526 24364
rect 19334 24284 19340 24336
rect 19392 24324 19398 24336
rect 19981 24327 20039 24333
rect 19981 24324 19993 24327
rect 19392 24296 19993 24324
rect 19392 24284 19398 24296
rect 19981 24293 19993 24296
rect 20027 24293 20039 24327
rect 19981 24287 20039 24293
rect 20717 24327 20775 24333
rect 20717 24293 20729 24327
rect 20763 24324 20775 24327
rect 22186 24324 22192 24336
rect 20763 24296 22192 24324
rect 20763 24293 20775 24296
rect 20717 24287 20775 24293
rect 22186 24284 22192 24296
rect 22244 24284 22250 24336
rect 11790 24256 11796 24268
rect 11751 24228 11796 24256
rect 11790 24216 11796 24228
rect 11848 24216 11854 24268
rect 15013 24259 15071 24265
rect 15013 24225 15025 24259
rect 15059 24256 15071 24259
rect 15838 24256 15844 24268
rect 15059 24228 15844 24256
rect 15059 24225 15071 24228
rect 15013 24219 15071 24225
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 20530 24256 20536 24268
rect 17920 24228 20536 24256
rect 17920 24216 17926 24228
rect 20530 24216 20536 24228
rect 20588 24256 20594 24268
rect 23584 24256 23612 24364
rect 28828 24364 46020 24392
rect 24302 24284 24308 24336
rect 24360 24324 24366 24336
rect 27890 24324 27896 24336
rect 24360 24296 27896 24324
rect 24360 24284 24366 24296
rect 27890 24284 27896 24296
rect 27948 24284 27954 24336
rect 28828 24265 28856 24364
rect 46014 24352 46020 24364
rect 46072 24352 46078 24404
rect 33226 24324 33232 24336
rect 33187 24296 33232 24324
rect 33226 24284 33232 24296
rect 33284 24284 33290 24336
rect 36906 24324 36912 24336
rect 36867 24296 36912 24324
rect 36906 24284 36912 24296
rect 36964 24284 36970 24336
rect 47762 24324 47768 24336
rect 46308 24296 47768 24324
rect 28813 24259 28871 24265
rect 20588 24228 20760 24256
rect 23584 24228 26372 24256
rect 20588 24216 20594 24228
rect 13354 24148 13360 24200
rect 13412 24188 13418 24200
rect 14366 24188 14372 24200
rect 13412 24160 14372 24188
rect 13412 24148 13418 24160
rect 14366 24148 14372 24160
rect 14424 24148 14430 24200
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24157 14611 24191
rect 16758 24188 16764 24200
rect 16422 24160 16764 24188
rect 14553 24151 14611 24157
rect 12066 24120 12072 24132
rect 12027 24092 12072 24120
rect 12066 24080 12072 24092
rect 12124 24080 12130 24132
rect 13998 24120 14004 24132
rect 13294 24092 14004 24120
rect 13998 24080 14004 24092
rect 14056 24080 14062 24132
rect 14568 24120 14596 24151
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24188 17371 24191
rect 17402 24188 17408 24200
rect 17359 24160 17408 24188
rect 17359 24157 17371 24160
rect 17313 24151 17371 24157
rect 17402 24148 17408 24160
rect 17460 24188 17466 24200
rect 18322 24188 18328 24200
rect 17460 24160 18328 24188
rect 17460 24148 17466 24160
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24188 19855 24191
rect 20070 24188 20076 24200
rect 19843 24160 20076 24188
rect 19843 24157 19855 24160
rect 19797 24151 19855 24157
rect 15194 24120 15200 24132
rect 14568 24092 15200 24120
rect 15194 24080 15200 24092
rect 15252 24080 15258 24132
rect 15289 24123 15347 24129
rect 15289 24089 15301 24123
rect 15335 24120 15347 24123
rect 15378 24120 15384 24132
rect 15335 24092 15384 24120
rect 15335 24089 15347 24092
rect 15289 24083 15347 24089
rect 15378 24080 15384 24092
rect 15436 24080 15442 24132
rect 19720 24120 19748 24151
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20732 24197 20760 24228
rect 20717 24191 20775 24197
rect 20717 24157 20729 24191
rect 20763 24157 20775 24191
rect 20990 24188 20996 24200
rect 20951 24160 20996 24188
rect 20717 24151 20775 24157
rect 20990 24148 20996 24160
rect 21048 24148 21054 24200
rect 21450 24188 21456 24200
rect 21411 24160 21456 24188
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 24762 24148 24768 24200
rect 24820 24188 24826 24200
rect 26344 24197 26372 24228
rect 28813 24225 28825 24259
rect 28859 24225 28871 24259
rect 30742 24256 30748 24268
rect 30703 24228 30748 24256
rect 28813 24219 28871 24225
rect 30742 24216 30748 24228
rect 30800 24216 30806 24268
rect 35434 24256 35440 24268
rect 35395 24228 35440 24256
rect 35434 24216 35440 24228
rect 35492 24216 35498 24268
rect 35802 24216 35808 24268
rect 35860 24256 35866 24268
rect 37461 24259 37519 24265
rect 37461 24256 37473 24259
rect 35860 24228 37473 24256
rect 35860 24216 35866 24228
rect 37461 24225 37473 24228
rect 37507 24225 37519 24259
rect 40310 24256 40316 24268
rect 40271 24228 40316 24256
rect 37461 24219 37519 24225
rect 40310 24216 40316 24228
rect 40368 24216 40374 24268
rect 46308 24265 46336 24296
rect 47762 24284 47768 24296
rect 47820 24284 47826 24336
rect 46293 24259 46351 24265
rect 46293 24225 46305 24259
rect 46339 24225 46351 24259
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 46293 24219 46351 24225
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 25317 24191 25375 24197
rect 25317 24188 25329 24191
rect 24820 24160 25329 24188
rect 24820 24148 24826 24160
rect 25317 24157 25329 24160
rect 25363 24157 25375 24191
rect 25317 24151 25375 24157
rect 26329 24191 26387 24197
rect 26329 24157 26341 24191
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 26510 24148 26516 24200
rect 26568 24188 26574 24200
rect 26973 24191 27031 24197
rect 26973 24188 26985 24191
rect 26568 24160 26985 24188
rect 26568 24148 26574 24160
rect 26973 24157 26985 24160
rect 27019 24157 27031 24191
rect 29546 24188 29552 24200
rect 29507 24160 29552 24188
rect 26973 24151 27031 24157
rect 29546 24148 29552 24160
rect 29604 24148 29610 24200
rect 30466 24188 30472 24200
rect 30427 24160 30472 24188
rect 30466 24148 30472 24160
rect 30524 24148 30530 24200
rect 32861 24191 32919 24197
rect 32861 24157 32873 24191
rect 32907 24188 32919 24191
rect 32950 24188 32956 24200
rect 32907 24160 32956 24188
rect 32907 24157 32919 24160
rect 32861 24151 32919 24157
rect 32950 24148 32956 24160
rect 33008 24148 33014 24200
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 34514 24188 34520 24200
rect 34011 24160 34520 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 34514 24148 34520 24160
rect 34572 24148 34578 24200
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 35161 24191 35219 24197
rect 35161 24188 35173 24191
rect 34848 24160 35173 24188
rect 34848 24148 34854 24160
rect 35161 24157 35173 24160
rect 35207 24157 35219 24191
rect 39850 24188 39856 24200
rect 39811 24160 39856 24188
rect 35161 24151 35219 24157
rect 39850 24148 39856 24160
rect 39908 24148 39914 24200
rect 20346 24120 20352 24132
rect 19720 24092 20352 24120
rect 20346 24080 20352 24092
rect 20404 24080 20410 24132
rect 26421 24123 26479 24129
rect 26421 24089 26433 24123
rect 26467 24120 26479 24123
rect 27157 24123 27215 24129
rect 27157 24120 27169 24123
rect 26467 24092 27169 24120
rect 26467 24089 26479 24092
rect 26421 24083 26479 24089
rect 27157 24089 27169 24092
rect 27203 24089 27215 24123
rect 27157 24083 27215 24089
rect 31754 24080 31760 24132
rect 31812 24080 31818 24132
rect 32674 24120 32680 24132
rect 32635 24092 32680 24120
rect 32674 24080 32680 24092
rect 32732 24080 32738 24132
rect 32766 24080 32772 24132
rect 32824 24120 32830 24132
rect 33045 24123 33103 24129
rect 33045 24120 33057 24123
rect 32824 24092 33057 24120
rect 32824 24080 32830 24092
rect 33045 24089 33057 24092
rect 33091 24089 33103 24123
rect 33045 24083 33103 24089
rect 33796 24092 34192 24120
rect 12342 24012 12348 24064
rect 12400 24052 12406 24064
rect 13541 24055 13599 24061
rect 13541 24052 13553 24055
rect 12400 24024 13553 24052
rect 12400 24012 12406 24024
rect 13541 24021 13553 24024
rect 13587 24052 13599 24055
rect 14090 24052 14096 24064
rect 13587 24024 14096 24052
rect 13587 24021 13599 24024
rect 13541 24015 13599 24021
rect 14090 24012 14096 24024
rect 14148 24012 14154 24064
rect 14553 24055 14611 24061
rect 14553 24021 14565 24055
rect 14599 24052 14611 24055
rect 15654 24052 15660 24064
rect 14599 24024 15660 24052
rect 14599 24021 14611 24024
rect 14553 24015 14611 24021
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 17126 24012 17132 24064
rect 17184 24052 17190 24064
rect 17497 24055 17555 24061
rect 17497 24052 17509 24055
rect 17184 24024 17509 24052
rect 17184 24012 17190 24024
rect 17497 24021 17509 24024
rect 17543 24052 17555 24055
rect 18322 24052 18328 24064
rect 17543 24024 18328 24052
rect 17543 24021 17555 24024
rect 17497 24015 17555 24021
rect 18322 24012 18328 24024
rect 18380 24012 18386 24064
rect 20806 24012 20812 24064
rect 20864 24052 20870 24064
rect 20901 24055 20959 24061
rect 20901 24052 20913 24055
rect 20864 24024 20913 24052
rect 20864 24012 20870 24024
rect 20901 24021 20913 24024
rect 20947 24021 20959 24055
rect 20901 24015 20959 24021
rect 21637 24055 21695 24061
rect 21637 24021 21649 24055
rect 21683 24052 21695 24055
rect 21818 24052 21824 24064
rect 21683 24024 21824 24052
rect 21683 24021 21695 24024
rect 21637 24015 21695 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 25406 24052 25412 24064
rect 25367 24024 25412 24052
rect 25406 24012 25412 24024
rect 25464 24012 25470 24064
rect 29638 24052 29644 24064
rect 29599 24024 29644 24052
rect 29638 24012 29644 24024
rect 29696 24012 29702 24064
rect 32122 24012 32128 24064
rect 32180 24052 32186 24064
rect 32217 24055 32275 24061
rect 32217 24052 32229 24055
rect 32180 24024 32229 24052
rect 32180 24012 32186 24024
rect 32217 24021 32229 24024
rect 32263 24052 32275 24055
rect 32953 24055 33011 24061
rect 32953 24052 32965 24055
rect 32263 24024 32965 24052
rect 32263 24021 32275 24024
rect 32217 24015 32275 24021
rect 32953 24021 32965 24024
rect 32999 24052 33011 24055
rect 33796 24052 33824 24092
rect 34054 24052 34060 24064
rect 32999 24024 33824 24052
rect 34015 24024 34060 24052
rect 32999 24021 33011 24024
rect 32953 24015 33011 24021
rect 34054 24012 34060 24024
rect 34112 24012 34118 24064
rect 34164 24052 34192 24092
rect 35986 24080 35992 24132
rect 36044 24080 36050 24132
rect 37642 24120 37648 24132
rect 37603 24092 37648 24120
rect 37642 24080 37648 24092
rect 37700 24080 37706 24132
rect 39298 24120 39304 24132
rect 39259 24092 39304 24120
rect 39298 24080 39304 24092
rect 39356 24080 39362 24132
rect 40034 24120 40040 24132
rect 39995 24092 40040 24120
rect 40034 24080 40040 24092
rect 40092 24080 40098 24132
rect 36078 24052 36084 24064
rect 34164 24024 36084 24052
rect 36078 24012 36084 24024
rect 36136 24012 36142 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1949 23851 2007 23857
rect 1949 23817 1961 23851
rect 1995 23848 2007 23851
rect 1995 23820 6914 23848
rect 1995 23817 2007 23820
rect 1949 23811 2007 23817
rect 6886 23780 6914 23820
rect 11698 23808 11704 23860
rect 11756 23848 11762 23860
rect 12069 23851 12127 23857
rect 12069 23848 12081 23851
rect 11756 23820 12081 23848
rect 11756 23808 11762 23820
rect 12069 23817 12081 23820
rect 12115 23848 12127 23851
rect 13446 23848 13452 23860
rect 12115 23820 13216 23848
rect 13407 23820 13452 23848
rect 12115 23817 12127 23820
rect 12069 23811 12127 23817
rect 12986 23780 12992 23792
rect 6886 23752 12992 23780
rect 12986 23740 12992 23752
rect 13044 23740 13050 23792
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 11974 23712 11980 23724
rect 11935 23684 11980 23712
rect 11974 23672 11980 23684
rect 12032 23672 12038 23724
rect 12342 23712 12348 23724
rect 12084 23684 12348 23712
rect 11606 23604 11612 23656
rect 11664 23644 11670 23656
rect 12084 23644 12112 23684
rect 12342 23672 12348 23684
rect 12400 23712 12406 23724
rect 13188 23721 13216 23820
rect 13446 23808 13452 23820
rect 13504 23808 13510 23860
rect 13998 23848 14004 23860
rect 13959 23820 14004 23848
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 14090 23808 14096 23860
rect 14148 23848 14154 23860
rect 14737 23851 14795 23857
rect 14737 23848 14749 23851
rect 14148 23820 14749 23848
rect 14148 23808 14154 23820
rect 14737 23817 14749 23820
rect 14783 23817 14795 23851
rect 14737 23811 14795 23817
rect 15105 23851 15163 23857
rect 15105 23817 15117 23851
rect 15151 23848 15163 23851
rect 15194 23848 15200 23860
rect 15151 23820 15200 23848
rect 15151 23817 15163 23820
rect 15105 23811 15163 23817
rect 15194 23808 15200 23820
rect 15252 23808 15258 23860
rect 20806 23848 20812 23860
rect 20767 23820 20812 23848
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 20993 23851 21051 23857
rect 20993 23817 21005 23851
rect 21039 23848 21051 23851
rect 21358 23848 21364 23860
rect 21039 23820 21364 23848
rect 21039 23817 21051 23820
rect 20993 23811 21051 23817
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 23569 23851 23627 23857
rect 23569 23848 23581 23851
rect 22066 23820 23581 23848
rect 14553 23783 14611 23789
rect 14553 23749 14565 23783
rect 14599 23780 14611 23783
rect 15010 23780 15016 23792
rect 14599 23752 15016 23780
rect 14599 23749 14611 23752
rect 14553 23743 14611 23749
rect 15010 23740 15016 23752
rect 15068 23740 15074 23792
rect 20441 23783 20499 23789
rect 20441 23749 20453 23783
rect 20487 23780 20499 23783
rect 20530 23780 20536 23792
rect 20487 23752 20536 23780
rect 20487 23749 20499 23752
rect 20441 23743 20499 23749
rect 20530 23740 20536 23752
rect 20588 23780 20594 23792
rect 22066 23780 22094 23820
rect 23569 23817 23581 23820
rect 23615 23817 23627 23851
rect 23569 23811 23627 23817
rect 26786 23808 26792 23860
rect 26844 23848 26850 23860
rect 29733 23851 29791 23857
rect 29733 23848 29745 23851
rect 26844 23820 29745 23848
rect 26844 23808 26850 23820
rect 29733 23817 29745 23820
rect 29779 23817 29791 23851
rect 30466 23848 30472 23860
rect 30427 23820 30472 23848
rect 29733 23811 29791 23817
rect 28258 23780 28264 23792
rect 20588 23752 22094 23780
rect 28219 23752 28264 23780
rect 20588 23740 20594 23752
rect 28258 23740 28264 23752
rect 28316 23740 28322 23792
rect 29638 23780 29644 23792
rect 29486 23752 29644 23780
rect 29638 23740 29644 23752
rect 29696 23740 29702 23792
rect 29748 23780 29776 23811
rect 30466 23808 30472 23820
rect 30524 23808 30530 23860
rect 33051 23851 33109 23857
rect 33051 23817 33063 23851
rect 33097 23848 33109 23851
rect 33502 23848 33508 23860
rect 33097 23820 33508 23848
rect 33097 23817 33109 23820
rect 33051 23811 33109 23817
rect 33502 23808 33508 23820
rect 33560 23808 33566 23860
rect 35437 23851 35495 23857
rect 35437 23848 35449 23851
rect 33796 23820 35449 23848
rect 31297 23783 31355 23789
rect 29748 23752 30512 23780
rect 12897 23715 12955 23721
rect 12897 23712 12909 23715
rect 12400 23684 12909 23712
rect 12400 23672 12406 23684
rect 12897 23681 12909 23684
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 13173 23715 13231 23721
rect 13173 23681 13185 23715
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13354 23712 13360 23724
rect 13311 23684 13360 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 11664 23616 12112 23644
rect 12161 23647 12219 23653
rect 11664 23604 11670 23616
rect 12161 23613 12173 23647
rect 12207 23644 12219 23647
rect 13096 23644 13124 23675
rect 12207 23616 13124 23644
rect 13188 23644 13216 23675
rect 13354 23672 13360 23684
rect 13412 23672 13418 23724
rect 13906 23712 13912 23724
rect 13867 23684 13912 23712
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 14274 23672 14280 23724
rect 14332 23712 14338 23724
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 14332 23684 14841 23712
rect 14332 23672 14338 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 14921 23715 14979 23721
rect 14921 23681 14933 23715
rect 14967 23681 14979 23715
rect 14921 23675 14979 23681
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23712 15807 23715
rect 16942 23712 16948 23724
rect 15795 23684 16948 23712
rect 15795 23681 15807 23684
rect 15749 23675 15807 23681
rect 13722 23644 13728 23656
rect 13188 23616 13728 23644
rect 12207 23613 12219 23616
rect 12161 23607 12219 23613
rect 13096 23576 13124 23616
rect 13722 23604 13728 23616
rect 13780 23644 13786 23656
rect 14936 23644 14964 23675
rect 16942 23672 16948 23684
rect 17000 23672 17006 23724
rect 17126 23712 17132 23724
rect 17087 23684 17132 23712
rect 17126 23672 17132 23684
rect 17184 23672 17190 23724
rect 19610 23672 19616 23724
rect 19668 23712 19674 23724
rect 19705 23715 19763 23721
rect 19705 23712 19717 23715
rect 19668 23684 19717 23712
rect 19668 23672 19674 23684
rect 19705 23681 19717 23684
rect 19751 23681 19763 23715
rect 19886 23712 19892 23724
rect 19847 23684 19892 23712
rect 19705 23675 19763 23681
rect 19886 23672 19892 23684
rect 19944 23672 19950 23724
rect 19978 23672 19984 23724
rect 20036 23712 20042 23724
rect 20622 23712 20628 23724
rect 20036 23684 20081 23712
rect 20583 23684 20628 23712
rect 20036 23672 20042 23684
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 21818 23712 21824 23724
rect 20772 23684 20817 23712
rect 21779 23684 21824 23712
rect 20772 23672 20778 23684
rect 21818 23672 21824 23684
rect 21876 23672 21882 23724
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23712 25835 23715
rect 25866 23712 25872 23724
rect 25823 23684 25872 23712
rect 25823 23681 25835 23684
rect 25777 23675 25835 23681
rect 25866 23672 25872 23684
rect 25924 23672 25930 23724
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23712 27491 23715
rect 27890 23712 27896 23724
rect 27479 23684 27896 23712
rect 27479 23681 27491 23684
rect 27433 23675 27491 23681
rect 27890 23672 27896 23684
rect 27948 23672 27954 23724
rect 30377 23715 30435 23721
rect 30377 23681 30389 23715
rect 30423 23681 30435 23715
rect 30484 23712 30512 23752
rect 31297 23749 31309 23783
rect 31343 23780 31355 23783
rect 32122 23780 32128 23792
rect 31343 23752 32128 23780
rect 31343 23749 31355 23752
rect 31297 23743 31355 23749
rect 32122 23740 32128 23752
rect 32180 23740 32186 23792
rect 32325 23783 32383 23789
rect 32325 23780 32337 23783
rect 32232 23752 32337 23780
rect 31481 23715 31539 23721
rect 31481 23712 31493 23715
rect 30484 23684 31493 23712
rect 30377 23675 30435 23681
rect 15654 23644 15660 23656
rect 13780 23616 14964 23644
rect 15615 23616 15660 23644
rect 13780 23604 13786 23616
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 16022 23604 16028 23656
rect 16080 23644 16086 23656
rect 21450 23644 21456 23656
rect 16080 23616 21456 23644
rect 16080 23604 16086 23616
rect 21450 23604 21456 23616
rect 21508 23604 21514 23656
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 27525 23647 27583 23653
rect 22152 23616 22197 23644
rect 22152 23604 22158 23616
rect 27525 23613 27537 23647
rect 27571 23644 27583 23647
rect 27985 23647 28043 23653
rect 27985 23644 27997 23647
rect 27571 23616 27997 23644
rect 27571 23613 27583 23616
rect 27525 23607 27583 23613
rect 27985 23613 27997 23616
rect 28031 23613 28043 23647
rect 30392 23644 30420 23675
rect 30834 23644 30840 23656
rect 27985 23607 28043 23613
rect 28092 23616 30840 23644
rect 14274 23576 14280 23588
rect 13096 23548 14280 23576
rect 14274 23536 14280 23548
rect 14332 23536 14338 23588
rect 16117 23579 16175 23585
rect 16117 23545 16129 23579
rect 16163 23576 16175 23579
rect 16390 23576 16396 23588
rect 16163 23548 16396 23576
rect 16163 23545 16175 23548
rect 16117 23539 16175 23545
rect 16390 23536 16396 23548
rect 16448 23536 16454 23588
rect 18046 23576 18052 23588
rect 16500 23548 18052 23576
rect 12342 23508 12348 23520
rect 12303 23480 12348 23508
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 16500 23508 16528 23548
rect 18046 23536 18052 23548
rect 18104 23536 18110 23588
rect 27890 23536 27896 23588
rect 27948 23576 27954 23588
rect 28092 23576 28120 23616
rect 30834 23604 30840 23616
rect 30892 23604 30898 23656
rect 31294 23576 31300 23588
rect 27948 23548 28120 23576
rect 31255 23548 31300 23576
rect 27948 23536 27954 23548
rect 31294 23536 31300 23548
rect 31352 23536 31358 23588
rect 13044 23480 16528 23508
rect 13044 23468 13050 23480
rect 17126 23468 17132 23520
rect 17184 23508 17190 23520
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 17184 23480 17233 23508
rect 17184 23468 17190 23480
rect 17221 23477 17233 23480
rect 17267 23477 17279 23511
rect 19518 23508 19524 23520
rect 19479 23480 19524 23508
rect 17221 23471 17279 23477
rect 19518 23468 19524 23480
rect 19576 23468 19582 23520
rect 25222 23468 25228 23520
rect 25280 23508 25286 23520
rect 25961 23511 26019 23517
rect 25961 23508 25973 23511
rect 25280 23480 25973 23508
rect 25280 23468 25286 23480
rect 25961 23477 25973 23480
rect 26007 23477 26019 23511
rect 31404 23508 31432 23684
rect 31481 23681 31493 23684
rect 31527 23681 31539 23715
rect 31481 23675 31539 23681
rect 31570 23672 31576 23724
rect 31628 23712 31634 23724
rect 32232 23712 32260 23752
rect 32325 23749 32337 23752
rect 32371 23749 32383 23783
rect 32325 23743 32383 23749
rect 32674 23740 32680 23792
rect 32732 23780 32738 23792
rect 32953 23783 33011 23789
rect 32953 23780 32965 23783
rect 32732 23752 32965 23780
rect 32732 23740 32738 23752
rect 32953 23749 32965 23752
rect 32999 23780 33011 23783
rect 33796 23780 33824 23820
rect 35437 23817 35449 23820
rect 35483 23848 35495 23851
rect 35526 23848 35532 23860
rect 35483 23820 35532 23848
rect 35483 23817 35495 23820
rect 35437 23811 35495 23817
rect 35526 23808 35532 23820
rect 35584 23808 35590 23860
rect 35986 23848 35992 23860
rect 35947 23820 35992 23848
rect 35986 23808 35992 23820
rect 36044 23808 36050 23860
rect 37553 23851 37611 23857
rect 37553 23817 37565 23851
rect 37599 23848 37611 23851
rect 37642 23848 37648 23860
rect 37599 23820 37648 23848
rect 37599 23817 37611 23820
rect 37553 23811 37611 23817
rect 37642 23808 37648 23820
rect 37700 23808 37706 23860
rect 39301 23851 39359 23857
rect 39301 23817 39313 23851
rect 39347 23848 39359 23851
rect 40034 23848 40040 23860
rect 39347 23820 40040 23848
rect 39347 23817 39359 23820
rect 39301 23811 39359 23817
rect 40034 23808 40040 23820
rect 40092 23808 40098 23860
rect 46566 23808 46572 23860
rect 46624 23848 46630 23860
rect 47673 23851 47731 23857
rect 47673 23848 47685 23851
rect 46624 23820 47685 23848
rect 46624 23808 46630 23820
rect 47673 23817 47685 23820
rect 47719 23817 47731 23851
rect 47673 23811 47731 23817
rect 33962 23780 33968 23792
rect 32999 23752 33824 23780
rect 33923 23752 33968 23780
rect 32999 23749 33011 23752
rect 32953 23743 33011 23749
rect 33962 23740 33968 23752
rect 34020 23740 34026 23792
rect 34054 23740 34060 23792
rect 34112 23780 34118 23792
rect 44910 23780 44916 23792
rect 34112 23752 34454 23780
rect 41386 23752 44916 23780
rect 34112 23740 34118 23752
rect 31628 23684 32260 23712
rect 31628 23672 31634 23684
rect 33042 23672 33048 23724
rect 33100 23712 33106 23724
rect 33137 23715 33195 23721
rect 33137 23712 33149 23715
rect 33100 23684 33149 23712
rect 33100 23672 33106 23684
rect 33137 23681 33149 23684
rect 33183 23681 33195 23715
rect 33137 23675 33195 23681
rect 33229 23715 33287 23721
rect 33229 23681 33241 23715
rect 33275 23681 33287 23715
rect 33229 23675 33287 23681
rect 35897 23715 35955 23721
rect 35897 23681 35909 23715
rect 35943 23681 35955 23715
rect 37458 23712 37464 23724
rect 37419 23684 37464 23712
rect 35897 23675 35955 23681
rect 31478 23536 31484 23588
rect 31536 23576 31542 23588
rect 32493 23579 32551 23585
rect 32493 23576 32505 23579
rect 31536 23548 32505 23576
rect 31536 23536 31542 23548
rect 32493 23545 32505 23548
rect 32539 23576 32551 23579
rect 33244 23576 33272 23675
rect 33686 23644 33692 23656
rect 33647 23616 33692 23644
rect 33686 23604 33692 23616
rect 33744 23604 33750 23656
rect 34514 23604 34520 23656
rect 34572 23644 34578 23656
rect 35912 23644 35940 23675
rect 37458 23672 37464 23684
rect 37516 23672 37522 23724
rect 39206 23712 39212 23724
rect 39167 23684 39212 23712
rect 39206 23672 39212 23684
rect 39264 23712 39270 23724
rect 41386 23712 41414 23752
rect 44910 23740 44916 23752
rect 44968 23740 44974 23792
rect 39264 23684 41414 23712
rect 42797 23715 42855 23721
rect 39264 23672 39270 23684
rect 42797 23681 42809 23715
rect 42843 23681 42855 23715
rect 42978 23712 42984 23724
rect 42939 23684 42984 23712
rect 42797 23675 42855 23681
rect 34572 23616 35940 23644
rect 42812 23644 42840 23675
rect 42978 23672 42984 23684
rect 43036 23672 43042 23724
rect 45925 23715 45983 23721
rect 45925 23681 45937 23715
rect 45971 23681 45983 23715
rect 47026 23712 47032 23724
rect 46987 23684 47032 23712
rect 45925 23675 45983 23681
rect 43438 23644 43444 23656
rect 42812 23616 43444 23644
rect 34572 23604 34578 23616
rect 43438 23604 43444 23616
rect 43496 23604 43502 23656
rect 45940 23644 45968 23675
rect 47026 23672 47032 23684
rect 47084 23672 47090 23724
rect 47578 23712 47584 23724
rect 47539 23684 47584 23712
rect 47578 23672 47584 23684
rect 47636 23672 47642 23724
rect 48038 23644 48044 23656
rect 45940 23616 48044 23644
rect 48038 23604 48044 23616
rect 48096 23604 48102 23656
rect 32539 23548 33272 23576
rect 32539 23545 32551 23548
rect 32493 23539 32551 23545
rect 32309 23511 32367 23517
rect 32309 23508 32321 23511
rect 31404 23480 32321 23508
rect 25961 23471 26019 23477
rect 32309 23477 32321 23480
rect 32355 23508 32367 23511
rect 32766 23508 32772 23520
rect 32355 23480 32772 23508
rect 32355 23477 32367 23480
rect 32309 23471 32367 23477
rect 32766 23468 32772 23480
rect 32824 23468 32830 23520
rect 33778 23468 33784 23520
rect 33836 23508 33842 23520
rect 37826 23508 37832 23520
rect 33836 23480 37832 23508
rect 33836 23468 33842 23480
rect 37826 23468 37832 23480
rect 37884 23468 37890 23520
rect 42794 23508 42800 23520
rect 42755 23480 42800 23508
rect 42794 23468 42800 23480
rect 42852 23468 42858 23520
rect 45738 23508 45744 23520
rect 45699 23480 45744 23508
rect 45738 23468 45744 23480
rect 45796 23468 45802 23520
rect 46566 23468 46572 23520
rect 46624 23508 46630 23520
rect 46845 23511 46903 23517
rect 46845 23508 46857 23511
rect 46624 23480 46857 23508
rect 46624 23468 46630 23480
rect 46845 23477 46857 23480
rect 46891 23477 46903 23511
rect 46845 23471 46903 23477
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 12066 23264 12072 23316
rect 12124 23304 12130 23316
rect 12345 23307 12403 23313
rect 12345 23304 12357 23307
rect 12124 23276 12357 23304
rect 12124 23264 12130 23276
rect 12345 23273 12357 23276
rect 12391 23273 12403 23307
rect 12345 23267 12403 23273
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 16942 23304 16948 23316
rect 16632 23276 16948 23304
rect 16632 23264 16638 23276
rect 16942 23264 16948 23276
rect 17000 23304 17006 23316
rect 17862 23304 17868 23316
rect 17000 23276 17868 23304
rect 17000 23264 17006 23276
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 22094 23264 22100 23316
rect 22152 23304 22158 23316
rect 22189 23307 22247 23313
rect 22189 23304 22201 23307
rect 22152 23276 22201 23304
rect 22152 23264 22158 23276
rect 22189 23273 22201 23276
rect 22235 23273 22247 23307
rect 23198 23304 23204 23316
rect 23159 23276 23204 23304
rect 22189 23267 22247 23273
rect 23198 23264 23204 23276
rect 23256 23264 23262 23316
rect 29546 23304 29552 23316
rect 23952 23276 29552 23304
rect 16022 23168 16028 23180
rect 15580 23140 16028 23168
rect 12342 23100 12348 23112
rect 12303 23072 12348 23100
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 13446 23100 13452 23112
rect 12575 23072 13452 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 15580 23109 15608 23140
rect 16022 23128 16028 23140
rect 16080 23128 16086 23180
rect 16390 23168 16396 23180
rect 16351 23140 16396 23168
rect 16390 23128 16396 23140
rect 16448 23128 16454 23180
rect 19518 23128 19524 23180
rect 19576 23168 19582 23180
rect 20533 23171 20591 23177
rect 20533 23168 20545 23171
rect 19576 23140 20545 23168
rect 19576 23128 19582 23140
rect 20533 23137 20545 23140
rect 20579 23137 20591 23171
rect 20533 23131 20591 23137
rect 23952 23112 23980 23276
rect 29546 23264 29552 23276
rect 29604 23304 29610 23316
rect 29733 23307 29791 23313
rect 29733 23304 29745 23307
rect 29604 23276 29745 23304
rect 29604 23264 29610 23276
rect 29733 23273 29745 23276
rect 29779 23273 29791 23307
rect 29733 23267 29791 23273
rect 31665 23307 31723 23313
rect 31665 23273 31677 23307
rect 31711 23304 31723 23307
rect 31754 23304 31760 23316
rect 31711 23276 31760 23304
rect 31711 23273 31723 23276
rect 31665 23267 31723 23273
rect 24489 23171 24547 23177
rect 24489 23137 24501 23171
rect 24535 23168 24547 23171
rect 27798 23168 27804 23180
rect 24535 23140 27804 23168
rect 24535 23137 24547 23140
rect 24489 23131 24547 23137
rect 27798 23128 27804 23140
rect 27856 23128 27862 23180
rect 27982 23168 27988 23180
rect 27943 23140 27988 23168
rect 27982 23128 27988 23140
rect 28040 23128 28046 23180
rect 15565 23103 15623 23109
rect 15565 23069 15577 23103
rect 15611 23069 15623 23103
rect 15565 23063 15623 23069
rect 15657 23103 15715 23109
rect 15657 23069 15669 23103
rect 15703 23100 15715 23103
rect 16117 23103 16175 23109
rect 16117 23100 16129 23103
rect 15703 23072 16129 23100
rect 15703 23069 15715 23072
rect 15657 23063 15715 23069
rect 16117 23069 16129 23072
rect 16163 23069 16175 23103
rect 18322 23100 18328 23112
rect 18283 23072 18328 23100
rect 16117 23063 16175 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19705 23103 19763 23109
rect 19705 23100 19717 23103
rect 19392 23072 19717 23100
rect 19392 23060 19398 23072
rect 19705 23069 19717 23072
rect 19751 23100 19763 23103
rect 19886 23100 19892 23112
rect 19751 23072 19892 23100
rect 19751 23069 19763 23072
rect 19705 23063 19763 23069
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23100 20131 23103
rect 20806 23100 20812 23112
rect 20119 23072 20812 23100
rect 20119 23069 20131 23072
rect 20073 23063 20131 23069
rect 20806 23060 20812 23072
rect 20864 23100 20870 23112
rect 20901 23103 20959 23109
rect 20901 23100 20913 23103
rect 20864 23072 20913 23100
rect 20864 23060 20870 23072
rect 20901 23069 20913 23072
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 21450 23100 21456 23112
rect 21048 23072 21093 23100
rect 21411 23072 21456 23100
rect 21048 23060 21054 23072
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 22186 23100 22192 23112
rect 22147 23072 22192 23100
rect 22186 23060 22192 23072
rect 22244 23060 22250 23112
rect 22370 23100 22376 23112
rect 22331 23072 22376 23100
rect 22370 23060 22376 23072
rect 22428 23060 22434 23112
rect 23109 23103 23167 23109
rect 23109 23069 23121 23103
rect 23155 23100 23167 23103
rect 23934 23100 23940 23112
rect 23155 23072 23940 23100
rect 23155 23069 23167 23072
rect 23109 23063 23167 23069
rect 23934 23060 23940 23072
rect 23992 23060 23998 23112
rect 26786 23100 26792 23112
rect 26747 23072 26792 23100
rect 26786 23060 26792 23072
rect 26844 23060 26850 23112
rect 29549 23103 29607 23109
rect 29549 23069 29561 23103
rect 29595 23100 29607 23103
rect 29638 23100 29644 23112
rect 29595 23072 29644 23100
rect 29595 23069 29607 23072
rect 29549 23063 29607 23069
rect 17126 22992 17132 23044
rect 17184 22992 17190 23044
rect 19521 23035 19579 23041
rect 19521 23001 19533 23035
rect 19567 23032 19579 23035
rect 19610 23032 19616 23044
rect 19567 23004 19616 23032
rect 19567 23001 19579 23004
rect 19521 22995 19579 23001
rect 19610 22992 19616 23004
rect 19668 23032 19674 23044
rect 20162 23032 20168 23044
rect 19668 23004 20168 23032
rect 19668 22992 19674 23004
rect 20162 22992 20168 23004
rect 20220 22992 20226 23044
rect 24762 23032 24768 23044
rect 24723 23004 24768 23032
rect 24762 22992 24768 23004
rect 24820 22992 24826 23044
rect 25406 22992 25412 23044
rect 25464 22992 25470 23044
rect 26970 23032 26976 23044
rect 26068 23004 26372 23032
rect 26931 23004 26976 23032
rect 18322 22924 18328 22976
rect 18380 22964 18386 22976
rect 18417 22967 18475 22973
rect 18417 22964 18429 22967
rect 18380 22936 18429 22964
rect 18380 22924 18386 22936
rect 18417 22933 18429 22936
rect 18463 22933 18475 22967
rect 18417 22927 18475 22933
rect 19426 22924 19432 22976
rect 19484 22964 19490 22976
rect 19797 22967 19855 22973
rect 19797 22964 19809 22967
rect 19484 22936 19809 22964
rect 19484 22924 19490 22936
rect 19797 22933 19809 22936
rect 19843 22933 19855 22967
rect 19797 22927 19855 22933
rect 19889 22967 19947 22973
rect 19889 22933 19901 22967
rect 19935 22964 19947 22967
rect 20530 22964 20536 22976
rect 19935 22936 20536 22964
rect 19935 22933 19947 22936
rect 19889 22927 19947 22933
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 20806 22964 20812 22976
rect 20767 22936 20812 22964
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 21637 22967 21695 22973
rect 21637 22933 21649 22967
rect 21683 22964 21695 22967
rect 21818 22964 21824 22976
rect 21683 22936 21824 22964
rect 21683 22933 21695 22936
rect 21637 22927 21695 22933
rect 21818 22924 21824 22936
rect 21876 22924 21882 22976
rect 23290 22924 23296 22976
rect 23348 22964 23354 22976
rect 26068 22964 26096 23004
rect 23348 22936 26096 22964
rect 23348 22924 23354 22936
rect 26142 22924 26148 22976
rect 26200 22964 26206 22976
rect 26237 22967 26295 22973
rect 26237 22964 26249 22967
rect 26200 22936 26249 22964
rect 26200 22924 26206 22936
rect 26237 22933 26249 22936
rect 26283 22933 26295 22967
rect 26344 22964 26372 23004
rect 26970 22992 26976 23004
rect 27028 22992 27034 23044
rect 29564 22964 29592 23063
rect 29638 23060 29644 23072
rect 29696 23060 29702 23112
rect 29748 23032 29776 23267
rect 31754 23264 31760 23276
rect 31812 23264 31818 23316
rect 33686 23304 33692 23316
rect 33647 23276 33692 23304
rect 33686 23264 33692 23276
rect 33744 23264 33750 23316
rect 34790 23304 34796 23316
rect 34751 23276 34796 23304
rect 34790 23264 34796 23276
rect 34848 23264 34854 23316
rect 38102 23264 38108 23316
rect 38160 23304 38166 23316
rect 38654 23304 38660 23316
rect 38160 23276 38660 23304
rect 38160 23264 38166 23276
rect 38654 23264 38660 23276
rect 38712 23264 38718 23316
rect 42889 23307 42947 23313
rect 42889 23273 42901 23307
rect 42935 23304 42947 23307
rect 42978 23304 42984 23316
rect 42935 23276 42984 23304
rect 42935 23273 42947 23276
rect 42889 23267 42947 23273
rect 42978 23264 42984 23276
rect 43036 23264 43042 23316
rect 29914 23196 29920 23248
rect 29972 23236 29978 23248
rect 48133 23239 48191 23245
rect 48133 23236 48145 23239
rect 29972 23208 48145 23236
rect 29972 23196 29978 23208
rect 48133 23205 48145 23208
rect 48179 23205 48191 23239
rect 48133 23199 48191 23205
rect 30852 23140 33732 23168
rect 30852 23112 30880 23140
rect 30834 23100 30840 23112
rect 30795 23072 30840 23100
rect 30834 23060 30840 23072
rect 30892 23060 30898 23112
rect 33704 23109 33732 23140
rect 38378 23128 38384 23180
rect 38436 23168 38442 23180
rect 38841 23171 38899 23177
rect 38841 23168 38853 23171
rect 38436 23140 38853 23168
rect 38436 23128 38442 23140
rect 38841 23137 38853 23140
rect 38887 23137 38899 23171
rect 38841 23131 38899 23137
rect 39850 23128 39856 23180
rect 39908 23168 39914 23180
rect 39945 23171 40003 23177
rect 39945 23168 39957 23171
rect 39908 23140 39957 23168
rect 39908 23128 39914 23140
rect 39945 23137 39957 23140
rect 39991 23137 40003 23171
rect 39945 23131 40003 23137
rect 42334 23128 42340 23180
rect 42392 23168 42398 23180
rect 45465 23171 45523 23177
rect 42392 23140 42748 23168
rect 42392 23128 42398 23140
rect 31573 23103 31631 23109
rect 31573 23069 31585 23103
rect 31619 23069 31631 23103
rect 31573 23063 31631 23069
rect 33689 23103 33747 23109
rect 33689 23069 33701 23103
rect 33735 23100 33747 23103
rect 34701 23103 34759 23109
rect 34701 23100 34713 23103
rect 33735 23072 34713 23100
rect 33735 23069 33747 23072
rect 33689 23063 33747 23069
rect 34701 23069 34713 23072
rect 34747 23069 34759 23103
rect 34701 23063 34759 23069
rect 37001 23103 37059 23109
rect 37001 23069 37013 23103
rect 37047 23069 37059 23103
rect 38930 23100 38936 23112
rect 38891 23072 38936 23100
rect 37001 23063 37059 23069
rect 31588 23032 31616 23063
rect 32122 23032 32128 23044
rect 29748 23004 32128 23032
rect 32122 22992 32128 23004
rect 32180 22992 32186 23044
rect 33870 22992 33876 23044
rect 33928 23032 33934 23044
rect 37016 23032 37044 23063
rect 38930 23060 38936 23072
rect 38988 23060 38994 23112
rect 42720 23109 42748 23140
rect 45465 23137 45477 23171
rect 45511 23168 45523 23171
rect 45738 23168 45744 23180
rect 45511 23140 45744 23168
rect 45511 23137 45523 23140
rect 45465 23131 45523 23137
rect 45738 23128 45744 23140
rect 45796 23128 45802 23180
rect 46382 23168 46388 23180
rect 46343 23140 46388 23168
rect 46382 23128 46388 23140
rect 46440 23128 46446 23180
rect 42613 23103 42671 23109
rect 42613 23069 42625 23103
rect 42659 23069 42671 23103
rect 42613 23063 42671 23069
rect 42705 23103 42763 23109
rect 42705 23069 42717 23103
rect 42751 23100 42763 23103
rect 43349 23103 43407 23109
rect 43349 23100 43361 23103
rect 42751 23072 43361 23100
rect 42751 23069 42763 23072
rect 42705 23063 42763 23069
rect 43349 23069 43361 23072
rect 43395 23069 43407 23103
rect 43349 23063 43407 23069
rect 43533 23103 43591 23109
rect 43533 23069 43545 23103
rect 43579 23069 43591 23103
rect 43533 23063 43591 23069
rect 40126 23032 40132 23044
rect 33928 23004 39712 23032
rect 40087 23004 40132 23032
rect 33928 22992 33934 23004
rect 26344 22936 29592 22964
rect 26237 22927 26295 22933
rect 30926 22924 30932 22976
rect 30984 22964 30990 22976
rect 31021 22967 31079 22973
rect 31021 22964 31033 22967
rect 30984 22936 31033 22964
rect 30984 22924 30990 22936
rect 31021 22933 31033 22936
rect 31067 22933 31079 22967
rect 31021 22927 31079 22933
rect 37185 22967 37243 22973
rect 37185 22933 37197 22967
rect 37231 22964 37243 22967
rect 37274 22964 37280 22976
rect 37231 22936 37280 22964
rect 37231 22933 37243 22936
rect 37185 22927 37243 22933
rect 37274 22924 37280 22936
rect 37332 22924 37338 22976
rect 39301 22967 39359 22973
rect 39301 22933 39313 22967
rect 39347 22964 39359 22967
rect 39574 22964 39580 22976
rect 39347 22936 39580 22964
rect 39347 22933 39359 22936
rect 39301 22927 39359 22933
rect 39574 22924 39580 22936
rect 39632 22924 39638 22976
rect 39684 22964 39712 23004
rect 40126 22992 40132 23004
rect 40184 22992 40190 23044
rect 41782 23032 41788 23044
rect 41743 23004 41788 23032
rect 41782 22992 41788 23004
rect 41840 22992 41846 23044
rect 41874 22992 41880 23044
rect 41932 23032 41938 23044
rect 42628 23032 42656 23063
rect 43548 23032 43576 23063
rect 45002 23060 45008 23112
rect 45060 23100 45066 23112
rect 45281 23103 45339 23109
rect 45281 23100 45293 23103
rect 45060 23072 45293 23100
rect 45060 23060 45066 23072
rect 45281 23069 45293 23072
rect 45327 23069 45339 23103
rect 47302 23100 47308 23112
rect 45281 23063 45339 23069
rect 46676 23072 47308 23100
rect 46676 23032 46704 23072
rect 47302 23060 47308 23072
rect 47360 23060 47366 23112
rect 47946 23032 47952 23044
rect 41932 23004 46704 23032
rect 47907 23004 47952 23032
rect 41932 22992 41938 23004
rect 47946 22992 47952 23004
rect 48004 22992 48010 23044
rect 43254 22964 43260 22976
rect 39684 22936 43260 22964
rect 43254 22924 43260 22936
rect 43312 22924 43318 22976
rect 43438 22964 43444 22976
rect 43399 22936 43444 22964
rect 43438 22924 43444 22936
rect 43496 22924 43502 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 16022 22760 16028 22772
rect 15983 22732 16028 22760
rect 16022 22720 16028 22732
rect 16080 22760 16086 22772
rect 16206 22760 16212 22772
rect 16080 22732 16212 22760
rect 16080 22720 16086 22732
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 16761 22763 16819 22769
rect 16761 22729 16773 22763
rect 16807 22760 16819 22763
rect 16850 22760 16856 22772
rect 16807 22732 16856 22760
rect 16807 22729 16819 22732
rect 16761 22723 16819 22729
rect 16850 22720 16856 22732
rect 16908 22720 16914 22772
rect 17862 22720 17868 22772
rect 17920 22760 17926 22772
rect 19061 22763 19119 22769
rect 17920 22732 18920 22760
rect 17920 22720 17926 22732
rect 15470 22692 15476 22704
rect 15120 22664 15476 22692
rect 11698 22624 11704 22636
rect 11659 22596 11704 22624
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 13449 22627 13507 22633
rect 13449 22593 13461 22627
rect 13495 22624 13507 22627
rect 14642 22624 14648 22636
rect 13495 22596 14648 22624
rect 13495 22593 13507 22596
rect 13449 22587 13507 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 15120 22633 15148 22664
rect 15470 22652 15476 22664
rect 15528 22692 15534 22704
rect 17678 22692 17684 22704
rect 15528 22664 17684 22692
rect 15528 22652 15534 22664
rect 17678 22652 17684 22664
rect 17736 22652 17742 22704
rect 18322 22652 18328 22704
rect 18380 22652 18386 22704
rect 18892 22692 18920 22732
rect 19061 22729 19073 22763
rect 19107 22760 19119 22763
rect 19334 22760 19340 22772
rect 19107 22732 19340 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 19426 22720 19432 22772
rect 19484 22720 19490 22772
rect 19889 22763 19947 22769
rect 19889 22729 19901 22763
rect 19935 22760 19947 22763
rect 20070 22760 20076 22772
rect 19935 22732 20076 22760
rect 19935 22729 19947 22732
rect 19889 22723 19947 22729
rect 20070 22720 20076 22732
rect 20128 22760 20134 22772
rect 20901 22763 20959 22769
rect 20901 22760 20913 22763
rect 20128 22732 20913 22760
rect 20128 22720 20134 22732
rect 20901 22729 20913 22732
rect 20947 22729 20959 22763
rect 20901 22723 20959 22729
rect 23569 22763 23627 22769
rect 23569 22729 23581 22763
rect 23615 22760 23627 22763
rect 24762 22760 24768 22772
rect 23615 22732 24256 22760
rect 24723 22732 24768 22760
rect 23615 22729 23627 22732
rect 23569 22723 23627 22729
rect 19444 22692 19472 22720
rect 19521 22695 19579 22701
rect 19521 22692 19533 22695
rect 18892 22664 19533 22692
rect 19521 22661 19533 22664
rect 19567 22661 19579 22695
rect 19797 22695 19855 22701
rect 19797 22692 19809 22695
rect 19521 22655 19579 22661
rect 19628 22664 19809 22692
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22593 15163 22627
rect 15838 22624 15844 22636
rect 15799 22596 15844 22624
rect 15105 22587 15163 22593
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 16666 22624 16672 22636
rect 16627 22596 16672 22624
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 11793 22559 11851 22565
rect 11793 22525 11805 22559
rect 11839 22556 11851 22559
rect 11974 22556 11980 22568
rect 11839 22528 11980 22556
rect 11839 22525 11851 22528
rect 11793 22519 11851 22525
rect 11974 22516 11980 22528
rect 12032 22556 12038 22568
rect 12526 22556 12532 22568
rect 12032 22528 12532 22556
rect 12032 22516 12038 22528
rect 12526 22516 12532 22528
rect 12584 22516 12590 22568
rect 15194 22516 15200 22568
rect 15252 22516 15258 22568
rect 17310 22556 17316 22568
rect 17271 22528 17316 22556
rect 17310 22516 17316 22528
rect 17368 22516 17374 22568
rect 17589 22559 17647 22565
rect 17589 22525 17601 22559
rect 17635 22556 17647 22559
rect 18598 22556 18604 22568
rect 17635 22528 18604 22556
rect 17635 22525 17647 22528
rect 17589 22519 17647 22525
rect 18598 22516 18604 22528
rect 18656 22516 18662 22568
rect 19628 22556 19656 22664
rect 19797 22661 19809 22664
rect 19843 22692 19855 22695
rect 20530 22692 20536 22704
rect 19843 22664 20536 22692
rect 19843 22661 19855 22664
rect 19797 22655 19855 22661
rect 20530 22652 20536 22664
rect 20588 22652 20594 22704
rect 20806 22652 20812 22704
rect 20864 22692 20870 22704
rect 22097 22695 22155 22701
rect 22097 22692 22109 22695
rect 20864 22664 22109 22692
rect 20864 22652 20870 22664
rect 22097 22661 22109 22664
rect 22143 22661 22155 22695
rect 24121 22695 24179 22701
rect 24121 22692 24133 22695
rect 23322 22664 24133 22692
rect 22097 22655 22155 22661
rect 24121 22661 24133 22664
rect 24167 22661 24179 22695
rect 24121 22655 24179 22661
rect 24228 22692 24256 22732
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 25961 22763 26019 22769
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 26970 22760 26976 22772
rect 26007 22732 26976 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 26970 22720 26976 22732
rect 27028 22720 27034 22772
rect 27249 22763 27307 22769
rect 27249 22729 27261 22763
rect 27295 22760 27307 22763
rect 27338 22760 27344 22772
rect 27295 22732 27344 22760
rect 27295 22729 27307 22732
rect 27249 22723 27307 22729
rect 27338 22720 27344 22732
rect 27396 22720 27402 22772
rect 27798 22720 27804 22772
rect 27856 22760 27862 22772
rect 32858 22760 32864 22772
rect 27856 22732 32864 22760
rect 27856 22720 27862 22732
rect 32858 22720 32864 22732
rect 32916 22720 32922 22772
rect 39850 22720 39856 22772
rect 39908 22760 39914 22772
rect 40037 22763 40095 22769
rect 40037 22760 40049 22763
rect 39908 22732 40049 22760
rect 39908 22720 39914 22732
rect 40037 22729 40049 22732
rect 40083 22729 40095 22763
rect 40037 22723 40095 22729
rect 41782 22720 41788 22772
rect 41840 22760 41846 22772
rect 46382 22760 46388 22772
rect 41840 22732 46388 22760
rect 41840 22720 41846 22732
rect 46382 22720 46388 22732
rect 46440 22720 46446 22772
rect 48038 22760 48044 22772
rect 47999 22732 48044 22760
rect 48038 22720 48044 22732
rect 48096 22720 48102 22772
rect 26510 22692 26516 22704
rect 24228 22664 26516 22692
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22593 19763 22627
rect 20622 22624 20628 22636
rect 20583 22596 20628 22624
rect 19705 22587 19763 22593
rect 19260 22528 19656 22556
rect 15212 22488 15240 22516
rect 15212 22460 17448 22488
rect 11790 22380 11796 22432
rect 11848 22420 11854 22432
rect 12069 22423 12127 22429
rect 12069 22420 12081 22423
rect 11848 22392 12081 22420
rect 11848 22380 11854 22392
rect 12069 22389 12081 22392
rect 12115 22389 12127 22423
rect 12069 22383 12127 22389
rect 12342 22380 12348 22432
rect 12400 22420 12406 22432
rect 13633 22423 13691 22429
rect 13633 22420 13645 22423
rect 12400 22392 13645 22420
rect 12400 22380 12406 22392
rect 13633 22389 13645 22392
rect 13679 22420 13691 22423
rect 13722 22420 13728 22432
rect 13679 22392 13728 22420
rect 13679 22389 13691 22392
rect 13633 22383 13691 22389
rect 13722 22380 13728 22392
rect 13780 22380 13786 22432
rect 15194 22420 15200 22432
rect 15155 22392 15200 22420
rect 15194 22380 15200 22392
rect 15252 22380 15258 22432
rect 17420 22420 17448 22460
rect 19260 22420 19288 22528
rect 19720 22488 19748 22587
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 21818 22624 21824 22636
rect 20772 22596 20817 22624
rect 21779 22596 21824 22624
rect 20772 22584 20778 22596
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 23934 22584 23940 22636
rect 23992 22624 23998 22636
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 23992 22596 24041 22624
rect 23992 22584 23998 22596
rect 24029 22593 24041 22596
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 20162 22516 20168 22568
rect 20220 22556 20226 22568
rect 24228 22556 24256 22664
rect 26510 22652 26516 22664
rect 26568 22652 26574 22704
rect 38102 22692 38108 22704
rect 38063 22664 38108 22692
rect 38102 22652 38108 22664
rect 38160 22652 38166 22704
rect 45830 22692 45836 22704
rect 44744 22664 45836 22692
rect 24670 22624 24676 22636
rect 24631 22596 24676 22624
rect 24670 22584 24676 22596
rect 24728 22584 24734 22636
rect 25869 22627 25927 22633
rect 25869 22593 25881 22627
rect 25915 22593 25927 22627
rect 25869 22587 25927 22593
rect 20220 22528 24256 22556
rect 20220 22516 20226 22528
rect 19720 22460 20208 22488
rect 17420 22392 19288 22420
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19978 22420 19984 22432
rect 19392 22392 19984 22420
rect 19392 22380 19398 22392
rect 19978 22380 19984 22392
rect 20036 22420 20042 22432
rect 20073 22423 20131 22429
rect 20073 22420 20085 22423
rect 20036 22392 20085 22420
rect 20036 22380 20042 22392
rect 20073 22389 20085 22392
rect 20119 22389 20131 22423
rect 20180 22420 20208 22460
rect 25590 22448 25596 22500
rect 25648 22488 25654 22500
rect 25884 22488 25912 22587
rect 26142 22584 26148 22636
rect 26200 22624 26206 22636
rect 27065 22627 27123 22633
rect 27065 22624 27077 22627
rect 26200 22596 27077 22624
rect 26200 22584 26206 22596
rect 27065 22593 27077 22596
rect 27111 22624 27123 22627
rect 27801 22627 27859 22633
rect 27801 22624 27813 22627
rect 27111 22596 27813 22624
rect 27111 22593 27123 22596
rect 27065 22587 27123 22593
rect 27801 22593 27813 22596
rect 27847 22593 27859 22627
rect 27801 22587 27859 22593
rect 31113 22627 31171 22633
rect 31113 22593 31125 22627
rect 31159 22624 31171 22627
rect 31846 22624 31852 22636
rect 31159 22596 31852 22624
rect 31159 22593 31171 22596
rect 31113 22587 31171 22593
rect 31846 22584 31852 22596
rect 31904 22584 31910 22636
rect 32122 22624 32128 22636
rect 32083 22596 32128 22624
rect 32122 22584 32128 22596
rect 32180 22584 32186 22636
rect 33137 22627 33195 22633
rect 33137 22593 33149 22627
rect 33183 22624 33195 22627
rect 33870 22624 33876 22636
rect 33183 22596 33876 22624
rect 33183 22593 33195 22596
rect 33137 22587 33195 22593
rect 33870 22584 33876 22596
rect 33928 22584 33934 22636
rect 35161 22627 35219 22633
rect 35161 22593 35173 22627
rect 35207 22624 35219 22627
rect 35342 22624 35348 22636
rect 35207 22596 35348 22624
rect 35207 22593 35219 22596
rect 35161 22587 35219 22593
rect 35342 22584 35348 22596
rect 35400 22584 35406 22636
rect 37274 22624 37280 22636
rect 37235 22596 37280 22624
rect 37274 22584 37280 22596
rect 37332 22584 37338 22636
rect 39669 22627 39727 22633
rect 39669 22593 39681 22627
rect 39715 22593 39727 22627
rect 39669 22587 39727 22593
rect 31205 22559 31263 22565
rect 31205 22525 31217 22559
rect 31251 22556 31263 22559
rect 31478 22556 31484 22568
rect 31251 22528 31484 22556
rect 31251 22525 31263 22528
rect 31205 22519 31263 22525
rect 31478 22516 31484 22528
rect 31536 22516 31542 22568
rect 39574 22556 39580 22568
rect 39535 22528 39580 22556
rect 39574 22516 39580 22528
rect 39632 22516 39638 22568
rect 39684 22556 39712 22587
rect 40034 22584 40040 22636
rect 40092 22624 40098 22636
rect 40497 22627 40555 22633
rect 40497 22624 40509 22627
rect 40092 22596 40509 22624
rect 40092 22584 40098 22596
rect 40497 22593 40509 22596
rect 40543 22593 40555 22627
rect 40497 22587 40555 22593
rect 41693 22627 41751 22633
rect 41693 22593 41705 22627
rect 41739 22593 41751 22627
rect 41874 22624 41880 22636
rect 41835 22596 41880 22624
rect 41693 22587 41751 22593
rect 40218 22556 40224 22568
rect 39684 22528 40224 22556
rect 40218 22516 40224 22528
rect 40276 22516 40282 22568
rect 41708 22556 41736 22587
rect 41874 22584 41880 22596
rect 41932 22584 41938 22636
rect 42794 22584 42800 22636
rect 42852 22624 42858 22636
rect 44744 22633 44772 22664
rect 45830 22652 45836 22664
rect 45888 22652 45894 22704
rect 42981 22627 43039 22633
rect 42981 22624 42993 22627
rect 42852 22596 42993 22624
rect 42852 22584 42858 22596
rect 42981 22593 42993 22596
rect 43027 22593 43039 22627
rect 42981 22587 43039 22593
rect 44729 22627 44787 22633
rect 44729 22593 44741 22627
rect 44775 22593 44787 22627
rect 44729 22587 44787 22593
rect 47581 22627 47639 22633
rect 47581 22593 47593 22627
rect 47627 22593 47639 22627
rect 47581 22587 47639 22593
rect 42334 22556 42340 22568
rect 41708 22528 42340 22556
rect 42334 22516 42340 22528
rect 42392 22516 42398 22568
rect 42886 22556 42892 22568
rect 42847 22528 42892 22556
rect 42886 22516 42892 22528
rect 42944 22516 42950 22568
rect 43809 22559 43867 22565
rect 43809 22525 43821 22559
rect 43855 22556 43867 22559
rect 45186 22556 45192 22568
rect 43855 22528 45192 22556
rect 43855 22525 43867 22528
rect 43809 22519 43867 22525
rect 45186 22516 45192 22528
rect 45244 22516 45250 22568
rect 45373 22559 45431 22565
rect 45373 22525 45385 22559
rect 45419 22525 45431 22559
rect 46382 22556 46388 22568
rect 46343 22528 46388 22556
rect 45373 22519 45431 22525
rect 33870 22488 33876 22500
rect 25648 22460 33876 22488
rect 25648 22448 25654 22460
rect 33870 22448 33876 22460
rect 33928 22488 33934 22500
rect 35894 22488 35900 22500
rect 33928 22460 35900 22488
rect 33928 22448 33934 22460
rect 35894 22448 35900 22460
rect 35952 22448 35958 22500
rect 44545 22491 44603 22497
rect 44545 22457 44557 22491
rect 44591 22488 44603 22491
rect 45388 22488 45416 22519
rect 46382 22516 46388 22528
rect 46440 22516 46446 22568
rect 44591 22460 45416 22488
rect 44591 22457 44603 22460
rect 44545 22451 44603 22457
rect 45922 22448 45928 22500
rect 45980 22488 45986 22500
rect 47596 22488 47624 22587
rect 45980 22460 47624 22488
rect 45980 22448 45986 22460
rect 20346 22420 20352 22432
rect 20180 22392 20352 22420
rect 20073 22383 20131 22389
rect 20346 22380 20352 22392
rect 20404 22420 20410 22432
rect 22186 22420 22192 22432
rect 20404 22392 22192 22420
rect 20404 22380 20410 22392
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 27890 22380 27896 22432
rect 27948 22420 27954 22432
rect 27985 22423 28043 22429
rect 27985 22420 27997 22423
rect 27948 22392 27997 22420
rect 27948 22380 27954 22392
rect 27985 22389 27997 22392
rect 28031 22389 28043 22423
rect 27985 22383 28043 22389
rect 31202 22380 31208 22432
rect 31260 22420 31266 22432
rect 31481 22423 31539 22429
rect 31481 22420 31493 22423
rect 31260 22392 31493 22420
rect 31260 22380 31266 22392
rect 31481 22389 31493 22392
rect 31527 22389 31539 22423
rect 32214 22420 32220 22432
rect 32175 22392 32220 22420
rect 31481 22383 31539 22389
rect 32214 22380 32220 22392
rect 32272 22380 32278 22432
rect 32950 22380 32956 22432
rect 33008 22420 33014 22432
rect 33321 22423 33379 22429
rect 33321 22420 33333 22423
rect 33008 22392 33333 22420
rect 33008 22380 33014 22392
rect 33321 22389 33333 22392
rect 33367 22389 33379 22423
rect 33321 22383 33379 22389
rect 33686 22380 33692 22432
rect 33744 22420 33750 22432
rect 34057 22423 34115 22429
rect 34057 22420 34069 22423
rect 33744 22392 34069 22420
rect 33744 22380 33750 22392
rect 34057 22389 34069 22392
rect 34103 22389 34115 22423
rect 34057 22383 34115 22389
rect 34790 22380 34796 22432
rect 34848 22420 34854 22432
rect 34977 22423 35035 22429
rect 34977 22420 34989 22423
rect 34848 22392 34989 22420
rect 34848 22380 34854 22392
rect 34977 22389 34989 22392
rect 35023 22389 35035 22423
rect 40586 22420 40592 22432
rect 40547 22392 40592 22420
rect 34977 22383 35035 22389
rect 40586 22380 40592 22392
rect 40644 22380 40650 22432
rect 40862 22380 40868 22432
rect 40920 22420 40926 22432
rect 40957 22423 41015 22429
rect 40957 22420 40969 22423
rect 40920 22392 40969 22420
rect 40920 22380 40926 22392
rect 40957 22389 40969 22392
rect 41003 22389 41015 22423
rect 41782 22420 41788 22432
rect 41743 22392 41788 22420
rect 40957 22383 41015 22389
rect 41782 22380 41788 22392
rect 41840 22380 41846 22432
rect 45094 22380 45100 22432
rect 45152 22420 45158 22432
rect 45646 22420 45652 22432
rect 45152 22392 45652 22420
rect 45152 22380 45158 22392
rect 45646 22380 45652 22392
rect 45704 22380 45710 22432
rect 47210 22380 47216 22432
rect 47268 22420 47274 22432
rect 47673 22423 47731 22429
rect 47673 22420 47685 22423
rect 47268 22392 47685 22420
rect 47268 22380 47274 22392
rect 47673 22389 47685 22392
rect 47719 22389 47731 22423
rect 47673 22383 47731 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 11790 22225 11796 22228
rect 11780 22219 11796 22225
rect 11780 22185 11792 22219
rect 11780 22179 11796 22185
rect 11790 22176 11796 22179
rect 11848 22176 11854 22228
rect 17310 22176 17316 22228
rect 17368 22216 17374 22228
rect 17405 22219 17463 22225
rect 17405 22216 17417 22219
rect 17368 22188 17417 22216
rect 17368 22176 17374 22188
rect 17405 22185 17417 22188
rect 17451 22185 17463 22219
rect 26142 22216 26148 22228
rect 17405 22179 17463 22185
rect 17512 22188 26148 22216
rect 14642 22108 14648 22160
rect 14700 22148 14706 22160
rect 15838 22148 15844 22160
rect 14700 22120 15844 22148
rect 14700 22108 14706 22120
rect 15838 22108 15844 22120
rect 15896 22148 15902 22160
rect 17512 22148 17540 22188
rect 26142 22176 26148 22188
rect 26200 22176 26206 22228
rect 31202 22225 31208 22228
rect 31192 22219 31208 22225
rect 31192 22185 31204 22219
rect 31192 22179 31208 22185
rect 31202 22176 31208 22179
rect 31260 22176 31266 22228
rect 34977 22219 35035 22225
rect 34977 22216 34989 22219
rect 34900 22188 34989 22216
rect 15896 22120 17540 22148
rect 15896 22108 15902 22120
rect 18598 22108 18604 22160
rect 18656 22148 18662 22160
rect 25958 22148 25964 22160
rect 18656 22120 19656 22148
rect 18656 22108 18662 22120
rect 11790 22040 11796 22092
rect 11848 22080 11854 22092
rect 13541 22083 13599 22089
rect 13541 22080 13553 22083
rect 11848 22052 13553 22080
rect 11848 22040 11854 22052
rect 13541 22049 13553 22052
rect 13587 22049 13599 22083
rect 13541 22043 13599 22049
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22080 15071 22083
rect 15194 22080 15200 22092
rect 15059 22052 15200 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 19334 22080 19340 22092
rect 15344 22052 15389 22080
rect 19295 22052 19340 22080
rect 15344 22040 15350 22052
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19628 22080 19656 22120
rect 25608 22120 25964 22148
rect 19797 22083 19855 22089
rect 19797 22080 19809 22083
rect 19628 22052 19809 22080
rect 19797 22049 19809 22052
rect 19843 22049 19855 22083
rect 19797 22043 19855 22049
rect 22186 22040 22192 22092
rect 22244 22080 22250 22092
rect 25608 22080 25636 22120
rect 25958 22108 25964 22120
rect 26016 22108 26022 22160
rect 34900 22094 34928 22188
rect 34977 22185 34989 22188
rect 35023 22216 35035 22219
rect 35161 22219 35219 22225
rect 35023 22188 35112 22216
rect 35023 22185 35035 22188
rect 34977 22179 35035 22185
rect 35084 22148 35112 22188
rect 35161 22185 35173 22219
rect 35207 22216 35219 22219
rect 35342 22216 35348 22228
rect 35207 22188 35348 22216
rect 35207 22185 35219 22188
rect 35161 22179 35219 22185
rect 35342 22176 35348 22188
rect 35400 22176 35406 22228
rect 35529 22219 35587 22225
rect 35529 22185 35541 22219
rect 35575 22216 35587 22219
rect 35618 22216 35624 22228
rect 35575 22188 35624 22216
rect 35575 22185 35587 22188
rect 35529 22179 35587 22185
rect 35544 22148 35572 22179
rect 35618 22176 35624 22188
rect 35676 22176 35682 22228
rect 40126 22176 40132 22228
rect 40184 22216 40190 22228
rect 40681 22219 40739 22225
rect 40681 22216 40693 22219
rect 40184 22188 40693 22216
rect 40184 22176 40190 22188
rect 40681 22185 40693 22188
rect 40727 22185 40739 22219
rect 40681 22179 40739 22185
rect 45186 22176 45192 22228
rect 45244 22216 45250 22228
rect 45462 22216 45468 22228
rect 45244 22188 45468 22216
rect 45244 22176 45250 22188
rect 45462 22176 45468 22188
rect 45520 22176 45526 22228
rect 45646 22216 45652 22228
rect 45607 22188 45652 22216
rect 45646 22176 45652 22188
rect 45704 22176 45710 22228
rect 45830 22216 45836 22228
rect 45791 22188 45836 22216
rect 45830 22176 45836 22188
rect 45888 22176 45894 22228
rect 35084 22120 35572 22148
rect 42337 22151 42395 22157
rect 42337 22117 42349 22151
rect 42383 22117 42395 22151
rect 45922 22148 45928 22160
rect 42337 22111 42395 22117
rect 45388 22120 45928 22148
rect 22244 22052 25636 22080
rect 22244 22040 22250 22052
rect 28902 22040 28908 22092
rect 28960 22080 28966 22092
rect 30926 22080 30932 22092
rect 28960 22052 29592 22080
rect 30887 22052 30932 22080
rect 28960 22040 28966 22052
rect 11514 22012 11520 22024
rect 11475 21984 11520 22012
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 14829 22015 14887 22021
rect 14829 21981 14841 22015
rect 14875 21981 14887 22015
rect 14829 21975 14887 21981
rect 13078 21944 13084 21956
rect 13018 21916 13084 21944
rect 13078 21904 13084 21916
rect 13136 21904 13142 21956
rect 14844 21944 14872 21975
rect 16206 21972 16212 22024
rect 16264 22012 16270 22024
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 16264 21984 17233 22012
rect 16264 21972 16270 21984
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 19426 22012 19432 22024
rect 19387 21984 19432 22012
rect 17221 21975 17279 21981
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 22012 24639 22015
rect 24854 22012 24860 22024
rect 24627 21984 24860 22012
rect 24627 21981 24639 21984
rect 24581 21975 24639 21981
rect 24854 21972 24860 21984
rect 24912 21972 24918 22024
rect 25222 22012 25228 22024
rect 25183 21984 25228 22012
rect 25222 21972 25228 21984
rect 25280 21972 25286 22024
rect 25682 21972 25688 22024
rect 25740 22012 25746 22024
rect 27249 22015 27307 22021
rect 27249 22012 27261 22015
rect 25740 21984 27261 22012
rect 25740 21972 25746 21984
rect 27249 21981 27261 21984
rect 27295 21981 27307 22015
rect 27430 22012 27436 22024
rect 27391 21984 27436 22012
rect 27249 21975 27307 21981
rect 27430 21972 27436 21984
rect 27488 21972 27494 22024
rect 27890 21972 27896 22024
rect 27948 22012 27954 22024
rect 28077 22015 28135 22021
rect 28077 22012 28089 22015
rect 27948 21984 28089 22012
rect 27948 21972 27954 21984
rect 28077 21981 28089 21984
rect 28123 21981 28135 22015
rect 28994 22012 29000 22024
rect 28955 21984 29000 22012
rect 28077 21975 28135 21981
rect 28994 21972 29000 21984
rect 29052 21972 29058 22024
rect 29564 22021 29592 22052
rect 30926 22040 30932 22052
rect 30984 22040 30990 22092
rect 31754 22040 31760 22092
rect 31812 22080 31818 22092
rect 32677 22083 32735 22089
rect 32677 22080 32689 22083
rect 31812 22052 32689 22080
rect 31812 22040 31818 22052
rect 32677 22049 32689 22052
rect 32723 22080 32735 22083
rect 33042 22080 33048 22092
rect 32723 22052 33048 22080
rect 32723 22049 32735 22052
rect 32677 22043 32735 22049
rect 33042 22040 33048 22052
rect 33100 22040 33106 22092
rect 34333 22083 34391 22089
rect 34333 22049 34345 22083
rect 34379 22080 34391 22083
rect 34900 22080 35020 22094
rect 34379 22052 35020 22080
rect 34379 22049 34391 22052
rect 34333 22043 34391 22049
rect 40218 22040 40224 22092
rect 40276 22080 40282 22092
rect 42352 22080 42380 22111
rect 45388 22080 45416 22120
rect 45922 22108 45928 22120
rect 45980 22108 45986 22160
rect 40276 22052 42380 22080
rect 44284 22052 45416 22080
rect 40276 22040 40282 22052
rect 29549 22015 29607 22021
rect 29549 21981 29561 22015
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 32490 21972 32496 22024
rect 32548 22012 32554 22024
rect 32950 22012 32956 22024
rect 32548 21984 32956 22012
rect 32548 21972 32554 21984
rect 32950 21972 32956 21984
rect 33008 21972 33014 22024
rect 34698 22012 34704 22024
rect 34659 21984 34704 22012
rect 34698 21972 34704 21984
rect 34756 21972 34762 22024
rect 37093 22015 37151 22021
rect 37093 22012 37105 22015
rect 34808 21984 37105 22012
rect 16574 21944 16580 21956
rect 14844 21916 16580 21944
rect 16574 21904 16580 21916
rect 16632 21904 16638 21956
rect 24670 21904 24676 21956
rect 24728 21944 24734 21956
rect 27908 21944 27936 21972
rect 24728 21916 27936 21944
rect 24728 21904 24734 21916
rect 32214 21904 32220 21956
rect 32272 21904 32278 21956
rect 33778 21944 33784 21956
rect 32600 21916 32812 21944
rect 33739 21916 33784 21944
rect 24394 21876 24400 21888
rect 24355 21848 24400 21876
rect 24394 21836 24400 21848
rect 24452 21836 24458 21888
rect 25314 21876 25320 21888
rect 25275 21848 25320 21876
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 27433 21879 27491 21885
rect 27433 21845 27445 21879
rect 27479 21876 27491 21879
rect 27706 21876 27712 21888
rect 27479 21848 27712 21876
rect 27479 21845 27491 21848
rect 27433 21839 27491 21845
rect 27706 21836 27712 21848
rect 27764 21836 27770 21888
rect 28261 21879 28319 21885
rect 28261 21845 28273 21879
rect 28307 21876 28319 21879
rect 28442 21876 28448 21888
rect 28307 21848 28448 21876
rect 28307 21845 28319 21848
rect 28261 21839 28319 21845
rect 28442 21836 28448 21848
rect 28500 21836 28506 21888
rect 28810 21876 28816 21888
rect 28771 21848 28816 21876
rect 28810 21836 28816 21848
rect 28868 21836 28874 21888
rect 29641 21879 29699 21885
rect 29641 21845 29653 21879
rect 29687 21876 29699 21879
rect 29730 21876 29736 21888
rect 29687 21848 29736 21876
rect 29687 21845 29699 21848
rect 29641 21839 29699 21845
rect 29730 21836 29736 21848
rect 29788 21836 29794 21888
rect 30190 21836 30196 21888
rect 30248 21876 30254 21888
rect 32600 21876 32628 21916
rect 30248 21848 32628 21876
rect 32784 21876 32812 21916
rect 33778 21904 33784 21916
rect 33836 21904 33842 21956
rect 34808 21876 34836 21984
rect 37093 21981 37105 21984
rect 37139 21981 37151 22015
rect 37093 21975 37151 21981
rect 39945 22015 40003 22021
rect 39945 21981 39957 22015
rect 39991 22012 40003 22015
rect 40034 22012 40040 22024
rect 39991 21984 40040 22012
rect 39991 21981 40003 21984
rect 39945 21975 40003 21981
rect 40034 21972 40040 21984
rect 40092 21972 40098 22024
rect 40129 22015 40187 22021
rect 40129 21981 40141 22015
rect 40175 22012 40187 22015
rect 40586 22012 40592 22024
rect 40175 21984 40592 22012
rect 40175 21981 40187 21984
rect 40129 21975 40187 21981
rect 40586 21972 40592 21984
rect 40644 21972 40650 22024
rect 40862 22012 40868 22024
rect 40823 21984 40868 22012
rect 40862 21972 40868 21984
rect 40920 21972 40926 22024
rect 41782 21972 41788 22024
rect 41840 22012 41846 22024
rect 42521 22015 42579 22021
rect 42521 22012 42533 22015
rect 41840 21984 42533 22012
rect 41840 21972 41846 21984
rect 42521 21981 42533 21984
rect 42567 21981 42579 22015
rect 42521 21975 42579 21981
rect 42613 22015 42671 22021
rect 42613 21981 42625 22015
rect 42659 22012 42671 22015
rect 42794 22012 42800 22024
rect 42659 21984 42800 22012
rect 42659 21981 42671 21984
rect 42613 21975 42671 21981
rect 42794 21972 42800 21984
rect 42852 21972 42858 22024
rect 44284 22021 44312 22052
rect 45462 22040 45468 22092
rect 45520 22080 45526 22092
rect 46293 22083 46351 22089
rect 46293 22080 46305 22083
rect 45520 22052 46305 22080
rect 45520 22040 45526 22052
rect 46293 22049 46305 22052
rect 46339 22049 46351 22083
rect 46474 22080 46480 22092
rect 46435 22052 46480 22080
rect 46293 22043 46351 22049
rect 46474 22040 46480 22052
rect 46532 22040 46538 22092
rect 46750 22080 46756 22092
rect 46711 22052 46756 22080
rect 46750 22040 46756 22052
rect 46808 22040 46814 22092
rect 44269 22015 44327 22021
rect 44269 21981 44281 22015
rect 44315 21981 44327 22015
rect 44450 22012 44456 22024
rect 44411 21984 44456 22012
rect 44269 21975 44327 21981
rect 44450 21972 44456 21984
rect 44508 21972 44514 22024
rect 45281 22015 45339 22021
rect 45281 21981 45293 22015
rect 45327 21981 45339 22015
rect 45554 22012 45560 22024
rect 45515 21984 45560 22012
rect 45281 21975 45339 21981
rect 36265 21947 36323 21953
rect 36265 21913 36277 21947
rect 36311 21944 36323 21947
rect 36311 21916 36584 21944
rect 36311 21913 36323 21916
rect 36265 21907 36323 21913
rect 36354 21876 36360 21888
rect 32784 21848 34836 21876
rect 36315 21848 36360 21876
rect 30248 21836 30254 21848
rect 36354 21836 36360 21848
rect 36412 21836 36418 21888
rect 36556 21876 36584 21916
rect 36630 21904 36636 21956
rect 36688 21944 36694 21956
rect 37277 21947 37335 21953
rect 37277 21944 37289 21947
rect 36688 21916 37289 21944
rect 36688 21904 36694 21916
rect 37277 21913 37289 21916
rect 37323 21913 37335 21947
rect 37277 21907 37335 21913
rect 38933 21947 38991 21953
rect 38933 21913 38945 21947
rect 38979 21913 38991 21947
rect 40218 21944 40224 21956
rect 40179 21916 40224 21944
rect 38933 21907 38991 21913
rect 37182 21876 37188 21888
rect 36556 21848 37188 21876
rect 37182 21836 37188 21848
rect 37240 21836 37246 21888
rect 38948 21876 38976 21907
rect 40218 21904 40224 21916
rect 40276 21904 40282 21956
rect 42337 21947 42395 21953
rect 42337 21913 42349 21947
rect 42383 21944 42395 21947
rect 43438 21944 43444 21956
rect 42383 21916 43444 21944
rect 42383 21913 42395 21916
rect 42337 21907 42395 21913
rect 43438 21904 43444 21916
rect 43496 21904 43502 21956
rect 45094 21944 45100 21956
rect 43548 21916 45100 21944
rect 43548 21876 43576 21916
rect 45094 21904 45100 21916
rect 45152 21904 45158 21956
rect 45296 21944 45324 21975
rect 45554 21972 45560 21984
rect 45612 21972 45618 22024
rect 46014 21944 46020 21956
rect 45296 21916 46020 21944
rect 46014 21904 46020 21916
rect 46072 21904 46078 21956
rect 38948 21848 43576 21876
rect 44453 21879 44511 21885
rect 44453 21845 44465 21879
rect 44499 21876 44511 21879
rect 45646 21876 45652 21888
rect 44499 21848 45652 21876
rect 44499 21845 44511 21848
rect 44453 21839 44511 21845
rect 45646 21836 45652 21848
rect 45704 21876 45710 21888
rect 46290 21876 46296 21888
rect 45704 21848 46296 21876
rect 45704 21836 45710 21848
rect 46290 21836 46296 21848
rect 46348 21836 46354 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 11514 21632 11520 21684
rect 11572 21672 11578 21684
rect 11977 21675 12035 21681
rect 11977 21672 11989 21675
rect 11572 21644 11989 21672
rect 11572 21632 11578 21644
rect 11977 21641 11989 21644
rect 12023 21641 12035 21675
rect 13078 21672 13084 21684
rect 13039 21644 13084 21672
rect 11977 21635 12035 21641
rect 13078 21632 13084 21644
rect 13136 21632 13142 21684
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22373 21675 22431 21681
rect 22373 21672 22385 21675
rect 22244 21644 22385 21672
rect 22244 21632 22250 21644
rect 22373 21641 22385 21644
rect 22419 21641 22431 21675
rect 24670 21672 24676 21684
rect 22373 21635 22431 21641
rect 23400 21644 24676 21672
rect 3602 21564 3608 21616
rect 3660 21604 3666 21616
rect 14461 21607 14519 21613
rect 3660 21576 14228 21604
rect 3660 21564 3666 21576
rect 11790 21536 11796 21548
rect 11751 21508 11796 21536
rect 11790 21496 11796 21508
rect 11848 21536 11854 21548
rect 12342 21536 12348 21548
rect 11848 21508 12348 21536
rect 11848 21496 11854 21508
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21536 13047 21539
rect 13814 21536 13820 21548
rect 13035 21508 13820 21536
rect 13035 21505 13047 21508
rect 12989 21499 13047 21505
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14 21360 20 21412
rect 72 21400 78 21412
rect 11422 21400 11428 21412
rect 72 21372 11428 21400
rect 72 21360 78 21372
rect 11422 21360 11428 21372
rect 11480 21360 11486 21412
rect 14200 21400 14228 21576
rect 14461 21573 14473 21607
rect 14507 21604 14519 21607
rect 15378 21604 15384 21616
rect 14507 21576 15384 21604
rect 14507 21573 14519 21576
rect 14461 21567 14519 21573
rect 15378 21564 15384 21576
rect 15436 21564 15442 21616
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21536 17003 21539
rect 17773 21539 17831 21545
rect 17773 21536 17785 21539
rect 16991 21508 17785 21536
rect 16991 21505 17003 21508
rect 16945 21499 17003 21505
rect 17773 21505 17785 21508
rect 17819 21536 17831 21539
rect 18506 21536 18512 21548
rect 17819 21508 18512 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18506 21496 18512 21508
rect 18564 21496 18570 21548
rect 18874 21536 18880 21548
rect 18835 21508 18880 21536
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 22278 21536 22284 21548
rect 22239 21508 22284 21536
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 23400 21545 23428 21644
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 25130 21632 25136 21684
rect 25188 21672 25194 21684
rect 25590 21672 25596 21684
rect 25188 21644 25596 21672
rect 25188 21632 25194 21644
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 36630 21672 36636 21684
rect 25700 21644 36492 21672
rect 36591 21644 36636 21672
rect 24305 21607 24363 21613
rect 24305 21573 24317 21607
rect 24351 21604 24363 21607
rect 24394 21604 24400 21616
rect 24351 21576 24400 21604
rect 24351 21573 24363 21576
rect 24305 21567 24363 21573
rect 24394 21564 24400 21576
rect 24452 21564 24458 21616
rect 25314 21564 25320 21616
rect 25372 21564 25378 21616
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21468 14335 21471
rect 14458 21468 14464 21480
rect 14323 21440 14464 21468
rect 14323 21437 14335 21440
rect 14277 21431 14335 21437
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 14737 21471 14795 21477
rect 14737 21437 14749 21471
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23615 21440 24041 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 14752 21400 14780 21431
rect 24302 21428 24308 21480
rect 24360 21468 24366 21480
rect 25700 21468 25728 21644
rect 28721 21607 28779 21613
rect 28721 21573 28733 21607
rect 28767 21604 28779 21607
rect 28810 21604 28816 21616
rect 28767 21576 28816 21604
rect 28767 21573 28779 21576
rect 28721 21567 28779 21573
rect 28810 21564 28816 21576
rect 28868 21564 28874 21616
rect 29730 21564 29736 21616
rect 29788 21564 29794 21616
rect 33689 21607 33747 21613
rect 33689 21573 33701 21607
rect 33735 21604 33747 21607
rect 35897 21607 35955 21613
rect 35897 21604 35909 21607
rect 33735 21576 35909 21604
rect 33735 21573 33747 21576
rect 33689 21567 33747 21573
rect 35897 21573 35909 21576
rect 35943 21573 35955 21607
rect 35897 21567 35955 21573
rect 26878 21496 26884 21548
rect 26936 21536 26942 21548
rect 27246 21536 27252 21548
rect 26936 21508 27252 21536
rect 26936 21496 26942 21508
rect 27246 21496 27252 21508
rect 27304 21536 27310 21548
rect 27525 21539 27583 21545
rect 27525 21536 27537 21539
rect 27304 21508 27537 21536
rect 27304 21496 27310 21508
rect 27525 21505 27537 21508
rect 27571 21505 27583 21539
rect 28442 21536 28448 21548
rect 28403 21508 28448 21536
rect 27525 21499 27583 21505
rect 28442 21496 28448 21508
rect 28500 21496 28506 21548
rect 32490 21536 32496 21548
rect 32451 21508 32496 21536
rect 32490 21496 32496 21508
rect 32548 21496 32554 21548
rect 35342 21536 35348 21548
rect 35303 21508 35348 21536
rect 35342 21496 35348 21508
rect 35400 21496 35406 21548
rect 35805 21539 35863 21545
rect 35805 21505 35817 21539
rect 35851 21505 35863 21539
rect 35805 21499 35863 21505
rect 24360 21440 25728 21468
rect 24360 21428 24366 21440
rect 27154 21428 27160 21480
rect 27212 21468 27218 21480
rect 30190 21468 30196 21480
rect 27212 21440 30196 21468
rect 27212 21428 27218 21440
rect 30190 21428 30196 21440
rect 30248 21428 30254 21480
rect 32766 21468 32772 21480
rect 32727 21440 32772 21468
rect 32766 21428 32772 21440
rect 32824 21428 32830 21480
rect 33505 21471 33563 21477
rect 33505 21437 33517 21471
rect 33551 21437 33563 21471
rect 33505 21431 33563 21437
rect 14200 21372 14780 21400
rect 20898 21360 20904 21412
rect 20956 21400 20962 21412
rect 20956 21372 24164 21400
rect 20956 21360 20962 21372
rect 15746 21292 15752 21344
rect 15804 21332 15810 21344
rect 16666 21332 16672 21344
rect 15804 21304 16672 21332
rect 15804 21292 15810 21304
rect 16666 21292 16672 21304
rect 16724 21332 16730 21344
rect 17129 21335 17187 21341
rect 17129 21332 17141 21335
rect 16724 21304 17141 21332
rect 16724 21292 16730 21304
rect 17129 21301 17141 21304
rect 17175 21301 17187 21335
rect 17954 21332 17960 21344
rect 17915 21304 17960 21332
rect 17129 21295 17187 21301
rect 17954 21292 17960 21304
rect 18012 21292 18018 21344
rect 18966 21332 18972 21344
rect 18927 21304 18972 21332
rect 18966 21292 18972 21304
rect 19024 21292 19030 21344
rect 24136 21332 24164 21372
rect 30282 21360 30288 21412
rect 30340 21400 30346 21412
rect 33520 21400 33548 21431
rect 30340 21372 33548 21400
rect 35820 21400 35848 21499
rect 36464 21468 36492 21644
rect 36630 21632 36636 21644
rect 36688 21632 36694 21684
rect 40034 21632 40040 21684
rect 40092 21672 40098 21684
rect 45741 21675 45799 21681
rect 45741 21672 45753 21675
rect 40092 21644 45753 21672
rect 40092 21632 40098 21644
rect 45741 21641 45753 21644
rect 45787 21641 45799 21675
rect 45741 21635 45799 21641
rect 46014 21632 46020 21684
rect 46072 21672 46078 21684
rect 46072 21644 46612 21672
rect 46072 21632 46078 21644
rect 37274 21564 37280 21616
rect 37332 21604 37338 21616
rect 37645 21607 37703 21613
rect 37645 21604 37657 21607
rect 37332 21576 37657 21604
rect 37332 21564 37338 21576
rect 37645 21573 37657 21576
rect 37691 21573 37703 21607
rect 37645 21567 37703 21573
rect 38930 21564 38936 21616
rect 38988 21604 38994 21616
rect 43530 21604 43536 21616
rect 38988 21576 43536 21604
rect 38988 21564 38994 21576
rect 43530 21564 43536 21576
rect 43588 21564 43594 21616
rect 45462 21604 45468 21616
rect 45423 21576 45468 21604
rect 45462 21564 45468 21576
rect 45520 21564 45526 21616
rect 45557 21607 45615 21613
rect 45557 21573 45569 21607
rect 45603 21573 45615 21607
rect 45557 21567 45615 21573
rect 36541 21539 36599 21545
rect 36541 21505 36553 21539
rect 36587 21536 36599 21539
rect 37292 21536 37320 21564
rect 42702 21536 42708 21548
rect 36587 21508 37320 21536
rect 42663 21508 42708 21536
rect 36587 21505 36599 21508
rect 36541 21499 36599 21505
rect 42702 21496 42708 21508
rect 42760 21496 42766 21548
rect 42889 21539 42947 21545
rect 42889 21505 42901 21539
rect 42935 21505 42947 21539
rect 43806 21536 43812 21548
rect 43767 21508 43812 21536
rect 42889 21499 42947 21505
rect 36464 21440 41414 21468
rect 38194 21400 38200 21412
rect 35820 21372 38200 21400
rect 30340 21360 30346 21372
rect 25682 21332 25688 21344
rect 24136 21304 25688 21332
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 25777 21335 25835 21341
rect 25777 21301 25789 21335
rect 25823 21332 25835 21335
rect 25958 21332 25964 21344
rect 25823 21304 25964 21332
rect 25823 21301 25835 21304
rect 25777 21295 25835 21301
rect 25958 21292 25964 21304
rect 26016 21292 26022 21344
rect 27709 21335 27767 21341
rect 27709 21301 27721 21335
rect 27755 21332 27767 21335
rect 27890 21332 27896 21344
rect 27755 21304 27896 21332
rect 27755 21301 27767 21304
rect 27709 21295 27767 21301
rect 27890 21292 27896 21304
rect 27948 21292 27954 21344
rect 32766 21292 32772 21344
rect 32824 21332 32830 21344
rect 35820 21332 35848 21372
rect 38194 21360 38200 21372
rect 38252 21360 38258 21412
rect 41386 21400 41414 21440
rect 42610 21428 42616 21480
rect 42668 21468 42674 21480
rect 42904 21468 42932 21499
rect 43806 21496 43812 21508
rect 43864 21496 43870 21548
rect 43990 21536 43996 21548
rect 43951 21508 43996 21536
rect 43990 21496 43996 21508
rect 44048 21496 44054 21548
rect 45373 21539 45431 21545
rect 45373 21505 45385 21539
rect 45419 21505 45431 21539
rect 45572 21536 45600 21567
rect 45830 21536 45836 21548
rect 45572 21508 45836 21536
rect 45373 21499 45431 21505
rect 42668 21440 42932 21468
rect 45388 21468 45416 21499
rect 45830 21496 45836 21508
rect 45888 21496 45894 21548
rect 46032 21468 46060 21632
rect 46584 21616 46612 21644
rect 46566 21564 46572 21616
rect 46624 21604 46630 21616
rect 47765 21607 47823 21613
rect 47765 21604 47777 21607
rect 46624 21576 47777 21604
rect 46624 21564 46630 21576
rect 47765 21573 47777 21576
rect 47811 21573 47823 21607
rect 47765 21567 47823 21573
rect 46198 21536 46204 21548
rect 46159 21508 46204 21536
rect 46198 21496 46204 21508
rect 46256 21496 46262 21548
rect 46290 21496 46296 21548
rect 46348 21536 46354 21548
rect 47581 21539 47639 21545
rect 47581 21536 47593 21539
rect 46348 21508 47593 21536
rect 46348 21496 46354 21508
rect 47581 21505 47593 21508
rect 47627 21505 47639 21539
rect 47581 21499 47639 21505
rect 45388 21440 46060 21468
rect 42668 21428 42674 21440
rect 46106 21428 46112 21480
rect 46164 21468 46170 21480
rect 46477 21471 46535 21477
rect 46477 21468 46489 21471
rect 46164 21440 46489 21468
rect 46164 21428 46170 21440
rect 46477 21437 46489 21440
rect 46523 21437 46535 21471
rect 46477 21431 46535 21437
rect 44358 21400 44364 21412
rect 41386 21372 44364 21400
rect 44358 21360 44364 21372
rect 44416 21360 44422 21412
rect 44450 21360 44456 21412
rect 44508 21400 44514 21412
rect 45189 21403 45247 21409
rect 45189 21400 45201 21403
rect 44508 21372 45201 21400
rect 44508 21360 44514 21372
rect 45189 21369 45201 21372
rect 45235 21369 45247 21403
rect 45189 21363 45247 21369
rect 38930 21332 38936 21344
rect 32824 21304 35848 21332
rect 38891 21304 38936 21332
rect 32824 21292 32830 21304
rect 38930 21292 38936 21304
rect 38988 21292 38994 21344
rect 42705 21335 42763 21341
rect 42705 21301 42717 21335
rect 42751 21332 42763 21335
rect 43162 21332 43168 21344
rect 42751 21304 43168 21332
rect 42751 21301 42763 21304
rect 42705 21295 42763 21301
rect 43162 21292 43168 21304
rect 43220 21292 43226 21344
rect 43901 21335 43959 21341
rect 43901 21301 43913 21335
rect 43947 21332 43959 21335
rect 44266 21332 44272 21344
rect 43947 21304 44272 21332
rect 43947 21301 43959 21304
rect 43901 21295 43959 21301
rect 44266 21292 44272 21304
rect 44324 21292 44330 21344
rect 44726 21332 44732 21344
rect 44687 21304 44732 21332
rect 44726 21292 44732 21304
rect 44784 21292 44790 21344
rect 45204 21332 45232 21363
rect 45278 21360 45284 21412
rect 45336 21400 45342 21412
rect 47949 21403 48007 21409
rect 47949 21400 47961 21403
rect 45336 21372 47961 21400
rect 45336 21360 45342 21372
rect 47949 21369 47961 21372
rect 47995 21369 48007 21403
rect 47949 21363 48007 21369
rect 47210 21332 47216 21344
rect 45204 21304 47216 21332
rect 47210 21292 47216 21304
rect 47268 21292 47274 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 42705 21131 42763 21137
rect 2280 21100 33824 21128
rect 2280 21088 2286 21100
rect 24765 21063 24823 21069
rect 24765 21029 24777 21063
rect 24811 21060 24823 21063
rect 25409 21063 25467 21069
rect 25409 21060 25421 21063
rect 24811 21032 25421 21060
rect 24811 21029 24823 21032
rect 24765 21023 24823 21029
rect 25409 21029 25421 21032
rect 25455 21029 25467 21063
rect 25409 21023 25467 21029
rect 25682 21020 25688 21072
rect 25740 21060 25746 21072
rect 33410 21060 33416 21072
rect 25740 21032 33416 21060
rect 25740 21020 25746 21032
rect 33410 21020 33416 21032
rect 33468 21020 33474 21072
rect 3694 20952 3700 21004
rect 3752 20992 3758 21004
rect 11333 20995 11391 21001
rect 11333 20992 11345 20995
rect 3752 20964 11345 20992
rect 3752 20952 3758 20964
rect 11333 20961 11345 20964
rect 11379 20961 11391 20995
rect 11333 20955 11391 20961
rect 11422 20952 11428 21004
rect 11480 20992 11486 21004
rect 16853 20995 16911 21001
rect 16853 20992 16865 20995
rect 11480 20964 16865 20992
rect 11480 20952 11486 20964
rect 16853 20961 16865 20964
rect 16899 20961 16911 20995
rect 22830 20992 22836 21004
rect 22743 20964 22836 20992
rect 16853 20955 16911 20961
rect 22830 20952 22836 20964
rect 22888 20992 22894 21004
rect 24302 20992 24308 21004
rect 22888 20964 24308 20992
rect 22888 20952 22894 20964
rect 24302 20952 24308 20964
rect 24360 20952 24366 21004
rect 24854 20992 24860 21004
rect 24815 20964 24860 20992
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 25590 20992 25596 21004
rect 25551 20964 25596 20992
rect 25590 20952 25596 20964
rect 25648 20952 25654 21004
rect 25869 20995 25927 21001
rect 25869 20961 25881 20995
rect 25915 20992 25927 20995
rect 25958 20992 25964 21004
rect 25915 20964 25964 20992
rect 25915 20961 25927 20964
rect 25869 20955 25927 20961
rect 25958 20952 25964 20964
rect 26016 20952 26022 21004
rect 27706 20992 27712 21004
rect 27667 20964 27712 20992
rect 27706 20952 27712 20964
rect 27764 20952 27770 21004
rect 30282 20992 30288 21004
rect 27816 20964 30288 20992
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20893 10931 20927
rect 10873 20887 10931 20893
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20924 13231 20927
rect 13814 20924 13820 20936
rect 13219 20896 13820 20924
rect 13219 20893 13231 20896
rect 13173 20887 13231 20893
rect 10888 20788 10916 20887
rect 13814 20884 13820 20896
rect 13872 20924 13878 20936
rect 14366 20924 14372 20936
rect 13872 20896 14372 20924
rect 13872 20884 13878 20896
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14642 20924 14648 20936
rect 14603 20896 14648 20924
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 15746 20924 15752 20936
rect 15707 20896 15752 20924
rect 15746 20884 15752 20896
rect 15804 20884 15810 20936
rect 16390 20924 16396 20936
rect 16351 20896 16396 20924
rect 16390 20884 16396 20896
rect 16448 20884 16454 20936
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 19337 20927 19395 20933
rect 19337 20924 19349 20927
rect 18012 20896 19349 20924
rect 18012 20884 18018 20896
rect 19337 20893 19349 20896
rect 19383 20893 19395 20927
rect 19337 20887 19395 20893
rect 20346 20884 20352 20936
rect 20404 20884 20410 20936
rect 20717 20927 20775 20933
rect 20717 20893 20729 20927
rect 20763 20924 20775 20927
rect 22281 20927 22339 20933
rect 22281 20924 22293 20927
rect 20763 20896 22293 20924
rect 20763 20893 20775 20896
rect 20717 20887 20775 20893
rect 22281 20893 22293 20896
rect 22327 20924 22339 20927
rect 22554 20924 22560 20936
rect 22327 20896 22560 20924
rect 22327 20893 22339 20896
rect 22281 20887 22339 20893
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 25498 20884 25504 20936
rect 25556 20924 25562 20936
rect 25685 20927 25743 20933
rect 25685 20924 25697 20927
rect 25556 20896 25697 20924
rect 25556 20884 25562 20896
rect 25685 20893 25697 20896
rect 25731 20893 25743 20927
rect 25685 20887 25743 20893
rect 25777 20927 25835 20933
rect 25777 20893 25789 20927
rect 25823 20924 25835 20927
rect 25823 20896 25968 20924
rect 25823 20893 25835 20896
rect 25777 20887 25835 20893
rect 11054 20856 11060 20868
rect 11015 20828 11060 20856
rect 11054 20816 11060 20828
rect 11112 20816 11118 20868
rect 15841 20859 15899 20865
rect 15841 20825 15853 20859
rect 15887 20856 15899 20859
rect 16577 20859 16635 20865
rect 16577 20856 16589 20859
rect 15887 20828 16589 20856
rect 15887 20825 15899 20828
rect 15841 20819 15899 20825
rect 16577 20825 16589 20828
rect 16623 20825 16635 20859
rect 20364 20856 20392 20884
rect 21266 20856 21272 20868
rect 20364 20828 21272 20856
rect 16577 20819 16635 20825
rect 21266 20816 21272 20828
rect 21324 20816 21330 20868
rect 24397 20859 24455 20865
rect 24397 20825 24409 20859
rect 24443 20856 24455 20859
rect 25314 20856 25320 20868
rect 24443 20828 25320 20856
rect 24443 20825 24455 20828
rect 24397 20819 24455 20825
rect 25314 20816 25320 20828
rect 25372 20816 25378 20868
rect 25940 20856 25968 20896
rect 26050 20884 26056 20936
rect 26108 20924 26114 20936
rect 26789 20927 26847 20933
rect 26789 20924 26801 20927
rect 26108 20896 26801 20924
rect 26108 20884 26114 20896
rect 26789 20893 26801 20896
rect 26835 20893 26847 20927
rect 26789 20887 26847 20893
rect 26970 20884 26976 20936
rect 27028 20924 27034 20936
rect 27430 20924 27436 20936
rect 27028 20896 27436 20924
rect 27028 20884 27034 20896
rect 27430 20884 27436 20896
rect 27488 20884 27494 20936
rect 27816 20933 27844 20964
rect 30282 20952 30288 20964
rect 30340 20952 30346 21004
rect 31205 20995 31263 21001
rect 31205 20961 31217 20995
rect 31251 20992 31263 20995
rect 31754 20992 31760 21004
rect 31251 20964 31760 20992
rect 31251 20961 31263 20964
rect 31205 20955 31263 20961
rect 31754 20952 31760 20964
rect 31812 20952 31818 21004
rect 27801 20927 27859 20933
rect 27801 20893 27813 20927
rect 27847 20893 27859 20927
rect 27801 20887 27859 20893
rect 26142 20856 26148 20868
rect 25940 20828 26148 20856
rect 11882 20788 11888 20800
rect 10888 20760 11888 20788
rect 11882 20748 11888 20760
rect 11940 20748 11946 20800
rect 13262 20788 13268 20800
rect 13223 20760 13268 20788
rect 13262 20748 13268 20760
rect 13320 20748 13326 20800
rect 14921 20791 14979 20797
rect 14921 20757 14933 20791
rect 14967 20788 14979 20791
rect 16666 20788 16672 20800
rect 14967 20760 16672 20788
rect 14967 20757 14979 20760
rect 14921 20751 14979 20757
rect 16666 20748 16672 20760
rect 16724 20788 16730 20800
rect 17494 20788 17500 20800
rect 16724 20760 17500 20788
rect 16724 20748 16730 20760
rect 17494 20748 17500 20760
rect 17552 20748 17558 20800
rect 19429 20791 19487 20797
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 20346 20788 20352 20800
rect 19475 20760 20352 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 25774 20748 25780 20800
rect 25832 20788 25838 20800
rect 25940 20788 25968 20828
rect 26142 20816 26148 20828
rect 26200 20856 26206 20868
rect 27816 20856 27844 20887
rect 27890 20884 27896 20936
rect 27948 20924 27954 20936
rect 28629 20927 28687 20933
rect 28629 20924 28641 20927
rect 27948 20896 28641 20924
rect 27948 20884 27954 20896
rect 28629 20893 28641 20896
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28902 20884 28908 20936
rect 28960 20924 28966 20936
rect 29641 20927 29699 20933
rect 29641 20924 29653 20927
rect 28960 20896 29653 20924
rect 28960 20884 28966 20896
rect 29641 20893 29653 20896
rect 29687 20893 29699 20927
rect 33686 20924 33692 20936
rect 33647 20896 33692 20924
rect 29641 20887 29699 20893
rect 33686 20884 33692 20896
rect 33744 20884 33750 20936
rect 33796 20924 33824 21100
rect 42705 21097 42717 21131
rect 42751 21128 42763 21131
rect 42794 21128 42800 21140
rect 42751 21100 42800 21128
rect 42751 21097 42763 21100
rect 42705 21091 42763 21097
rect 42794 21088 42800 21100
rect 42852 21088 42858 21140
rect 44358 21088 44364 21140
rect 44416 21128 44422 21140
rect 47578 21128 47584 21140
rect 44416 21100 47584 21128
rect 44416 21088 44422 21100
rect 47578 21088 47584 21100
rect 47636 21088 47642 21140
rect 35434 21060 35440 21072
rect 33980 21032 35440 21060
rect 33980 21001 34008 21032
rect 35434 21020 35440 21032
rect 35492 21060 35498 21072
rect 47486 21060 47492 21072
rect 35492 21032 47492 21060
rect 35492 21020 35498 21032
rect 47486 21020 47492 21032
rect 47544 21020 47550 21072
rect 33965 20995 34023 21001
rect 33965 20961 33977 20995
rect 34011 20961 34023 20995
rect 38930 20992 38936 21004
rect 33965 20955 34023 20961
rect 34072 20964 38936 20992
rect 34072 20924 34100 20964
rect 38930 20952 38936 20964
rect 38988 20952 38994 21004
rect 42260 20964 43116 20992
rect 42260 20936 42288 20964
rect 37274 20924 37280 20936
rect 33796 20896 34100 20924
rect 37235 20896 37280 20924
rect 37274 20884 37280 20896
rect 37332 20884 37338 20936
rect 38010 20924 38016 20936
rect 37971 20896 38016 20924
rect 38010 20884 38016 20896
rect 38068 20884 38074 20936
rect 42061 20927 42119 20933
rect 42061 20893 42073 20927
rect 42107 20893 42119 20927
rect 42242 20924 42248 20936
rect 42203 20896 42248 20924
rect 42061 20887 42119 20893
rect 26200 20828 27844 20856
rect 26200 20816 26206 20828
rect 28718 20816 28724 20868
rect 28776 20856 28782 20868
rect 31386 20856 31392 20868
rect 28776 20828 29960 20856
rect 31347 20828 31392 20856
rect 28776 20816 28782 20828
rect 25832 20760 25968 20788
rect 27157 20791 27215 20797
rect 25832 20748 25838 20760
rect 27157 20757 27169 20791
rect 27203 20788 27215 20791
rect 27890 20788 27896 20800
rect 27203 20760 27896 20788
rect 27203 20757 27215 20760
rect 27157 20751 27215 20757
rect 27890 20748 27896 20760
rect 27948 20748 27954 20800
rect 28166 20788 28172 20800
rect 28127 20760 28172 20788
rect 28166 20748 28172 20760
rect 28224 20748 28230 20800
rect 28534 20748 28540 20800
rect 28592 20788 28598 20800
rect 28813 20791 28871 20797
rect 28813 20788 28825 20791
rect 28592 20760 28825 20788
rect 28592 20748 28598 20760
rect 28813 20757 28825 20760
rect 28859 20757 28871 20791
rect 28813 20751 28871 20757
rect 29733 20791 29791 20797
rect 29733 20757 29745 20791
rect 29779 20788 29791 20791
rect 29822 20788 29828 20800
rect 29779 20760 29828 20788
rect 29779 20757 29791 20760
rect 29733 20751 29791 20757
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 29932 20788 29960 20828
rect 31386 20816 31392 20828
rect 31444 20816 31450 20868
rect 33042 20856 33048 20868
rect 33003 20828 33048 20856
rect 33042 20816 33048 20828
rect 33100 20816 33106 20868
rect 34978 20859 35036 20865
rect 34978 20825 34990 20859
rect 35024 20825 35036 20859
rect 34978 20819 35036 20825
rect 34992 20788 35020 20819
rect 35066 20816 35072 20868
rect 35124 20856 35130 20868
rect 35986 20856 35992 20868
rect 35124 20828 35169 20856
rect 35947 20828 35992 20856
rect 35124 20816 35130 20828
rect 35986 20816 35992 20828
rect 36044 20816 36050 20868
rect 29932 20760 35020 20788
rect 42076 20788 42104 20887
rect 42242 20884 42248 20896
rect 42300 20884 42306 20936
rect 42886 20924 42892 20936
rect 42847 20896 42892 20924
rect 42886 20884 42892 20896
rect 42944 20884 42950 20936
rect 43088 20933 43116 20964
rect 44726 20952 44732 21004
rect 44784 20992 44790 21004
rect 46293 20995 46351 21001
rect 46293 20992 46305 20995
rect 44784 20964 46305 20992
rect 44784 20952 44790 20964
rect 46293 20961 46305 20964
rect 46339 20961 46351 20995
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 46293 20955 46351 20961
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 42981 20927 43039 20933
rect 42981 20893 42993 20927
rect 43027 20893 43039 20927
rect 42981 20887 43039 20893
rect 43073 20927 43131 20933
rect 43073 20893 43085 20927
rect 43119 20893 43131 20927
rect 43073 20887 43131 20893
rect 42153 20859 42211 20865
rect 42153 20825 42165 20859
rect 42199 20856 42211 20859
rect 42996 20856 43024 20887
rect 43162 20884 43168 20936
rect 43220 20924 43226 20936
rect 43714 20924 43720 20936
rect 43220 20896 43265 20924
rect 43675 20896 43720 20924
rect 43220 20884 43226 20896
rect 43714 20884 43720 20896
rect 43772 20884 43778 20936
rect 43898 20924 43904 20936
rect 43859 20896 43904 20924
rect 43898 20884 43904 20896
rect 43956 20884 43962 20936
rect 45189 20927 45247 20933
rect 45189 20893 45201 20927
rect 45235 20924 45247 20927
rect 45278 20924 45284 20936
rect 45235 20896 45284 20924
rect 45235 20893 45247 20896
rect 45189 20887 45247 20893
rect 45278 20884 45284 20896
rect 45336 20884 45342 20936
rect 45649 20927 45707 20933
rect 45649 20893 45661 20927
rect 45695 20893 45707 20927
rect 45649 20887 45707 20893
rect 42199 20828 42932 20856
rect 42996 20828 43208 20856
rect 42199 20825 42211 20828
rect 42153 20819 42211 20825
rect 42904 20800 42932 20828
rect 43180 20800 43208 20828
rect 43530 20816 43536 20868
rect 43588 20856 43594 20868
rect 45664 20856 45692 20887
rect 43588 20828 45692 20856
rect 45741 20859 45799 20865
rect 43588 20816 43594 20828
rect 45741 20825 45753 20859
rect 45787 20856 45799 20859
rect 46477 20859 46535 20865
rect 46477 20856 46489 20859
rect 45787 20828 46489 20856
rect 45787 20825 45799 20828
rect 45741 20819 45799 20825
rect 46477 20825 46489 20828
rect 46523 20825 46535 20859
rect 46477 20819 46535 20825
rect 42794 20788 42800 20800
rect 42076 20760 42800 20788
rect 42794 20748 42800 20760
rect 42852 20748 42858 20800
rect 42886 20748 42892 20800
rect 42944 20748 42950 20800
rect 43162 20748 43168 20800
rect 43220 20788 43226 20800
rect 43806 20788 43812 20800
rect 43220 20760 43812 20788
rect 43220 20748 43226 20760
rect 43806 20748 43812 20760
rect 43864 20748 43870 20800
rect 45005 20791 45063 20797
rect 45005 20757 45017 20791
rect 45051 20788 45063 20791
rect 45370 20788 45376 20800
rect 45051 20760 45376 20788
rect 45051 20757 45063 20760
rect 45005 20751 45063 20757
rect 45370 20748 45376 20760
rect 45428 20748 45434 20800
rect 45554 20748 45560 20800
rect 45612 20788 45618 20800
rect 46014 20788 46020 20800
rect 45612 20760 46020 20788
rect 45612 20748 45618 20760
rect 46014 20748 46020 20760
rect 46072 20748 46078 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 10873 20587 10931 20593
rect 10873 20553 10885 20587
rect 10919 20584 10931 20587
rect 11054 20584 11060 20596
rect 10919 20556 11060 20584
rect 10919 20553 10931 20556
rect 10873 20547 10931 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 11164 20556 19104 20584
rect 3970 20476 3976 20528
rect 4028 20516 4034 20528
rect 11164 20516 11192 20556
rect 13262 20516 13268 20528
rect 4028 20488 11192 20516
rect 13018 20488 13268 20516
rect 4028 20476 4034 20488
rect 13262 20476 13268 20488
rect 13320 20476 13326 20528
rect 15378 20516 15384 20528
rect 15339 20488 15384 20516
rect 15378 20476 15384 20488
rect 15436 20476 15442 20528
rect 18966 20516 18972 20528
rect 18927 20488 18972 20516
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 19076 20516 19104 20556
rect 19150 20544 19156 20596
rect 19208 20584 19214 20596
rect 22646 20584 22652 20596
rect 19208 20556 22652 20584
rect 19208 20544 19214 20556
rect 22646 20544 22652 20556
rect 22704 20584 22710 20596
rect 23385 20587 23443 20593
rect 23385 20584 23397 20587
rect 22704 20556 23397 20584
rect 22704 20544 22710 20556
rect 23385 20553 23397 20556
rect 23431 20553 23443 20587
rect 23385 20547 23443 20553
rect 25590 20544 25596 20596
rect 25648 20584 25654 20596
rect 25961 20587 26019 20593
rect 25961 20584 25973 20587
rect 25648 20556 25973 20584
rect 25648 20544 25654 20556
rect 25961 20553 25973 20556
rect 26007 20584 26019 20587
rect 26050 20584 26056 20596
rect 26007 20556 26056 20584
rect 26007 20553 26019 20556
rect 25961 20547 26019 20553
rect 26050 20544 26056 20556
rect 26108 20544 26114 20596
rect 26970 20584 26976 20596
rect 26931 20556 26976 20584
rect 26970 20544 26976 20556
rect 27028 20544 27034 20596
rect 28077 20587 28135 20593
rect 28077 20553 28089 20587
rect 28123 20584 28135 20587
rect 28994 20584 29000 20596
rect 28123 20556 29000 20584
rect 28123 20553 28135 20556
rect 28077 20547 28135 20553
rect 28994 20544 29000 20556
rect 29052 20544 29058 20596
rect 30282 20584 30288 20596
rect 30243 20556 30288 20584
rect 30282 20544 30288 20556
rect 30340 20544 30346 20596
rect 31386 20584 31392 20596
rect 31347 20556 31392 20584
rect 31386 20544 31392 20556
rect 31444 20544 31450 20596
rect 41877 20587 41935 20593
rect 41877 20553 41889 20587
rect 41923 20584 41935 20587
rect 42242 20584 42248 20596
rect 41923 20556 42248 20584
rect 41923 20553 41935 20556
rect 41877 20547 41935 20553
rect 42242 20544 42248 20556
rect 42300 20544 42306 20596
rect 42978 20544 42984 20596
rect 43036 20584 43042 20596
rect 44269 20587 44327 20593
rect 44269 20584 44281 20587
rect 43036 20556 44281 20584
rect 43036 20544 43042 20556
rect 44269 20553 44281 20556
rect 44315 20553 44327 20587
rect 44269 20547 44327 20553
rect 46474 20544 46480 20596
rect 46532 20584 46538 20596
rect 47673 20587 47731 20593
rect 47673 20584 47685 20587
rect 46532 20556 47685 20584
rect 46532 20544 46538 20556
rect 47673 20553 47685 20556
rect 47719 20553 47731 20587
rect 47673 20547 47731 20553
rect 25774 20516 25780 20528
rect 19076 20488 25084 20516
rect 25735 20488 25780 20516
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 11422 20448 11428 20460
rect 10827 20420 11428 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 11422 20408 11428 20420
rect 11480 20408 11486 20460
rect 13722 20448 13728 20460
rect 13683 20420 13728 20448
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 15746 20448 15752 20460
rect 15335 20420 15752 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 15746 20408 15752 20420
rect 15804 20448 15810 20460
rect 16206 20448 16212 20460
rect 15804 20420 16212 20448
rect 15804 20408 15810 20420
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 16761 20451 16819 20457
rect 16761 20417 16773 20451
rect 16807 20448 16819 20451
rect 17402 20448 17408 20460
rect 16807 20420 17408 20448
rect 16807 20417 16819 20420
rect 16761 20411 16819 20417
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 17494 20408 17500 20460
rect 17552 20448 17558 20460
rect 17552 20420 17597 20448
rect 17552 20408 17558 20420
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 22244 20420 22293 20448
rect 22244 20408 22250 20420
rect 22281 20417 22293 20420
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 23201 20451 23259 20457
rect 23201 20417 23213 20451
rect 23247 20448 23259 20451
rect 23290 20448 23296 20460
rect 23247 20420 23296 20448
rect 23247 20417 23259 20420
rect 23201 20411 23259 20417
rect 23290 20408 23296 20420
rect 23348 20408 23354 20460
rect 23937 20451 23995 20457
rect 23937 20417 23949 20451
rect 23983 20448 23995 20451
rect 24670 20448 24676 20460
rect 23983 20420 24676 20448
rect 23983 20417 23995 20420
rect 23937 20411 23995 20417
rect 24670 20408 24676 20420
rect 24728 20408 24734 20460
rect 25056 20448 25084 20488
rect 25774 20476 25780 20488
rect 25832 20476 25838 20528
rect 25866 20476 25872 20528
rect 25924 20516 25930 20528
rect 26510 20516 26516 20528
rect 25924 20488 26516 20516
rect 25924 20476 25930 20488
rect 26510 20476 26516 20488
rect 26568 20516 26574 20528
rect 26988 20516 27016 20544
rect 27982 20516 27988 20528
rect 26568 20488 27016 20516
rect 27080 20488 27988 20516
rect 26568 20476 26574 20488
rect 27080 20448 27108 20488
rect 27982 20476 27988 20488
rect 28040 20476 28046 20528
rect 28166 20476 28172 20528
rect 28224 20516 28230 20528
rect 28813 20519 28871 20525
rect 28813 20516 28825 20519
rect 28224 20488 28825 20516
rect 28224 20476 28230 20488
rect 28813 20485 28825 20488
rect 28859 20485 28871 20519
rect 28813 20479 28871 20485
rect 29822 20476 29828 20528
rect 29880 20476 29886 20528
rect 33870 20516 33876 20528
rect 33831 20488 33876 20516
rect 33870 20476 33876 20488
rect 33928 20476 33934 20528
rect 34698 20476 34704 20528
rect 34756 20516 34762 20528
rect 35529 20519 35587 20525
rect 35529 20516 35541 20519
rect 34756 20488 35541 20516
rect 34756 20476 34762 20488
rect 35529 20485 35541 20488
rect 35575 20516 35587 20519
rect 35618 20516 35624 20528
rect 35575 20488 35624 20516
rect 35575 20485 35587 20488
rect 35529 20479 35587 20485
rect 35618 20476 35624 20488
rect 35676 20476 35682 20528
rect 35986 20476 35992 20528
rect 36044 20516 36050 20528
rect 36449 20519 36507 20525
rect 36449 20516 36461 20519
rect 36044 20488 36461 20516
rect 36044 20476 36050 20488
rect 36449 20485 36461 20488
rect 36495 20485 36507 20519
rect 43714 20516 43720 20528
rect 36449 20479 36507 20485
rect 41386 20488 43720 20516
rect 25056 20420 27108 20448
rect 27154 20408 27160 20460
rect 27212 20448 27218 20460
rect 27706 20448 27712 20460
rect 27212 20420 27257 20448
rect 27667 20420 27712 20448
rect 27212 20408 27218 20420
rect 27706 20408 27712 20420
rect 27764 20408 27770 20460
rect 27890 20448 27896 20460
rect 27851 20420 27896 20448
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 28534 20448 28540 20460
rect 28495 20420 28540 20448
rect 28534 20408 28540 20420
rect 28592 20408 28598 20460
rect 31294 20448 31300 20460
rect 31255 20420 31300 20448
rect 31294 20408 31300 20420
rect 31352 20408 31358 20460
rect 33505 20451 33563 20457
rect 33505 20448 33517 20451
rect 31726 20420 33517 20448
rect 11514 20380 11520 20392
rect 11475 20352 11520 20380
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 11793 20383 11851 20389
rect 11793 20349 11805 20383
rect 11839 20380 11851 20383
rect 12342 20380 12348 20392
rect 11839 20352 12348 20380
rect 11839 20349 11851 20352
rect 11793 20343 11851 20349
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 18785 20383 18843 20389
rect 18785 20349 18797 20383
rect 18831 20380 18843 20383
rect 19426 20380 19432 20392
rect 18831 20352 19432 20380
rect 18831 20349 18843 20352
rect 18785 20343 18843 20349
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20349 19579 20383
rect 22462 20380 22468 20392
rect 22423 20352 22468 20380
rect 19521 20343 19579 20349
rect 13265 20315 13323 20321
rect 13265 20281 13277 20315
rect 13311 20312 13323 20315
rect 19334 20312 19340 20324
rect 13311 20284 19340 20312
rect 13311 20281 13323 20284
rect 13265 20275 13323 20281
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 13280 20244 13308 20275
rect 19334 20272 19340 20284
rect 19392 20272 19398 20324
rect 13722 20244 13728 20256
rect 11940 20216 13308 20244
rect 13683 20216 13728 20244
rect 11940 20204 11946 20216
rect 13722 20204 13728 20216
rect 13780 20204 13786 20256
rect 16942 20244 16948 20256
rect 16903 20216 16948 20244
rect 16942 20204 16948 20216
rect 17000 20204 17006 20256
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 17497 20247 17555 20253
rect 17497 20244 17509 20247
rect 17276 20216 17509 20244
rect 17276 20204 17282 20216
rect 17497 20213 17509 20216
rect 17543 20213 17555 20247
rect 17497 20207 17555 20213
rect 18414 20204 18420 20256
rect 18472 20244 18478 20256
rect 19536 20244 19564 20343
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 22554 20340 22560 20392
rect 22612 20380 22618 20392
rect 31726 20380 31754 20420
rect 33505 20417 33517 20420
rect 33551 20448 33563 20451
rect 33686 20448 33692 20460
rect 33551 20420 33692 20448
rect 33551 20417 33563 20420
rect 33505 20411 33563 20417
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 36464 20448 36492 20479
rect 41386 20448 41414 20488
rect 43714 20476 43720 20488
rect 43772 20476 43778 20528
rect 43898 20476 43904 20528
rect 43956 20516 43962 20528
rect 45370 20516 45376 20528
rect 43956 20488 44588 20516
rect 45331 20488 45376 20516
rect 43956 20476 43962 20488
rect 36464 20420 41414 20448
rect 41693 20451 41751 20457
rect 41693 20417 41705 20451
rect 41739 20417 41751 20451
rect 41693 20411 41751 20417
rect 41877 20451 41935 20457
rect 41877 20417 41889 20451
rect 41923 20448 41935 20451
rect 42610 20448 42616 20460
rect 41923 20420 42616 20448
rect 41923 20417 41935 20420
rect 41877 20411 41935 20417
rect 35434 20380 35440 20392
rect 22612 20352 31754 20380
rect 35395 20352 35440 20380
rect 22612 20340 22618 20352
rect 35434 20340 35440 20352
rect 35492 20340 35498 20392
rect 41708 20380 41736 20411
rect 42610 20408 42616 20420
rect 42668 20408 42674 20460
rect 42981 20451 43039 20457
rect 42981 20417 42993 20451
rect 43027 20448 43039 20451
rect 43070 20448 43076 20460
rect 43027 20420 43076 20448
rect 43027 20417 43039 20420
rect 42981 20411 43039 20417
rect 43070 20408 43076 20420
rect 43128 20408 43134 20460
rect 43732 20448 43760 20476
rect 44560 20457 44588 20488
rect 45370 20476 45376 20488
rect 45428 20476 45434 20528
rect 44361 20451 44419 20457
rect 44361 20448 44373 20451
rect 43732 20420 44373 20448
rect 44361 20417 44373 20420
rect 44407 20417 44419 20451
rect 44361 20411 44419 20417
rect 44545 20451 44603 20457
rect 44545 20417 44557 20451
rect 44591 20417 44603 20451
rect 44545 20411 44603 20417
rect 46566 20408 46572 20460
rect 46624 20448 46630 20460
rect 47581 20451 47639 20457
rect 47581 20448 47593 20451
rect 46624 20420 47593 20448
rect 46624 20408 46630 20420
rect 47581 20417 47593 20420
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 42702 20380 42708 20392
rect 41708 20352 42708 20380
rect 42702 20340 42708 20352
rect 42760 20340 42766 20392
rect 42886 20380 42892 20392
rect 42847 20352 42892 20380
rect 42886 20340 42892 20352
rect 42944 20340 42950 20392
rect 43530 20380 43536 20392
rect 43491 20352 43536 20380
rect 43530 20340 43536 20352
rect 43588 20380 43594 20392
rect 45189 20383 45247 20389
rect 45189 20380 45201 20383
rect 43588 20352 45201 20380
rect 43588 20340 43594 20352
rect 45189 20349 45201 20352
rect 45235 20349 45247 20383
rect 46382 20380 46388 20392
rect 46343 20352 46388 20380
rect 45189 20343 45247 20349
rect 46382 20340 46388 20352
rect 46440 20340 46446 20392
rect 22480 20312 22508 20340
rect 25038 20312 25044 20324
rect 22480 20284 25044 20312
rect 25038 20272 25044 20284
rect 25096 20272 25102 20324
rect 25590 20312 25596 20324
rect 25551 20284 25596 20312
rect 25590 20272 25596 20284
rect 25648 20272 25654 20324
rect 25774 20272 25780 20324
rect 25832 20312 25838 20324
rect 27154 20312 27160 20324
rect 25832 20284 27160 20312
rect 25832 20272 25838 20284
rect 27154 20272 27160 20284
rect 27212 20272 27218 20324
rect 32214 20272 32220 20324
rect 32272 20312 32278 20324
rect 42518 20312 42524 20324
rect 32272 20284 42524 20312
rect 32272 20272 32278 20284
rect 42518 20272 42524 20284
rect 42576 20272 42582 20324
rect 44085 20315 44143 20321
rect 44085 20281 44097 20315
rect 44131 20312 44143 20315
rect 44131 20284 44220 20312
rect 44131 20281 44143 20284
rect 44085 20275 44143 20281
rect 44192 20256 44220 20284
rect 18472 20216 19564 20244
rect 18472 20204 18478 20216
rect 23750 20204 23756 20256
rect 23808 20244 23814 20256
rect 24029 20247 24087 20253
rect 24029 20244 24041 20247
rect 23808 20216 24041 20244
rect 23808 20204 23814 20216
rect 24029 20213 24041 20216
rect 24075 20213 24087 20247
rect 24029 20207 24087 20213
rect 25314 20204 25320 20256
rect 25372 20244 25378 20256
rect 26145 20247 26203 20253
rect 26145 20244 26157 20247
rect 25372 20216 26157 20244
rect 25372 20204 25378 20216
rect 26145 20213 26157 20216
rect 26191 20213 26203 20247
rect 26145 20207 26203 20213
rect 26326 20204 26332 20256
rect 26384 20244 26390 20256
rect 31294 20244 31300 20256
rect 26384 20216 31300 20244
rect 26384 20204 26390 20216
rect 31294 20204 31300 20216
rect 31352 20244 31358 20256
rect 37458 20244 37464 20256
rect 31352 20216 37464 20244
rect 31352 20204 31358 20216
rect 37458 20204 37464 20216
rect 37516 20244 37522 20256
rect 42886 20244 42892 20256
rect 37516 20216 42892 20244
rect 37516 20204 37522 20216
rect 42886 20204 42892 20216
rect 42944 20204 42950 20256
rect 44174 20204 44180 20256
rect 44232 20204 44238 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 11609 20043 11667 20049
rect 11609 20040 11621 20043
rect 11572 20012 11621 20040
rect 11572 20000 11578 20012
rect 11609 20009 11621 20012
rect 11655 20009 11667 20043
rect 12342 20040 12348 20052
rect 12303 20012 12348 20040
rect 11609 20003 11667 20009
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 15562 20040 15568 20052
rect 15523 20012 15568 20040
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 15896 20012 19533 20040
rect 15896 20000 15902 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 19521 20003 19579 20009
rect 19705 20043 19763 20049
rect 19705 20009 19717 20043
rect 19751 20040 19763 20043
rect 20530 20040 20536 20052
rect 19751 20012 20536 20040
rect 19751 20009 19763 20012
rect 19705 20003 19763 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 22186 20040 22192 20052
rect 22066 20012 22192 20040
rect 13265 19975 13323 19981
rect 13265 19941 13277 19975
rect 13311 19941 13323 19975
rect 13265 19935 13323 19941
rect 13280 19904 13308 19935
rect 18506 19932 18512 19984
rect 18564 19972 18570 19984
rect 22066 19972 22094 20012
rect 22186 20000 22192 20012
rect 22244 20040 22250 20052
rect 32490 20040 32496 20052
rect 22244 20012 32496 20040
rect 22244 20000 22250 20012
rect 32490 20000 32496 20012
rect 32548 20000 32554 20052
rect 43806 20040 43812 20052
rect 38626 20012 43812 20040
rect 18564 19944 22094 19972
rect 25317 19975 25375 19981
rect 18564 19932 18570 19944
rect 25317 19941 25329 19975
rect 25363 19972 25375 19975
rect 25590 19972 25596 19984
rect 25363 19944 25596 19972
rect 25363 19941 25375 19944
rect 25317 19935 25375 19941
rect 25590 19932 25596 19944
rect 25648 19972 25654 19984
rect 25958 19972 25964 19984
rect 25648 19944 25964 19972
rect 25648 19932 25654 19944
rect 25958 19932 25964 19944
rect 26016 19972 26022 19984
rect 26329 19975 26387 19981
rect 26329 19972 26341 19975
rect 26016 19944 26341 19972
rect 26016 19932 26022 19944
rect 26329 19941 26341 19944
rect 26375 19941 26387 19975
rect 26329 19935 26387 19941
rect 36354 19932 36360 19984
rect 36412 19972 36418 19984
rect 38626 19972 38654 20012
rect 43806 20000 43812 20012
rect 43864 20000 43870 20052
rect 43990 20040 43996 20052
rect 43951 20012 43996 20040
rect 43990 20000 43996 20012
rect 44048 20000 44054 20052
rect 36412 19944 38654 19972
rect 36412 19932 36418 19944
rect 42518 19932 42524 19984
rect 42576 19972 42582 19984
rect 46106 19972 46112 19984
rect 42576 19944 46112 19972
rect 42576 19932 42582 19944
rect 46106 19932 46112 19944
rect 46164 19932 46170 19984
rect 12366 19876 13308 19904
rect 16945 19907 17003 19913
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 11790 19836 11796 19848
rect 11751 19808 11796 19836
rect 2041 19799 2099 19805
rect 11790 19796 11796 19808
rect 11848 19796 11854 19848
rect 12366 19845 12394 19876
rect 16945 19873 16957 19907
rect 16991 19904 17003 19907
rect 17218 19904 17224 19916
rect 16991 19876 17224 19904
rect 16991 19873 17003 19876
rect 16945 19867 17003 19873
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 19150 19904 19156 19916
rect 18656 19876 19156 19904
rect 18656 19864 18662 19876
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 20346 19904 20352 19916
rect 20307 19876 20352 19904
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 22005 19907 22063 19913
rect 22005 19873 22017 19907
rect 22051 19904 22063 19907
rect 22051 19876 43576 19904
rect 22051 19873 22063 19876
rect 22005 19867 22063 19873
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19805 12403 19839
rect 12526 19836 12532 19848
rect 12487 19808 12532 19836
rect 12345 19799 12403 19805
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14366 19836 14372 19848
rect 14139 19808 14372 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14366 19796 14372 19808
rect 14424 19836 14430 19848
rect 16850 19836 16856 19848
rect 14424 19808 16856 19836
rect 14424 19796 14430 19808
rect 16850 19796 16856 19808
rect 16908 19796 16914 19848
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19058 19836 19064 19848
rect 18748 19808 19064 19836
rect 18748 19796 18754 19808
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19978 19796 19984 19848
rect 20036 19836 20042 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 20036 19808 20177 19836
rect 20036 19796 20042 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 25682 19796 25688 19848
rect 25740 19836 25746 19848
rect 25740 19808 25785 19836
rect 25740 19796 25746 19808
rect 26234 19796 26240 19848
rect 26292 19836 26298 19848
rect 26605 19839 26663 19845
rect 26605 19836 26617 19839
rect 26292 19808 26617 19836
rect 26292 19796 26298 19808
rect 26605 19805 26617 19808
rect 26651 19805 26663 19839
rect 32398 19836 32404 19848
rect 32359 19808 32404 19836
rect 26605 19799 26663 19805
rect 32398 19796 32404 19808
rect 32456 19796 32462 19848
rect 34701 19839 34759 19845
rect 34701 19805 34713 19839
rect 34747 19805 34759 19839
rect 34701 19799 34759 19805
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 13265 19771 13323 19777
rect 13265 19768 13277 19771
rect 11940 19740 13277 19768
rect 11940 19728 11946 19740
rect 13265 19737 13277 19740
rect 13311 19737 13323 19771
rect 13265 19731 13323 19737
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 15470 19768 15476 19780
rect 15427 19740 15476 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 15597 19771 15655 19777
rect 15597 19737 15609 19771
rect 15643 19768 15655 19771
rect 16758 19768 16764 19780
rect 15643 19740 16764 19768
rect 15643 19737 15655 19740
rect 15597 19731 15655 19737
rect 16758 19728 16764 19740
rect 16816 19728 16822 19780
rect 17218 19768 17224 19780
rect 17179 19740 17224 19768
rect 17218 19728 17224 19740
rect 17276 19728 17282 19780
rect 18966 19768 18972 19780
rect 18446 19740 18972 19768
rect 18966 19728 18972 19740
rect 19024 19728 19030 19780
rect 19334 19768 19340 19780
rect 19295 19740 19340 19768
rect 19334 19728 19340 19740
rect 19392 19728 19398 19780
rect 22554 19768 22560 19780
rect 19444 19740 20392 19768
rect 22515 19740 22560 19768
rect 13449 19703 13507 19709
rect 13449 19669 13461 19703
rect 13495 19700 13507 19703
rect 13814 19700 13820 19712
rect 13495 19672 13820 19700
rect 13495 19669 13507 19672
rect 13449 19663 13507 19669
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 14182 19700 14188 19712
rect 14143 19672 14188 19700
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 15746 19700 15752 19712
rect 15707 19672 15752 19700
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 16390 19660 16396 19712
rect 16448 19700 16454 19712
rect 18046 19700 18052 19712
rect 16448 19672 18052 19700
rect 16448 19660 16454 19672
rect 18046 19660 18052 19672
rect 18104 19700 18110 19712
rect 18690 19700 18696 19712
rect 18104 19672 18696 19700
rect 18104 19660 18110 19672
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 18782 19660 18788 19712
rect 18840 19700 18846 19712
rect 19444 19700 19472 19740
rect 18840 19672 19472 19700
rect 19547 19703 19605 19709
rect 18840 19660 18846 19672
rect 19547 19669 19559 19703
rect 19593 19700 19605 19703
rect 20254 19700 20260 19712
rect 19593 19672 20260 19700
rect 19593 19669 19605 19672
rect 19547 19663 19605 19669
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20364 19700 20392 19740
rect 22554 19728 22560 19740
rect 22612 19728 22618 19780
rect 25501 19771 25559 19777
rect 25501 19737 25513 19771
rect 25547 19768 25559 19771
rect 25774 19768 25780 19780
rect 25547 19740 25780 19768
rect 25547 19737 25559 19740
rect 25501 19731 25559 19737
rect 25774 19728 25780 19740
rect 25832 19728 25838 19780
rect 25866 19728 25872 19780
rect 25924 19768 25930 19780
rect 26326 19768 26332 19780
rect 25924 19740 25969 19768
rect 26176 19740 26332 19768
rect 25924 19728 25930 19740
rect 22186 19700 22192 19712
rect 20364 19672 22192 19700
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 22428 19672 22661 19700
rect 22428 19660 22434 19672
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 22649 19663 22707 19669
rect 25593 19703 25651 19709
rect 25593 19669 25605 19703
rect 25639 19700 25651 19703
rect 26176 19700 26204 19740
rect 26326 19728 26332 19740
rect 26384 19768 26390 19780
rect 26697 19771 26755 19777
rect 26697 19768 26709 19771
rect 26384 19740 26709 19768
rect 26384 19728 26390 19740
rect 26697 19737 26709 19740
rect 26743 19737 26755 19771
rect 34716 19768 34744 19799
rect 35434 19796 35440 19848
rect 35492 19836 35498 19848
rect 42429 19839 42487 19845
rect 35492 19808 41414 19836
rect 35492 19796 35498 19808
rect 36354 19768 36360 19780
rect 34716 19740 36360 19768
rect 26697 19731 26755 19737
rect 36354 19728 36360 19740
rect 36412 19728 36418 19780
rect 26510 19700 26516 19712
rect 25639 19672 26204 19700
rect 26471 19672 26516 19700
rect 25639 19669 25651 19672
rect 25593 19663 25651 19669
rect 26510 19660 26516 19672
rect 26568 19660 26574 19712
rect 26786 19660 26792 19712
rect 26844 19700 26850 19712
rect 26881 19703 26939 19709
rect 26881 19700 26893 19703
rect 26844 19672 26893 19700
rect 26844 19660 26850 19672
rect 26881 19669 26893 19672
rect 26927 19669 26939 19703
rect 26881 19663 26939 19669
rect 32217 19703 32275 19709
rect 32217 19669 32229 19703
rect 32263 19700 32275 19703
rect 33226 19700 33232 19712
rect 32263 19672 33232 19700
rect 32263 19669 32275 19672
rect 32217 19663 32275 19669
rect 33226 19660 33232 19672
rect 33284 19660 33290 19712
rect 33502 19660 33508 19712
rect 33560 19700 33566 19712
rect 34793 19703 34851 19709
rect 34793 19700 34805 19703
rect 33560 19672 34805 19700
rect 33560 19660 33566 19672
rect 34793 19669 34805 19672
rect 34839 19669 34851 19703
rect 41386 19700 41414 19808
rect 42429 19805 42441 19839
rect 42475 19836 42487 19839
rect 42702 19836 42708 19848
rect 42475 19808 42708 19836
rect 42475 19805 42487 19808
rect 42429 19799 42487 19805
rect 42702 19796 42708 19808
rect 42760 19796 42766 19848
rect 42794 19796 42800 19848
rect 42852 19836 42858 19848
rect 42852 19808 42897 19836
rect 42852 19796 42858 19808
rect 42610 19768 42616 19780
rect 42571 19740 42616 19768
rect 42610 19728 42616 19740
rect 42668 19728 42674 19780
rect 43438 19700 43444 19712
rect 41386 19672 43444 19700
rect 34793 19663 34851 19669
rect 43438 19660 43444 19672
rect 43496 19660 43502 19712
rect 43548 19700 43576 19876
rect 43714 19864 43720 19916
rect 43772 19864 43778 19916
rect 43806 19864 43812 19916
rect 43864 19904 43870 19916
rect 46566 19904 46572 19916
rect 43864 19876 46572 19904
rect 43864 19864 43870 19876
rect 46566 19864 46572 19876
rect 46624 19864 46630 19916
rect 43625 19839 43683 19845
rect 43625 19805 43637 19839
rect 43671 19836 43683 19839
rect 43732 19836 43760 19864
rect 43671 19808 43760 19836
rect 45833 19839 45891 19845
rect 43671 19805 43683 19808
rect 43625 19799 43683 19805
rect 45833 19805 45845 19839
rect 45879 19836 45891 19839
rect 46293 19839 46351 19845
rect 46293 19836 46305 19839
rect 45879 19808 46305 19836
rect 45879 19805 45891 19808
rect 45833 19799 45891 19805
rect 46293 19805 46305 19808
rect 46339 19805 46351 19839
rect 46293 19799 46351 19805
rect 43714 19728 43720 19780
rect 43772 19768 43778 19780
rect 43809 19771 43867 19777
rect 43809 19768 43821 19771
rect 43772 19740 43821 19768
rect 43772 19728 43778 19740
rect 43809 19737 43821 19740
rect 43855 19768 43867 19771
rect 43898 19768 43904 19780
rect 43855 19740 43904 19768
rect 43855 19737 43867 19740
rect 43809 19731 43867 19737
rect 43898 19728 43904 19740
rect 43956 19728 43962 19780
rect 46477 19771 46535 19777
rect 46477 19737 46489 19771
rect 46523 19768 46535 19771
rect 47670 19768 47676 19780
rect 46523 19740 47676 19768
rect 46523 19737 46535 19740
rect 46477 19731 46535 19737
rect 47670 19728 47676 19740
rect 47728 19728 47734 19780
rect 48130 19768 48136 19780
rect 48091 19740 48136 19768
rect 48130 19728 48136 19740
rect 48188 19728 48194 19780
rect 45922 19700 45928 19712
rect 43548 19672 45928 19700
rect 45922 19660 45928 19672
rect 45980 19660 45986 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 20073 19499 20131 19505
rect 3476 19468 19840 19496
rect 3476 19456 3482 19468
rect 19812 19440 19840 19468
rect 20073 19465 20085 19499
rect 20119 19496 20131 19499
rect 20119 19468 20300 19496
rect 20119 19465 20131 19468
rect 20073 19459 20131 19465
rect 13722 19428 13728 19440
rect 13188 19400 13728 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 13188 19369 13216 19400
rect 13722 19388 13728 19400
rect 13780 19388 13786 19440
rect 14182 19388 14188 19440
rect 14240 19388 14246 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14936 19400 15393 19428
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19329 13231 19363
rect 13173 19323 13231 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19292 13507 19295
rect 14090 19292 14096 19304
rect 13495 19264 14096 19292
rect 13495 19261 13507 19264
rect 13449 19255 13507 19261
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14936 19301 14964 19400
rect 15381 19397 15393 19400
rect 15427 19397 15439 19431
rect 15381 19391 15439 19397
rect 15562 19388 15568 19440
rect 15620 19437 15626 19440
rect 15620 19431 15639 19437
rect 15627 19397 15639 19431
rect 15620 19391 15639 19397
rect 15620 19388 15626 19391
rect 17218 19388 17224 19440
rect 17276 19428 17282 19440
rect 17405 19431 17463 19437
rect 17405 19428 17417 19431
rect 17276 19400 17417 19428
rect 17276 19388 17282 19400
rect 17405 19397 17417 19400
rect 17451 19397 17463 19431
rect 18782 19428 18788 19440
rect 17405 19391 17463 19397
rect 17512 19400 18788 19428
rect 15838 19360 15844 19372
rect 15028 19332 15844 19360
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14516 19264 14933 19292
rect 14516 19252 14522 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14182 19156 14188 19168
rect 13872 19128 14188 19156
rect 13872 19116 13878 19128
rect 14182 19116 14188 19128
rect 14240 19156 14246 19168
rect 15028 19156 15056 19332
rect 15764 19233 15792 19332
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 16758 19360 16764 19372
rect 16671 19332 16764 19360
rect 16758 19320 16764 19332
rect 16816 19360 16822 19372
rect 17512 19360 17540 19400
rect 18782 19388 18788 19400
rect 18840 19388 18846 19440
rect 19794 19388 19800 19440
rect 19852 19388 19858 19440
rect 19981 19431 20039 19437
rect 19981 19397 19993 19431
rect 20027 19428 20039 19431
rect 20162 19428 20168 19440
rect 20027 19400 20168 19428
rect 20027 19397 20039 19400
rect 19981 19391 20039 19397
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 16816 19332 17540 19360
rect 17589 19363 17647 19369
rect 16816 19320 16822 19332
rect 17589 19329 17601 19363
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19360 17923 19363
rect 17911 19332 18000 19360
rect 17911 19329 17923 19332
rect 17865 19323 17923 19329
rect 17604 19292 17632 19323
rect 16868 19264 17632 19292
rect 17972 19292 18000 19332
rect 18046 19320 18052 19372
rect 18104 19360 18110 19372
rect 18104 19332 18149 19360
rect 18104 19320 18110 19332
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18869 19363 18927 19369
rect 18869 19360 18881 19363
rect 18656 19332 18881 19360
rect 18656 19320 18662 19332
rect 18869 19329 18881 19332
rect 18915 19329 18927 19363
rect 18869 19323 18927 19329
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19116 19332 19717 19360
rect 19116 19320 19122 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19886 19360 19892 19372
rect 19847 19332 19892 19360
rect 19705 19323 19763 19329
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 20272 19360 20300 19468
rect 20530 19456 20536 19508
rect 20588 19496 20594 19508
rect 43070 19496 43076 19508
rect 20588 19468 35204 19496
rect 43031 19468 43076 19496
rect 20588 19456 20594 19468
rect 20622 19388 20628 19440
rect 20680 19428 20686 19440
rect 20901 19431 20959 19437
rect 20901 19428 20913 19431
rect 20680 19400 20913 19428
rect 20680 19388 20686 19400
rect 20901 19397 20913 19400
rect 20947 19397 20959 19431
rect 20901 19391 20959 19397
rect 21821 19431 21879 19437
rect 21821 19397 21833 19431
rect 21867 19397 21879 19431
rect 21821 19391 21879 19397
rect 20806 19360 20812 19372
rect 20272 19332 20812 19360
rect 20806 19320 20812 19332
rect 20864 19360 20870 19372
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20864 19332 21005 19360
rect 20864 19320 20870 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21836 19360 21864 19391
rect 22002 19388 22008 19440
rect 22060 19437 22066 19440
rect 22060 19431 22079 19437
rect 22067 19397 22079 19431
rect 22278 19428 22284 19440
rect 22060 19391 22079 19397
rect 22112 19400 22284 19428
rect 22060 19388 22066 19391
rect 22112 19360 22140 19400
rect 22278 19388 22284 19400
rect 22336 19388 22342 19440
rect 25866 19428 25872 19440
rect 25254 19400 25872 19428
rect 25866 19388 25872 19400
rect 25924 19388 25930 19440
rect 25961 19431 26019 19437
rect 25961 19397 25973 19431
rect 26007 19397 26019 19431
rect 25961 19391 26019 19397
rect 21140 19332 21185 19360
rect 21836 19332 22140 19360
rect 21140 19320 21146 19332
rect 22186 19320 22192 19372
rect 22244 19320 22250 19372
rect 22925 19363 22983 19369
rect 22925 19329 22937 19363
rect 22971 19360 22983 19363
rect 23382 19360 23388 19372
rect 22971 19332 23388 19360
rect 22971 19329 22983 19332
rect 22925 19323 22983 19329
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 23750 19360 23756 19372
rect 23711 19332 23756 19360
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 21269 19295 21327 19301
rect 21269 19292 21281 19295
rect 17972 19264 19104 19292
rect 15749 19227 15807 19233
rect 15749 19193 15761 19227
rect 15795 19193 15807 19227
rect 15749 19187 15807 19193
rect 16868 19168 16896 19264
rect 18966 19224 18972 19236
rect 18927 19196 18972 19224
rect 18966 19184 18972 19196
rect 19024 19184 19030 19236
rect 19076 19224 19104 19264
rect 20272 19264 21281 19292
rect 20272 19224 20300 19264
rect 21269 19261 21281 19264
rect 21315 19261 21327 19295
rect 21269 19255 21327 19261
rect 19076 19196 20300 19224
rect 20717 19227 20775 19233
rect 20717 19193 20729 19227
rect 20763 19224 20775 19227
rect 20990 19224 20996 19236
rect 20763 19196 20996 19224
rect 20763 19193 20775 19196
rect 20717 19187 20775 19193
rect 20990 19184 20996 19196
rect 21048 19184 21054 19236
rect 22204 19233 22232 19320
rect 23017 19295 23075 19301
rect 23017 19261 23029 19295
rect 23063 19261 23075 19295
rect 24029 19295 24087 19301
rect 24029 19292 24041 19295
rect 23017 19255 23075 19261
rect 23860 19264 24041 19292
rect 22189 19227 22247 19233
rect 22189 19193 22201 19227
rect 22235 19193 22247 19227
rect 22189 19187 22247 19193
rect 14240 19128 15056 19156
rect 14240 19116 14246 19128
rect 15470 19116 15476 19168
rect 15528 19156 15534 19168
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 15528 19128 15577 19156
rect 15528 19116 15534 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 16850 19156 16856 19168
rect 16811 19128 16856 19156
rect 15565 19119 15623 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 20254 19156 20260 19168
rect 20167 19128 20260 19156
rect 20254 19116 20260 19128
rect 20312 19156 20318 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 20312 19128 22017 19156
rect 20312 19116 20318 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 23032 19156 23060 19255
rect 23293 19227 23351 19233
rect 23293 19193 23305 19227
rect 23339 19224 23351 19227
rect 23860 19224 23888 19264
rect 24029 19261 24041 19264
rect 24075 19261 24087 19295
rect 25976 19292 26004 19391
rect 26142 19388 26148 19440
rect 26200 19437 26206 19440
rect 26200 19431 26219 19437
rect 26207 19397 26219 19431
rect 32214 19428 32220 19440
rect 32175 19400 32220 19428
rect 26200 19391 26219 19397
rect 26200 19388 26206 19391
rect 32214 19388 32220 19400
rect 32272 19388 32278 19440
rect 32309 19431 32367 19437
rect 32309 19397 32321 19431
rect 32355 19428 32367 19431
rect 33318 19428 33324 19440
rect 32355 19400 33324 19428
rect 32355 19397 32367 19400
rect 32309 19391 32367 19397
rect 33318 19388 33324 19400
rect 33376 19388 33382 19440
rect 33502 19428 33508 19440
rect 33463 19400 33508 19428
rect 33502 19388 33508 19400
rect 33560 19388 33566 19440
rect 35176 19437 35204 19468
rect 43070 19456 43076 19468
rect 43128 19456 43134 19508
rect 43438 19456 43444 19508
rect 43496 19496 43502 19508
rect 45557 19499 45615 19505
rect 43496 19468 45140 19496
rect 43496 19456 43502 19468
rect 35161 19431 35219 19437
rect 35161 19397 35173 19431
rect 35207 19397 35219 19431
rect 35161 19391 35219 19397
rect 42886 19388 42892 19440
rect 42944 19428 42950 19440
rect 45002 19428 45008 19440
rect 42944 19400 44772 19428
rect 44963 19400 45008 19428
rect 42944 19388 42950 19400
rect 26050 19320 26056 19372
rect 26108 19360 26114 19372
rect 26786 19360 26792 19372
rect 26108 19332 26792 19360
rect 26108 19320 26114 19332
rect 26786 19320 26792 19332
rect 26844 19320 26850 19372
rect 42978 19360 42984 19372
rect 42939 19332 42984 19360
rect 42978 19320 42984 19332
rect 43036 19320 43042 19372
rect 43162 19360 43168 19372
rect 43123 19332 43168 19360
rect 43162 19320 43168 19332
rect 43220 19320 43226 19372
rect 43990 19360 43996 19372
rect 43951 19332 43996 19360
rect 43990 19320 43996 19332
rect 44048 19320 44054 19372
rect 44266 19320 44272 19372
rect 44324 19320 44330 19372
rect 44744 19360 44772 19400
rect 45002 19388 45008 19400
rect 45060 19388 45066 19440
rect 45112 19428 45140 19468
rect 45557 19465 45569 19499
rect 45603 19496 45615 19499
rect 45646 19496 45652 19508
rect 45603 19468 45652 19496
rect 45603 19465 45615 19468
rect 45557 19459 45615 19465
rect 45646 19456 45652 19468
rect 45704 19456 45710 19508
rect 47670 19496 47676 19508
rect 47631 19468 47676 19496
rect 47670 19456 47676 19468
rect 47728 19456 47734 19508
rect 46750 19428 46756 19440
rect 45112 19400 46756 19428
rect 46750 19388 46756 19400
rect 46808 19388 46814 19440
rect 45738 19360 45744 19372
rect 44744 19332 45600 19360
rect 45699 19332 45744 19360
rect 26510 19292 26516 19304
rect 25976 19264 26516 19292
rect 24029 19255 24087 19261
rect 26510 19252 26516 19264
rect 26568 19252 26574 19304
rect 32490 19292 32496 19304
rect 32451 19264 32496 19292
rect 32490 19252 32496 19264
rect 32548 19252 32554 19304
rect 33226 19252 33232 19304
rect 33284 19292 33290 19304
rect 33321 19295 33379 19301
rect 33321 19292 33333 19295
rect 33284 19264 33333 19292
rect 33284 19252 33290 19264
rect 33321 19261 33333 19264
rect 33367 19261 33379 19295
rect 45572 19292 45600 19332
rect 45738 19320 45744 19332
rect 45796 19320 45802 19372
rect 46845 19363 46903 19369
rect 46845 19360 46857 19363
rect 45848 19332 46857 19360
rect 45848 19292 45876 19332
rect 46845 19329 46857 19332
rect 46891 19329 46903 19363
rect 46845 19323 46903 19329
rect 47486 19320 47492 19372
rect 47544 19360 47550 19372
rect 47581 19363 47639 19369
rect 47581 19360 47593 19363
rect 47544 19332 47593 19360
rect 47544 19320 47550 19332
rect 47581 19329 47593 19332
rect 47627 19329 47639 19363
rect 47581 19323 47639 19329
rect 45572 19264 45876 19292
rect 33321 19255 33379 19261
rect 26326 19224 26332 19236
rect 23339 19196 23888 19224
rect 26287 19196 26332 19224
rect 23339 19193 23351 19196
rect 23293 19187 23351 19193
rect 26326 19184 26332 19196
rect 26384 19184 26390 19236
rect 25314 19156 25320 19168
rect 23032 19128 25320 19156
rect 22005 19119 22063 19125
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 25498 19156 25504 19168
rect 25459 19128 25504 19156
rect 25498 19116 25504 19128
rect 25556 19156 25562 19168
rect 26145 19159 26203 19165
rect 26145 19156 26157 19159
rect 25556 19128 26157 19156
rect 25556 19116 25562 19128
rect 26145 19125 26157 19128
rect 26191 19125 26203 19159
rect 26145 19119 26203 19125
rect 46290 19116 46296 19168
rect 46348 19156 46354 19168
rect 46385 19159 46443 19165
rect 46385 19156 46397 19159
rect 46348 19128 46397 19156
rect 46348 19116 46354 19128
rect 46385 19125 46397 19128
rect 46431 19125 46443 19159
rect 46934 19156 46940 19168
rect 46895 19128 46940 19156
rect 46385 19119 46443 19125
rect 46934 19116 46940 19128
rect 46992 19116 46998 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 14090 18952 14096 18964
rect 14051 18924 14096 18952
rect 2225 18915 2283 18921
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 14516 18924 14657 18952
rect 14516 18912 14522 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 21082 18952 21088 18964
rect 20995 18924 21088 18952
rect 14645 18915 14703 18921
rect 21082 18912 21088 18924
rect 21140 18952 21146 18964
rect 22373 18955 22431 18961
rect 22373 18952 22385 18955
rect 21140 18924 22385 18952
rect 21140 18912 21146 18924
rect 22373 18921 22385 18924
rect 22419 18921 22431 18955
rect 22373 18915 22431 18921
rect 25866 18912 25872 18964
rect 25924 18952 25930 18964
rect 25961 18955 26019 18961
rect 25961 18952 25973 18955
rect 25924 18924 25973 18952
rect 25924 18912 25930 18924
rect 25961 18921 25973 18924
rect 26007 18921 26019 18955
rect 25961 18915 26019 18921
rect 28905 18955 28963 18961
rect 28905 18921 28917 18955
rect 28951 18952 28963 18955
rect 29822 18952 29828 18964
rect 28951 18924 29828 18952
rect 28951 18921 28963 18924
rect 28905 18915 28963 18921
rect 29822 18912 29828 18924
rect 29880 18952 29886 18964
rect 30282 18952 30288 18964
rect 29880 18924 30288 18952
rect 29880 18912 29886 18924
rect 30282 18912 30288 18924
rect 30340 18912 30346 18964
rect 30745 18955 30803 18961
rect 30745 18921 30757 18955
rect 30791 18952 30803 18955
rect 32398 18952 32404 18964
rect 30791 18924 32404 18952
rect 30791 18921 30803 18924
rect 30745 18915 30803 18921
rect 32398 18912 32404 18924
rect 32456 18912 32462 18964
rect 32582 18952 32588 18964
rect 32543 18924 32588 18952
rect 32582 18912 32588 18924
rect 32640 18912 32646 18964
rect 33318 18952 33324 18964
rect 33279 18924 33324 18952
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 45830 18952 45836 18964
rect 45791 18924 45836 18952
rect 45830 18912 45836 18924
rect 45888 18912 45894 18964
rect 13538 18844 13544 18896
rect 13596 18884 13602 18896
rect 16850 18884 16856 18896
rect 13596 18856 16856 18884
rect 13596 18844 13602 18856
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 14737 18819 14795 18825
rect 4948 18788 14412 18816
rect 4948 18776 4954 18788
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 2314 18748 2320 18760
rect 2179 18720 2320 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 2314 18708 2320 18720
rect 2372 18748 2378 18760
rect 13630 18748 13636 18760
rect 2372 18720 13636 18748
rect 2372 18708 2378 18720
rect 13630 18708 13636 18720
rect 13688 18708 13694 18760
rect 14182 18708 14188 18760
rect 14240 18757 14246 18760
rect 14240 18751 14276 18757
rect 14264 18717 14276 18751
rect 14240 18711 14276 18717
rect 14240 18708 14246 18711
rect 14384 18680 14412 18788
rect 14737 18785 14749 18819
rect 14783 18816 14795 18819
rect 15194 18816 15200 18828
rect 14783 18788 15200 18816
rect 14783 18785 14795 18788
rect 14737 18779 14795 18785
rect 15194 18776 15200 18788
rect 15252 18816 15258 18828
rect 15746 18816 15752 18828
rect 15252 18788 15752 18816
rect 15252 18776 15258 18788
rect 15746 18776 15752 18788
rect 15804 18776 15810 18828
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 15470 18748 15476 18760
rect 15427 18720 15476 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 15657 18751 15715 18757
rect 15657 18717 15669 18751
rect 15703 18748 15715 18751
rect 15856 18748 15884 18856
rect 16850 18844 16856 18856
rect 16908 18844 16914 18896
rect 19886 18844 19892 18896
rect 19944 18884 19950 18896
rect 20990 18884 20996 18896
rect 19944 18856 20996 18884
rect 19944 18844 19950 18856
rect 20990 18844 20996 18856
rect 21048 18844 21054 18896
rect 20714 18776 20720 18828
rect 20772 18816 20778 18828
rect 21100 18825 21128 18912
rect 22094 18844 22100 18896
rect 22152 18844 22158 18896
rect 25222 18844 25228 18896
rect 25280 18884 25286 18896
rect 25774 18884 25780 18896
rect 25280 18856 25780 18884
rect 25280 18844 25286 18856
rect 25774 18844 25780 18856
rect 25832 18844 25838 18896
rect 31849 18887 31907 18893
rect 31849 18884 31861 18887
rect 28828 18856 31861 18884
rect 21085 18819 21143 18825
rect 21085 18816 21097 18819
rect 20772 18788 21097 18816
rect 20772 18776 20778 18788
rect 21085 18785 21097 18788
rect 21131 18785 21143 18819
rect 21542 18816 21548 18828
rect 21503 18788 21548 18816
rect 21085 18779 21143 18785
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 22005 18819 22063 18825
rect 22005 18785 22017 18819
rect 22051 18816 22063 18819
rect 22112 18816 22140 18844
rect 22051 18788 22140 18816
rect 23308 18788 27384 18816
rect 22051 18785 22063 18788
rect 22005 18779 22063 18785
rect 16298 18748 16304 18760
rect 15703 18720 15884 18748
rect 16259 18720 16304 18748
rect 15703 18717 15715 18720
rect 15657 18711 15715 18717
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18748 17647 18751
rect 17954 18748 17960 18760
rect 17635 18720 17960 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 21177 18751 21235 18757
rect 21177 18748 21189 18751
rect 20956 18720 21189 18748
rect 20956 18708 20962 18720
rect 21177 18717 21189 18720
rect 21223 18748 21235 18751
rect 21910 18748 21916 18760
rect 21223 18720 21916 18748
rect 21223 18717 21235 18720
rect 21177 18711 21235 18717
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22094 18708 22100 18760
rect 22152 18748 22158 18760
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 22152 18720 22201 18748
rect 22152 18708 22158 18720
rect 22189 18717 22201 18720
rect 22235 18717 22247 18751
rect 22189 18711 22247 18717
rect 23308 18680 23336 18788
rect 23382 18708 23388 18760
rect 23440 18748 23446 18760
rect 23440 18720 25268 18748
rect 23440 18708 23446 18720
rect 14384 18652 23336 18680
rect 25038 18640 25044 18692
rect 25096 18680 25102 18692
rect 25133 18683 25191 18689
rect 25133 18680 25145 18683
rect 25096 18652 25145 18680
rect 25096 18640 25102 18652
rect 25133 18649 25145 18652
rect 25179 18649 25191 18683
rect 25240 18680 25268 18720
rect 25314 18708 25320 18760
rect 25372 18748 25378 18760
rect 25409 18751 25467 18757
rect 25409 18748 25421 18751
rect 25372 18720 25421 18748
rect 25372 18708 25378 18720
rect 25409 18717 25421 18720
rect 25455 18717 25467 18751
rect 25409 18711 25467 18717
rect 25774 18708 25780 18760
rect 25832 18748 25838 18760
rect 25869 18751 25927 18757
rect 25869 18748 25881 18751
rect 25832 18720 25881 18748
rect 25832 18708 25838 18720
rect 25869 18717 25881 18720
rect 25915 18717 25927 18751
rect 26878 18748 26884 18760
rect 26839 18720 26884 18748
rect 25869 18711 25927 18717
rect 26878 18708 26884 18720
rect 26936 18708 26942 18760
rect 25498 18680 25504 18692
rect 25240 18652 25504 18680
rect 25133 18643 25191 18649
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 13538 18612 13544 18624
rect 13136 18584 13544 18612
rect 13136 18572 13142 18584
rect 13538 18572 13544 18584
rect 13596 18612 13602 18624
rect 14277 18615 14335 18621
rect 14277 18612 14289 18615
rect 13596 18584 14289 18612
rect 13596 18572 13602 18584
rect 14277 18581 14289 18584
rect 14323 18581 14335 18615
rect 14277 18575 14335 18581
rect 15197 18615 15255 18621
rect 15197 18581 15209 18615
rect 15243 18612 15255 18615
rect 15378 18612 15384 18624
rect 15243 18584 15384 18612
rect 15243 18581 15255 18584
rect 15197 18575 15255 18581
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 15562 18612 15568 18624
rect 15523 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15712 18584 16129 18612
rect 15712 18572 15718 18584
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 17678 18612 17684 18624
rect 17639 18584 17684 18612
rect 16117 18575 16175 18581
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 25222 18612 25228 18624
rect 25280 18621 25286 18624
rect 25332 18621 25360 18652
rect 25498 18640 25504 18652
rect 25556 18640 25562 18692
rect 27356 18680 27384 18788
rect 28718 18708 28724 18760
rect 28776 18748 28782 18760
rect 28828 18757 28856 18856
rect 29564 18757 29592 18856
rect 31849 18853 31861 18856
rect 31895 18884 31907 18887
rect 32490 18884 32496 18896
rect 31895 18856 32496 18884
rect 31895 18853 31907 18856
rect 31849 18847 31907 18853
rect 32490 18844 32496 18856
rect 32548 18844 32554 18896
rect 33226 18844 33232 18896
rect 33284 18884 33290 18896
rect 33284 18856 34744 18884
rect 33284 18844 33290 18856
rect 29917 18819 29975 18825
rect 29917 18785 29929 18819
rect 29963 18816 29975 18819
rect 31297 18819 31355 18825
rect 29963 18788 30604 18816
rect 29963 18785 29975 18788
rect 29917 18779 29975 18785
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 28776 18720 28825 18748
rect 28776 18708 28782 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18717 29055 18751
rect 28997 18711 29055 18717
rect 29549 18751 29607 18757
rect 29549 18717 29561 18751
rect 29595 18717 29607 18751
rect 29549 18711 29607 18717
rect 29012 18680 29040 18711
rect 30282 18708 30288 18760
rect 30340 18748 30346 18760
rect 30576 18757 30604 18788
rect 31297 18785 31309 18819
rect 31343 18816 31355 18819
rect 31386 18816 31392 18828
rect 31343 18788 31392 18816
rect 31343 18785 31355 18788
rect 31297 18779 31355 18785
rect 31386 18776 31392 18788
rect 31444 18816 31450 18828
rect 34716 18825 34744 18856
rect 46750 18844 46756 18896
rect 46808 18884 46814 18896
rect 46808 18856 47072 18884
rect 46808 18844 46814 18856
rect 32861 18819 32919 18825
rect 31444 18788 32812 18816
rect 31444 18776 31450 18788
rect 30377 18751 30435 18757
rect 30377 18748 30389 18751
rect 30340 18720 30389 18748
rect 30340 18708 30346 18720
rect 30377 18717 30389 18720
rect 30423 18717 30435 18751
rect 30377 18711 30435 18717
rect 30561 18751 30619 18757
rect 30561 18717 30573 18751
rect 30607 18717 30619 18751
rect 30561 18711 30619 18717
rect 32401 18751 32459 18757
rect 32401 18717 32413 18751
rect 32447 18717 32459 18751
rect 32401 18711 32459 18717
rect 29178 18680 29184 18692
rect 27356 18652 29184 18680
rect 29178 18640 29184 18652
rect 29236 18680 29242 18692
rect 29733 18683 29791 18689
rect 29733 18680 29745 18683
rect 29236 18652 29745 18680
rect 29236 18640 29242 18652
rect 29733 18649 29745 18652
rect 29779 18649 29791 18683
rect 29733 18643 29791 18649
rect 31389 18683 31447 18689
rect 31389 18649 31401 18683
rect 31435 18649 31447 18683
rect 31389 18643 31447 18649
rect 25189 18584 25228 18612
rect 25222 18572 25228 18584
rect 25280 18575 25289 18621
rect 25317 18615 25375 18621
rect 25317 18581 25329 18615
rect 25363 18581 25375 18615
rect 25317 18575 25375 18581
rect 25280 18572 25286 18575
rect 25866 18572 25872 18624
rect 25924 18612 25930 18624
rect 26973 18615 27031 18621
rect 26973 18612 26985 18615
rect 25924 18584 26985 18612
rect 25924 18572 25930 18584
rect 26973 18581 26985 18584
rect 27019 18581 27031 18615
rect 26973 18575 27031 18581
rect 29086 18572 29092 18624
rect 29144 18612 29150 18624
rect 31404 18612 31432 18643
rect 32416 18612 32444 18711
rect 32784 18680 32812 18788
rect 32861 18785 32873 18819
rect 32907 18816 32919 18819
rect 34701 18819 34759 18825
rect 32907 18788 33548 18816
rect 32907 18785 32919 18788
rect 32861 18779 32919 18785
rect 33520 18757 33548 18788
rect 34701 18785 34713 18819
rect 34747 18785 34759 18819
rect 34701 18779 34759 18785
rect 34885 18819 34943 18825
rect 34885 18785 34897 18819
rect 34931 18816 34943 18819
rect 35066 18816 35072 18828
rect 34931 18788 35072 18816
rect 34931 18785 34943 18788
rect 34885 18779 34943 18785
rect 35066 18776 35072 18788
rect 35124 18816 35130 18828
rect 45281 18819 45339 18825
rect 35124 18788 41414 18816
rect 35124 18776 35130 18788
rect 33505 18751 33563 18757
rect 33505 18717 33517 18751
rect 33551 18717 33563 18751
rect 41386 18748 41414 18788
rect 45281 18785 45293 18819
rect 45327 18816 45339 18819
rect 46106 18816 46112 18828
rect 45327 18788 46112 18816
rect 45327 18785 45339 18788
rect 45281 18779 45339 18785
rect 46106 18776 46112 18788
rect 46164 18776 46170 18828
rect 46290 18816 46296 18828
rect 46251 18788 46296 18816
rect 46290 18776 46296 18788
rect 46348 18776 46354 18828
rect 46477 18819 46535 18825
rect 46477 18785 46489 18819
rect 46523 18816 46535 18819
rect 46934 18816 46940 18828
rect 46523 18788 46940 18816
rect 46523 18785 46535 18788
rect 46477 18779 46535 18785
rect 46934 18776 46940 18788
rect 46992 18776 46998 18828
rect 47044 18825 47072 18856
rect 47029 18819 47087 18825
rect 47029 18785 47041 18819
rect 47075 18785 47087 18819
rect 47029 18779 47087 18785
rect 45465 18751 45523 18757
rect 45465 18748 45477 18751
rect 41386 18720 45477 18748
rect 33505 18711 33563 18717
rect 45465 18717 45477 18720
rect 45511 18748 45523 18751
rect 45830 18748 45836 18760
rect 45511 18720 45836 18748
rect 45511 18717 45523 18720
rect 45465 18711 45523 18717
rect 45830 18708 45836 18720
rect 45888 18708 45894 18760
rect 35434 18680 35440 18692
rect 32784 18652 35440 18680
rect 35434 18640 35440 18652
rect 35492 18640 35498 18692
rect 36538 18680 36544 18692
rect 36499 18652 36544 18680
rect 36538 18640 36544 18652
rect 36596 18640 36602 18692
rect 45370 18640 45376 18692
rect 45428 18680 45434 18692
rect 45649 18683 45707 18689
rect 45649 18680 45661 18683
rect 45428 18652 45661 18680
rect 45428 18640 45434 18652
rect 45649 18649 45661 18652
rect 45695 18680 45707 18683
rect 47854 18680 47860 18692
rect 45695 18652 47860 18680
rect 45695 18649 45707 18652
rect 45649 18643 45707 18649
rect 47854 18640 47860 18652
rect 47912 18640 47918 18692
rect 29144 18584 32444 18612
rect 29144 18572 29150 18584
rect 45554 18572 45560 18624
rect 45612 18612 45618 18624
rect 45612 18584 45657 18612
rect 45612 18572 45618 18584
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 4028 18380 31616 18408
rect 4028 18368 4034 18380
rect 15105 18343 15163 18349
rect 15105 18309 15117 18343
rect 15151 18340 15163 18343
rect 15194 18340 15200 18352
rect 15151 18312 15200 18340
rect 15151 18309 15163 18312
rect 15105 18303 15163 18309
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 17678 18340 17684 18352
rect 17639 18312 17684 18340
rect 17678 18300 17684 18312
rect 17736 18300 17742 18352
rect 21542 18300 21548 18352
rect 21600 18340 21606 18352
rect 22097 18343 22155 18349
rect 22097 18340 22109 18343
rect 21600 18312 22109 18340
rect 21600 18300 21606 18312
rect 22097 18309 22109 18312
rect 22143 18309 22155 18343
rect 22097 18303 22155 18309
rect 22738 18300 22744 18352
rect 22796 18300 22802 18352
rect 25866 18340 25872 18352
rect 25148 18312 25872 18340
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 11422 18232 11428 18284
rect 11480 18272 11486 18284
rect 11885 18275 11943 18281
rect 11885 18272 11897 18275
rect 11480 18244 11897 18272
rect 11480 18232 11486 18244
rect 11885 18241 11897 18244
rect 11931 18272 11943 18275
rect 12250 18272 12256 18284
rect 11931 18244 12256 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 25148 18281 25176 18312
rect 25866 18300 25872 18312
rect 25924 18300 25930 18352
rect 31588 18349 31616 18380
rect 35710 18368 35716 18420
rect 35768 18408 35774 18420
rect 45554 18408 45560 18420
rect 35768 18380 45560 18408
rect 35768 18368 35774 18380
rect 45554 18368 45560 18380
rect 45612 18368 45618 18420
rect 31573 18343 31631 18349
rect 31573 18309 31585 18343
rect 31619 18309 31631 18343
rect 31573 18303 31631 18309
rect 41785 18343 41843 18349
rect 41785 18309 41797 18343
rect 41831 18340 41843 18343
rect 42613 18343 42671 18349
rect 42613 18340 42625 18343
rect 41831 18312 42625 18340
rect 41831 18309 41843 18312
rect 41785 18303 41843 18309
rect 42613 18309 42625 18312
rect 42659 18309 42671 18343
rect 42613 18303 42671 18309
rect 25133 18275 25191 18281
rect 15528 18244 17172 18272
rect 15528 18232 15534 18244
rect 17144 18216 17172 18244
rect 25133 18241 25145 18275
rect 25179 18241 25191 18275
rect 25133 18235 25191 18241
rect 25222 18232 25228 18284
rect 25280 18272 25286 18284
rect 25777 18275 25835 18281
rect 25777 18272 25789 18275
rect 25280 18244 25789 18272
rect 25280 18232 25286 18244
rect 25777 18241 25789 18244
rect 25823 18241 25835 18275
rect 25777 18235 25835 18241
rect 25961 18275 26019 18281
rect 25961 18241 25973 18275
rect 26007 18272 26019 18275
rect 26050 18272 26056 18284
rect 26007 18244 26056 18272
rect 26007 18241 26019 18244
rect 25961 18235 26019 18241
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 28994 18272 29000 18284
rect 28955 18244 29000 18272
rect 28994 18232 29000 18244
rect 29052 18232 29058 18284
rect 29181 18275 29239 18281
rect 29181 18241 29193 18275
rect 29227 18272 29239 18275
rect 29454 18272 29460 18284
rect 29227 18244 29460 18272
rect 29227 18241 29239 18244
rect 29181 18235 29239 18241
rect 29454 18232 29460 18244
rect 29512 18232 29518 18284
rect 35066 18272 35072 18284
rect 35027 18244 35072 18272
rect 35066 18232 35072 18244
rect 35124 18272 35130 18284
rect 35434 18272 35440 18284
rect 35124 18244 35440 18272
rect 35124 18232 35130 18244
rect 35434 18232 35440 18244
rect 35492 18232 35498 18284
rect 38102 18232 38108 18284
rect 38160 18272 38166 18284
rect 41693 18275 41751 18281
rect 41693 18272 41705 18275
rect 38160 18244 41705 18272
rect 38160 18232 38166 18244
rect 41693 18241 41705 18244
rect 41739 18241 41751 18275
rect 41693 18235 41751 18241
rect 45097 18275 45155 18281
rect 45097 18241 45109 18275
rect 45143 18272 45155 18275
rect 45370 18272 45376 18284
rect 45143 18244 45376 18272
rect 45143 18241 45155 18244
rect 45097 18235 45155 18241
rect 45370 18232 45376 18244
rect 45428 18232 45434 18284
rect 45572 18281 45600 18368
rect 45557 18275 45615 18281
rect 45557 18241 45569 18275
rect 45603 18241 45615 18275
rect 45830 18272 45836 18284
rect 45743 18244 45836 18272
rect 45557 18235 45615 18241
rect 45830 18232 45836 18244
rect 45888 18232 45894 18284
rect 46106 18272 46112 18284
rect 46019 18244 46112 18272
rect 46106 18232 46112 18244
rect 46164 18272 46170 18284
rect 46164 18244 46336 18272
rect 46164 18232 46170 18244
rect 13078 18204 13084 18216
rect 13039 18176 13084 18204
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 16298 18204 16304 18216
rect 15611 18176 16304 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17497 18207 17555 18213
rect 17497 18204 17509 18207
rect 17184 18176 17509 18204
rect 17184 18164 17190 18176
rect 17497 18173 17509 18176
rect 17543 18173 17555 18207
rect 19150 18204 19156 18216
rect 19111 18176 19156 18204
rect 17497 18167 17555 18173
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 21821 18207 21879 18213
rect 21821 18173 21833 18207
rect 21867 18173 21879 18207
rect 21821 18167 21879 18173
rect 2041 18139 2099 18145
rect 2041 18105 2053 18139
rect 2087 18136 2099 18139
rect 15378 18136 15384 18148
rect 2087 18108 14596 18136
rect 15339 18108 15384 18136
rect 2087 18105 2099 18108
rect 2041 18099 2099 18105
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 11977 18071 12035 18077
rect 11977 18068 11989 18071
rect 11940 18040 11989 18068
rect 11940 18028 11946 18040
rect 11977 18037 11989 18040
rect 12023 18037 12035 18071
rect 13354 18068 13360 18080
rect 13315 18040 13360 18068
rect 11977 18031 12035 18037
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 14458 18068 14464 18080
rect 14419 18040 14464 18068
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 14568 18068 14596 18108
rect 15378 18096 15384 18108
rect 15436 18096 15442 18148
rect 17034 18068 17040 18080
rect 14568 18040 17040 18068
rect 17034 18028 17040 18040
rect 17092 18028 17098 18080
rect 21836 18068 21864 18167
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 23842 18204 23848 18216
rect 22152 18176 23848 18204
rect 22152 18164 22158 18176
rect 23842 18164 23848 18176
rect 23900 18164 23906 18216
rect 25038 18164 25044 18216
rect 25096 18204 25102 18216
rect 26510 18204 26516 18216
rect 25096 18176 26516 18204
rect 25096 18164 25102 18176
rect 26510 18164 26516 18176
rect 26568 18204 26574 18216
rect 26786 18204 26792 18216
rect 26568 18176 26792 18204
rect 26568 18164 26574 18176
rect 26786 18164 26792 18176
rect 26844 18164 26850 18216
rect 29733 18207 29791 18213
rect 29733 18173 29745 18207
rect 29779 18173 29791 18207
rect 29733 18167 29791 18173
rect 29917 18207 29975 18213
rect 29917 18173 29929 18207
rect 29963 18204 29975 18207
rect 31202 18204 31208 18216
rect 29963 18176 31208 18204
rect 29963 18173 29975 18176
rect 29917 18167 29975 18173
rect 29748 18136 29776 18167
rect 31202 18164 31208 18176
rect 31260 18164 31266 18216
rect 32769 18207 32827 18213
rect 32769 18204 32781 18207
rect 31726 18176 32781 18204
rect 30650 18136 30656 18148
rect 29748 18108 30656 18136
rect 30650 18096 30656 18108
rect 30708 18136 30714 18148
rect 31726 18136 31754 18176
rect 32769 18173 32781 18176
rect 32815 18173 32827 18207
rect 32769 18167 32827 18173
rect 32953 18207 33011 18213
rect 32953 18173 32965 18207
rect 32999 18204 33011 18207
rect 33870 18204 33876 18216
rect 32999 18176 33876 18204
rect 32999 18173 33011 18176
rect 32953 18167 33011 18173
rect 33870 18164 33876 18176
rect 33928 18164 33934 18216
rect 33965 18207 34023 18213
rect 33965 18173 33977 18207
rect 34011 18204 34023 18207
rect 36538 18204 36544 18216
rect 34011 18176 36544 18204
rect 34011 18173 34023 18176
rect 33965 18167 34023 18173
rect 30708 18108 31754 18136
rect 30708 18096 30714 18108
rect 32858 18096 32864 18148
rect 32916 18136 32922 18148
rect 33980 18136 34008 18167
rect 36538 18164 36544 18176
rect 36596 18164 36602 18216
rect 42429 18207 42487 18213
rect 42429 18173 42441 18207
rect 42475 18204 42487 18207
rect 43530 18204 43536 18216
rect 42475 18176 43536 18204
rect 42475 18173 42487 18176
rect 42429 18167 42487 18173
rect 43530 18164 43536 18176
rect 43588 18164 43594 18216
rect 43898 18204 43904 18216
rect 43859 18176 43904 18204
rect 43898 18164 43904 18176
rect 43956 18164 43962 18216
rect 45848 18204 45876 18232
rect 46198 18204 46204 18216
rect 45848 18176 46204 18204
rect 46198 18164 46204 18176
rect 46256 18164 46262 18216
rect 46308 18204 46336 18244
rect 47394 18232 47400 18284
rect 47452 18272 47458 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47452 18244 47593 18272
rect 47452 18232 47458 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 48038 18204 48044 18216
rect 46308 18176 48044 18204
rect 32916 18108 34008 18136
rect 32916 18096 32922 18108
rect 34514 18096 34520 18148
rect 34572 18136 34578 18148
rect 35529 18139 35587 18145
rect 35529 18136 35541 18139
rect 34572 18108 35541 18136
rect 34572 18096 34578 18108
rect 35529 18105 35541 18108
rect 35575 18105 35587 18139
rect 46308 18136 46336 18176
rect 48038 18164 48044 18176
rect 48096 18164 48102 18216
rect 35529 18099 35587 18105
rect 41386 18108 46336 18136
rect 22094 18068 22100 18080
rect 21836 18040 22100 18068
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 25038 18068 25044 18080
rect 24999 18040 25044 18068
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 25314 18028 25320 18080
rect 25372 18068 25378 18080
rect 25777 18071 25835 18077
rect 25777 18068 25789 18071
rect 25372 18040 25789 18068
rect 25372 18028 25378 18040
rect 25777 18037 25789 18040
rect 25823 18037 25835 18071
rect 25777 18031 25835 18037
rect 29089 18071 29147 18077
rect 29089 18037 29101 18071
rect 29135 18068 29147 18071
rect 29730 18068 29736 18080
rect 29135 18040 29736 18068
rect 29135 18037 29147 18040
rect 29089 18031 29147 18037
rect 29730 18028 29736 18040
rect 29788 18028 29794 18080
rect 35342 18068 35348 18080
rect 35255 18040 35348 18068
rect 35342 18028 35348 18040
rect 35400 18068 35406 18080
rect 41386 18068 41414 18108
rect 45554 18068 45560 18080
rect 35400 18040 41414 18068
rect 45515 18040 45560 18068
rect 35400 18028 35406 18040
rect 45554 18028 45560 18040
rect 45612 18028 45618 18080
rect 47026 18068 47032 18080
rect 46987 18040 47032 18068
rect 47026 18028 47032 18040
rect 47084 18028 47090 18080
rect 47670 18068 47676 18080
rect 47631 18040 47676 18068
rect 47670 18028 47676 18040
rect 47728 18028 47734 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 16666 17864 16672 17876
rect 14936 17836 16672 17864
rect 3970 17756 3976 17808
rect 4028 17796 4034 17808
rect 4028 17768 12204 17796
rect 4028 17756 4034 17768
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 11701 17731 11759 17737
rect 11701 17728 11713 17731
rect 11664 17700 11713 17728
rect 11664 17688 11670 17700
rect 11701 17697 11713 17700
rect 11747 17697 11759 17731
rect 11882 17728 11888 17740
rect 11843 17700 11888 17728
rect 11701 17691 11759 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 12176 17737 12204 17768
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17697 12219 17731
rect 12161 17691 12219 17697
rect 12250 17688 12256 17740
rect 12308 17728 12314 17740
rect 14936 17728 14964 17836
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 17126 17864 17132 17876
rect 17087 17836 17132 17864
rect 17126 17824 17132 17836
rect 17184 17824 17190 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22738 17864 22744 17876
rect 22152 17836 22197 17864
rect 22699 17836 22744 17864
rect 22152 17824 22158 17836
rect 22738 17824 22744 17836
rect 22796 17824 22802 17876
rect 26786 17864 26792 17876
rect 24872 17836 26464 17864
rect 26747 17836 26792 17864
rect 15654 17728 15660 17740
rect 12308 17700 14780 17728
rect 12308 17688 12314 17700
rect 14752 17524 14780 17700
rect 14844 17700 14964 17728
rect 15615 17700 15660 17728
rect 14844 17669 14872 17700
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 18874 17728 18880 17740
rect 17788 17700 18880 17728
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17660 14979 17663
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 14967 17632 15393 17660
rect 14967 17629 14979 17632
rect 14921 17623 14979 17629
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15381 17623 15439 17629
rect 16758 17620 16764 17672
rect 16816 17620 16822 17672
rect 17788 17524 17816 17700
rect 18874 17688 18880 17700
rect 18932 17728 18938 17740
rect 22370 17728 22376 17740
rect 18932 17700 22376 17728
rect 18932 17688 18938 17700
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 17920 17632 19257 17660
rect 17920 17620 17926 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 21174 17620 21180 17672
rect 21232 17660 21238 17672
rect 21913 17663 21971 17669
rect 21913 17660 21925 17663
rect 21232 17632 21925 17660
rect 21232 17620 21238 17632
rect 21913 17629 21925 17632
rect 21959 17629 21971 17663
rect 22646 17660 22652 17672
rect 22607 17632 22652 17660
rect 21913 17623 21971 17629
rect 22646 17620 22652 17632
rect 22704 17620 22710 17672
rect 24394 17660 24400 17672
rect 24307 17632 24400 17660
rect 24394 17620 24400 17632
rect 24452 17660 24458 17672
rect 24872 17660 24900 17836
rect 26436 17796 26464 17836
rect 26786 17824 26792 17836
rect 26844 17824 26850 17876
rect 31202 17864 31208 17876
rect 31163 17836 31208 17864
rect 31202 17824 31208 17836
rect 31260 17824 31266 17876
rect 33870 17864 33876 17876
rect 33831 17836 33876 17864
rect 33870 17824 33876 17836
rect 33928 17824 33934 17876
rect 35710 17824 35716 17876
rect 35768 17864 35774 17876
rect 36081 17867 36139 17873
rect 36081 17864 36093 17867
rect 35768 17836 36093 17864
rect 35768 17824 35774 17836
rect 36081 17833 36093 17836
rect 36127 17833 36139 17867
rect 36081 17827 36139 17833
rect 43990 17824 43996 17876
rect 44048 17864 44054 17876
rect 45649 17867 45707 17873
rect 45649 17864 45661 17867
rect 44048 17836 45661 17864
rect 44048 17824 44054 17836
rect 45649 17833 45661 17836
rect 45695 17833 45707 17867
rect 45649 17827 45707 17833
rect 26436 17768 31754 17796
rect 25038 17728 25044 17740
rect 24999 17700 25044 17728
rect 25038 17688 25044 17700
rect 25096 17688 25102 17740
rect 25314 17728 25320 17740
rect 25275 17700 25320 17728
rect 25314 17688 25320 17700
rect 25372 17688 25378 17740
rect 28718 17728 28724 17740
rect 28679 17700 28724 17728
rect 28718 17688 28724 17700
rect 28776 17688 28782 17740
rect 29822 17688 29828 17740
rect 29880 17728 29886 17740
rect 30650 17728 30656 17740
rect 29880 17700 29925 17728
rect 30611 17700 30656 17728
rect 29880 17688 29886 17700
rect 30650 17688 30656 17700
rect 30708 17688 30714 17740
rect 31726 17728 31754 17768
rect 35066 17756 35072 17808
rect 35124 17796 35130 17808
rect 35253 17799 35311 17805
rect 35253 17796 35265 17799
rect 35124 17768 35265 17796
rect 35124 17756 35130 17768
rect 35253 17765 35265 17768
rect 35299 17765 35311 17799
rect 44634 17796 44640 17808
rect 35253 17759 35311 17765
rect 41386 17768 44640 17796
rect 41386 17728 41414 17768
rect 44634 17756 44640 17768
rect 44692 17756 44698 17808
rect 44453 17731 44511 17737
rect 44453 17728 44465 17731
rect 31726 17700 41414 17728
rect 43456 17700 44465 17728
rect 29736 17672 29788 17678
rect 28350 17660 28356 17672
rect 24452 17632 24900 17660
rect 28311 17632 28356 17660
rect 24452 17620 24458 17632
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 28445 17663 28503 17669
rect 28445 17629 28457 17663
rect 28491 17660 28503 17663
rect 28534 17660 28540 17672
rect 28491 17632 28540 17660
rect 28491 17629 28503 17632
rect 28445 17623 28503 17629
rect 28534 17620 28540 17632
rect 28592 17620 28598 17672
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17660 28687 17663
rect 29178 17660 29184 17672
rect 28675 17632 29184 17660
rect 28675 17629 28687 17632
rect 28629 17623 28687 17629
rect 29178 17620 29184 17632
rect 29236 17620 29242 17672
rect 31110 17660 31116 17672
rect 31071 17632 31116 17660
rect 31110 17620 31116 17632
rect 31168 17620 31174 17672
rect 34057 17663 34115 17669
rect 34057 17629 34069 17663
rect 34103 17660 34115 17663
rect 34514 17660 34520 17672
rect 34103 17632 34520 17660
rect 34103 17629 34115 17632
rect 34057 17623 34115 17629
rect 34514 17620 34520 17632
rect 34572 17620 34578 17672
rect 35161 17663 35219 17669
rect 35161 17629 35173 17663
rect 35207 17629 35219 17663
rect 35342 17660 35348 17672
rect 35303 17632 35348 17660
rect 35161 17623 35219 17629
rect 29736 17614 29788 17620
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19521 17595 19579 17601
rect 19521 17592 19533 17595
rect 19484 17564 19533 17592
rect 19484 17552 19490 17564
rect 19521 17561 19533 17564
rect 19567 17561 19579 17595
rect 19521 17555 19579 17561
rect 20162 17552 20168 17604
rect 20220 17552 20226 17604
rect 26050 17552 26056 17604
rect 26108 17552 26114 17604
rect 35176 17592 35204 17623
rect 35342 17620 35348 17632
rect 35400 17620 35406 17672
rect 35434 17620 35440 17672
rect 35492 17660 35498 17672
rect 43456 17669 43484 17700
rect 44453 17697 44465 17700
rect 44499 17728 44511 17731
rect 45005 17731 45063 17737
rect 45005 17728 45017 17731
rect 44499 17700 45017 17728
rect 44499 17697 44511 17700
rect 44453 17691 44511 17697
rect 45005 17697 45017 17700
rect 45051 17697 45063 17731
rect 45005 17691 45063 17697
rect 46293 17731 46351 17737
rect 46293 17697 46305 17731
rect 46339 17728 46351 17731
rect 47026 17728 47032 17740
rect 46339 17700 47032 17728
rect 46339 17697 46351 17700
rect 46293 17691 46351 17697
rect 47026 17688 47032 17700
rect 47084 17688 47090 17740
rect 43441 17663 43499 17669
rect 35492 17632 35537 17660
rect 35492 17620 35498 17632
rect 43441 17629 43453 17663
rect 43487 17629 43499 17663
rect 43441 17623 43499 17629
rect 43625 17663 43683 17669
rect 43625 17629 43637 17663
rect 43671 17660 43683 17663
rect 45370 17660 45376 17672
rect 43671 17632 45376 17660
rect 43671 17629 43683 17632
rect 43625 17623 43683 17629
rect 45370 17620 45376 17632
rect 45428 17620 45434 17672
rect 45465 17663 45523 17669
rect 45465 17629 45477 17663
rect 45511 17629 45523 17663
rect 45465 17623 45523 17629
rect 35710 17592 35716 17604
rect 35176 17564 35716 17592
rect 35710 17552 35716 17564
rect 35768 17552 35774 17604
rect 44082 17592 44088 17604
rect 44043 17564 44088 17592
rect 44082 17552 44088 17564
rect 44140 17552 44146 17604
rect 44269 17595 44327 17601
rect 44269 17561 44281 17595
rect 44315 17561 44327 17595
rect 44269 17555 44327 17561
rect 20990 17524 20996 17536
rect 14752 17496 17816 17524
rect 20951 17496 20996 17524
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 23658 17484 23664 17536
rect 23716 17524 23722 17536
rect 24489 17527 24547 17533
rect 24489 17524 24501 17527
rect 23716 17496 24501 17524
rect 23716 17484 23722 17496
rect 24489 17493 24501 17496
rect 24535 17493 24547 17527
rect 24489 17487 24547 17493
rect 28626 17484 28632 17536
rect 28684 17524 28690 17536
rect 28721 17527 28779 17533
rect 28721 17524 28733 17527
rect 28684 17496 28733 17524
rect 28684 17484 28690 17496
rect 28721 17493 28733 17496
rect 28767 17524 28779 17527
rect 28810 17524 28816 17536
rect 28767 17496 28816 17524
rect 28767 17493 28779 17496
rect 28721 17487 28779 17493
rect 28810 17484 28816 17496
rect 28868 17484 28874 17536
rect 31110 17484 31116 17536
rect 31168 17524 31174 17536
rect 39206 17524 39212 17536
rect 31168 17496 39212 17524
rect 31168 17484 31174 17496
rect 39206 17484 39212 17496
rect 39264 17484 39270 17536
rect 43622 17524 43628 17536
rect 43583 17496 43628 17524
rect 43622 17484 43628 17496
rect 43680 17484 43686 17536
rect 44284 17524 44312 17555
rect 45278 17552 45284 17604
rect 45336 17592 45342 17604
rect 45480 17592 45508 17623
rect 45646 17620 45652 17672
rect 45704 17620 45710 17672
rect 45664 17592 45692 17620
rect 45336 17564 45508 17592
rect 45572 17564 45692 17592
rect 46477 17595 46535 17601
rect 45336 17552 45342 17564
rect 45572 17524 45600 17564
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 47670 17592 47676 17604
rect 46523 17564 47676 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 47670 17552 47676 17564
rect 47728 17552 47734 17604
rect 48133 17595 48191 17601
rect 48133 17561 48145 17595
rect 48179 17592 48191 17595
rect 48222 17592 48228 17604
rect 48179 17564 48228 17592
rect 48179 17561 48191 17564
rect 48133 17555 48191 17561
rect 48222 17552 48228 17564
rect 48280 17552 48286 17604
rect 44284 17496 45600 17524
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 16758 17320 16764 17332
rect 5500 17292 16620 17320
rect 16719 17292 16764 17320
rect 5500 17280 5506 17292
rect 13354 17212 13360 17264
rect 13412 17252 13418 17264
rect 13725 17255 13783 17261
rect 13725 17252 13737 17255
rect 13412 17224 13737 17252
rect 13412 17212 13418 17224
rect 13725 17221 13737 17224
rect 13771 17221 13783 17255
rect 13725 17215 13783 17221
rect 14458 17212 14464 17264
rect 14516 17212 14522 17264
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17184 12035 17187
rect 12250 17184 12256 17196
rect 12023 17156 12256 17184
rect 12023 17153 12035 17156
rect 11977 17147 12035 17153
rect 12250 17144 12256 17156
rect 12308 17144 12314 17196
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17116 13507 17119
rect 14182 17116 14188 17128
rect 13495 17088 14188 17116
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 12069 16983 12127 16989
rect 12069 16980 12081 16983
rect 11940 16952 12081 16980
rect 11940 16940 11946 16952
rect 12069 16949 12081 16952
rect 12115 16949 12127 16983
rect 12069 16943 12127 16949
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 13044 16952 15209 16980
rect 13044 16940 13050 16952
rect 15197 16949 15209 16952
rect 15243 16980 15255 16983
rect 15562 16980 15568 16992
rect 15243 16952 15568 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 16592 16980 16620 17292
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 17862 17320 17868 17332
rect 17823 17292 17868 17320
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 20070 17280 20076 17332
rect 20128 17320 20134 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 20128 17292 21097 17320
rect 20128 17280 20134 17292
rect 21085 17289 21097 17292
rect 21131 17289 21143 17323
rect 21085 17283 21143 17289
rect 26050 17280 26056 17332
rect 26108 17320 26114 17332
rect 26145 17323 26203 17329
rect 26145 17320 26157 17323
rect 26108 17292 26157 17320
rect 26108 17280 26114 17292
rect 26145 17289 26157 17292
rect 26191 17289 26203 17323
rect 28718 17320 28724 17332
rect 28679 17292 28724 17320
rect 26145 17283 26203 17289
rect 28718 17280 28724 17292
rect 28776 17280 28782 17332
rect 28810 17280 28816 17332
rect 28868 17320 28874 17332
rect 28868 17292 29684 17320
rect 28868 17280 28874 17292
rect 16942 17252 16948 17264
rect 16684 17224 16948 17252
rect 16684 17193 16712 17224
rect 16942 17212 16948 17224
rect 17000 17212 17006 17264
rect 20346 17212 20352 17264
rect 20404 17252 20410 17264
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 20404 17224 20729 17252
rect 20404 17212 20410 17224
rect 20717 17221 20729 17224
rect 20763 17221 20775 17255
rect 20917 17255 20975 17261
rect 20917 17252 20929 17255
rect 20717 17215 20775 17221
rect 20916 17221 20929 17252
rect 20963 17221 20975 17255
rect 23658 17252 23664 17264
rect 23619 17224 23664 17252
rect 20916 17215 20975 17221
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 17678 17184 17684 17196
rect 16816 17156 17684 17184
rect 16816 17144 16822 17156
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 20916 17184 20944 17215
rect 23658 17212 23664 17224
rect 23716 17212 23722 17264
rect 23842 17212 23848 17264
rect 23900 17252 23906 17264
rect 27890 17252 27896 17264
rect 23900 17224 27896 17252
rect 23900 17212 23906 17224
rect 27890 17212 27896 17224
rect 27948 17212 27954 17264
rect 28626 17252 28632 17264
rect 28587 17224 28632 17252
rect 28626 17212 28632 17224
rect 28684 17212 28690 17264
rect 19918 17156 20024 17184
rect 19996 17128 20024 17156
rect 20732 17156 20944 17184
rect 21821 17187 21879 17193
rect 20732 17128 20760 17156
rect 21821 17153 21833 17187
rect 21867 17184 21879 17187
rect 22370 17184 22376 17196
rect 21867 17156 22376 17184
rect 21867 17153 21879 17156
rect 21821 17147 21879 17153
rect 22370 17144 22376 17156
rect 22428 17144 22434 17196
rect 23382 17144 23388 17196
rect 23440 17184 23446 17196
rect 23477 17187 23535 17193
rect 23477 17184 23489 17187
rect 23440 17156 23489 17184
rect 23440 17144 23446 17156
rect 23477 17153 23489 17156
rect 23523 17153 23535 17187
rect 23477 17147 23535 17153
rect 25774 17144 25780 17196
rect 25832 17184 25838 17196
rect 26050 17184 26056 17196
rect 25832 17156 26056 17184
rect 25832 17144 25838 17156
rect 26050 17144 26056 17156
rect 26108 17144 26114 17196
rect 27522 17184 27528 17196
rect 26160 17156 27528 17184
rect 18506 17116 18512 17128
rect 18467 17088 18512 17116
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 18785 17119 18843 17125
rect 18785 17085 18797 17119
rect 18831 17116 18843 17119
rect 19334 17116 19340 17128
rect 18831 17088 19340 17116
rect 18831 17085 18843 17088
rect 18785 17079 18843 17085
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 19978 17076 19984 17128
rect 20036 17076 20042 17128
rect 20257 17119 20315 17125
rect 20257 17085 20269 17119
rect 20303 17116 20315 17119
rect 20346 17116 20352 17128
rect 20303 17088 20352 17116
rect 20303 17085 20315 17088
rect 20257 17079 20315 17085
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 20714 17076 20720 17128
rect 20772 17076 20778 17128
rect 25314 17116 25320 17128
rect 25275 17088 25320 17116
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 26160 17048 26188 17156
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 27706 17184 27712 17196
rect 27667 17156 27712 17184
rect 27706 17144 27712 17156
rect 27764 17144 27770 17196
rect 28853 17187 28911 17193
rect 28853 17184 28865 17187
rect 28828 17153 28865 17184
rect 28899 17153 28911 17187
rect 28828 17147 28911 17153
rect 28997 17187 29055 17193
rect 28997 17153 29009 17187
rect 29043 17184 29055 17187
rect 29086 17184 29092 17196
rect 29043 17156 29092 17184
rect 29043 17153 29055 17156
rect 28997 17147 29055 17153
rect 27617 17119 27675 17125
rect 27617 17085 27629 17119
rect 27663 17116 27675 17119
rect 28828 17116 28856 17147
rect 29086 17144 29092 17156
rect 29144 17144 29150 17196
rect 29656 17193 29684 17292
rect 36538 17280 36544 17332
rect 36596 17320 36602 17332
rect 41874 17320 41880 17332
rect 36596 17292 41880 17320
rect 36596 17280 36602 17292
rect 41874 17280 41880 17292
rect 41932 17320 41938 17332
rect 45738 17320 45744 17332
rect 41932 17292 45744 17320
rect 41932 17280 41938 17292
rect 45738 17280 45744 17292
rect 45796 17280 45802 17332
rect 35066 17252 35072 17264
rect 35027 17224 35072 17252
rect 35066 17212 35072 17224
rect 35124 17212 35130 17264
rect 44266 17252 44272 17264
rect 44227 17224 44272 17252
rect 44266 17212 44272 17224
rect 44324 17212 44330 17264
rect 45189 17255 45247 17261
rect 45189 17221 45201 17255
rect 45235 17252 45247 17255
rect 45554 17252 45560 17264
rect 45235 17224 45560 17252
rect 45235 17221 45247 17224
rect 45189 17215 45247 17221
rect 45554 17212 45560 17224
rect 45612 17212 45618 17264
rect 43628 17196 43680 17202
rect 29641 17187 29699 17193
rect 29288 17156 29592 17184
rect 29288 17116 29316 17156
rect 29454 17116 29460 17128
rect 27663 17088 29316 17116
rect 29415 17088 29460 17116
rect 27663 17085 27675 17088
rect 27617 17079 27675 17085
rect 29454 17076 29460 17088
rect 29512 17076 29518 17128
rect 29564 17116 29592 17156
rect 29641 17153 29653 17187
rect 29687 17153 29699 17187
rect 29641 17147 29699 17153
rect 30285 17187 30343 17193
rect 30285 17153 30297 17187
rect 30331 17153 30343 17187
rect 30285 17147 30343 17153
rect 30300 17116 30328 17147
rect 44284 17184 44312 17212
rect 45005 17187 45063 17193
rect 45005 17184 45017 17187
rect 44284 17156 45017 17184
rect 45005 17153 45017 17156
rect 45051 17153 45063 17187
rect 47578 17184 47584 17196
rect 47539 17156 47584 17184
rect 45005 17147 45063 17153
rect 47578 17144 47584 17156
rect 47636 17144 47642 17196
rect 43628 17138 43680 17144
rect 29564 17088 30328 17116
rect 30650 17076 30656 17128
rect 30708 17116 30714 17128
rect 34885 17119 34943 17125
rect 34885 17116 34897 17119
rect 30708 17088 34897 17116
rect 30708 17076 30714 17088
rect 34885 17085 34897 17088
rect 34931 17085 34943 17119
rect 36538 17116 36544 17128
rect 36499 17088 36544 17116
rect 34885 17079 34943 17085
rect 19812 17020 26188 17048
rect 28445 17051 28503 17057
rect 19812 16980 19840 17020
rect 28445 17017 28457 17051
rect 28491 17048 28503 17051
rect 34900 17048 34928 17079
rect 36538 17076 36544 17088
rect 36596 17076 36602 17128
rect 43717 17119 43775 17125
rect 43717 17085 43729 17119
rect 43763 17116 43775 17119
rect 45278 17116 45284 17128
rect 43763 17088 45284 17116
rect 43763 17085 43775 17088
rect 43717 17079 43775 17085
rect 42518 17048 42524 17060
rect 28491 17020 31754 17048
rect 34900 17020 42524 17048
rect 28491 17017 28503 17020
rect 28445 17011 28503 17017
rect 20898 16980 20904 16992
rect 16592 16952 19840 16980
rect 20859 16952 20904 16980
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 21358 16940 21364 16992
rect 21416 16980 21422 16992
rect 21913 16983 21971 16989
rect 21913 16980 21925 16983
rect 21416 16952 21925 16980
rect 21416 16940 21422 16952
rect 21913 16949 21925 16952
rect 21959 16949 21971 16983
rect 21913 16943 21971 16949
rect 24854 16940 24860 16992
rect 24912 16980 24918 16992
rect 25038 16980 25044 16992
rect 24912 16952 25044 16980
rect 24912 16940 24918 16952
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 28718 16940 28724 16992
rect 28776 16980 28782 16992
rect 29454 16980 29460 16992
rect 28776 16952 29460 16980
rect 28776 16940 28782 16952
rect 29454 16940 29460 16952
rect 29512 16940 29518 16992
rect 29822 16980 29828 16992
rect 29783 16952 29828 16980
rect 29822 16940 29828 16952
rect 29880 16940 29886 16992
rect 30374 16980 30380 16992
rect 30335 16952 30380 16980
rect 30374 16940 30380 16952
rect 30432 16940 30438 16992
rect 31726 16980 31754 17020
rect 42518 17008 42524 17020
rect 42576 17008 42582 17060
rect 43732 17048 43760 17079
rect 45278 17076 45284 17088
rect 45336 17076 45342 17128
rect 45738 17116 45744 17128
rect 45699 17088 45744 17116
rect 45738 17076 45744 17088
rect 45796 17076 45802 17128
rect 43364 17020 43760 17048
rect 43364 16980 43392 17020
rect 47670 16980 47676 16992
rect 31726 16952 43392 16980
rect 47631 16952 47676 16980
rect 47670 16940 47676 16952
rect 47728 16940 47734 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 17957 16779 18015 16785
rect 17957 16745 17969 16779
rect 18003 16776 18015 16779
rect 18506 16776 18512 16788
rect 18003 16748 18512 16776
rect 18003 16745 18015 16748
rect 17957 16739 18015 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19797 16779 19855 16785
rect 19797 16776 19809 16779
rect 19484 16748 19809 16776
rect 19484 16736 19490 16748
rect 19797 16745 19809 16748
rect 19843 16745 19855 16779
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 19797 16739 19855 16745
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25038 16776 25044 16788
rect 24999 16748 25044 16776
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 25685 16779 25743 16785
rect 25685 16745 25697 16779
rect 25731 16776 25743 16779
rect 25774 16776 25780 16788
rect 25731 16748 25780 16776
rect 25731 16745 25743 16748
rect 25685 16739 25743 16745
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 28813 16779 28871 16785
rect 28813 16745 28825 16779
rect 28859 16776 28871 16779
rect 28994 16776 29000 16788
rect 28859 16748 29000 16776
rect 28859 16745 28871 16748
rect 28813 16739 28871 16745
rect 28994 16736 29000 16748
rect 29052 16736 29058 16788
rect 12986 16708 12992 16720
rect 11716 16680 12992 16708
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 11716 16649 11744 16680
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 20254 16708 20260 16720
rect 20088 16680 20260 16708
rect 20088 16652 20116 16680
rect 20254 16668 20260 16680
rect 20312 16668 20318 16720
rect 23658 16668 23664 16720
rect 23716 16708 23722 16720
rect 25869 16711 25927 16717
rect 25869 16708 25881 16711
rect 23716 16680 25881 16708
rect 23716 16668 23722 16680
rect 25869 16677 25881 16680
rect 25915 16677 25927 16711
rect 25869 16671 25927 16677
rect 27617 16711 27675 16717
rect 27617 16677 27629 16711
rect 27663 16708 27675 16711
rect 29086 16708 29092 16720
rect 27663 16680 29092 16708
rect 27663 16677 27675 16680
rect 27617 16671 27675 16677
rect 29086 16668 29092 16680
rect 29144 16668 29150 16720
rect 29196 16680 31754 16708
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16609 11759 16643
rect 11882 16640 11888 16652
rect 11843 16612 11888 16640
rect 11701 16603 11759 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 16666 16640 16672 16652
rect 12492 16612 12537 16640
rect 14108 16612 16672 16640
rect 12492 16600 12498 16612
rect 14108 16581 14136 16612
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 17678 16600 17684 16652
rect 17736 16640 17742 16652
rect 19521 16643 19579 16649
rect 17736 16612 17908 16640
rect 17736 16600 17742 16612
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14182 16532 14188 16584
rect 14240 16572 14246 16584
rect 16206 16572 16212 16584
rect 14240 16544 14285 16572
rect 16167 16544 16212 16572
rect 14240 16532 14246 16544
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 17880 16581 17908 16612
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 20070 16640 20076 16652
rect 19567 16612 20076 16640
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 20346 16640 20352 16652
rect 20272 16612 20352 16640
rect 20272 16581 20300 16612
rect 20346 16600 20352 16612
rect 20404 16640 20410 16652
rect 21177 16643 21235 16649
rect 21177 16640 21189 16643
rect 20404 16612 21189 16640
rect 20404 16600 20410 16612
rect 21177 16609 21189 16612
rect 21223 16609 21235 16643
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 21177 16603 21235 16609
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 24394 16640 24400 16652
rect 23768 16612 24400 16640
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16572 20591 16575
rect 20714 16572 20720 16584
rect 20579 16544 20720 16572
rect 20579 16541 20591 16544
rect 20533 16535 20591 16541
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 19444 16504 19472 16535
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16574 23719 16575
rect 23768 16574 23796 16612
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 27522 16600 27528 16652
rect 27580 16640 27586 16652
rect 27580 16612 27660 16640
rect 27580 16600 27586 16612
rect 23707 16546 23796 16574
rect 23707 16541 23719 16546
rect 23661 16535 23719 16541
rect 24854 16532 24860 16584
rect 24912 16572 24918 16584
rect 24912 16544 25544 16572
rect 24912 16532 24918 16544
rect 20990 16504 20996 16516
rect 19444 16476 20996 16504
rect 20990 16464 20996 16476
rect 21048 16464 21054 16516
rect 23017 16507 23075 16513
rect 23017 16473 23029 16507
rect 23063 16504 23075 16507
rect 23382 16504 23388 16516
rect 23063 16476 23388 16504
rect 23063 16473 23075 16476
rect 23017 16467 23075 16473
rect 23382 16464 23388 16476
rect 23440 16464 23446 16516
rect 23566 16464 23572 16516
rect 23624 16504 23630 16516
rect 25516 16513 25544 16544
rect 25590 16532 25596 16584
rect 25648 16572 25654 16584
rect 25774 16572 25780 16584
rect 25648 16544 25780 16572
rect 25648 16532 25654 16544
rect 25774 16532 25780 16544
rect 25832 16532 25838 16584
rect 27632 16581 27660 16612
rect 27706 16600 27712 16652
rect 27764 16640 27770 16652
rect 27764 16612 27844 16640
rect 27764 16600 27770 16612
rect 27816 16581 27844 16612
rect 27890 16600 27896 16652
rect 27948 16640 27954 16652
rect 29196 16640 29224 16680
rect 30650 16640 30656 16652
rect 27948 16612 29224 16640
rect 30611 16612 30656 16640
rect 27948 16600 27954 16612
rect 30650 16600 30656 16612
rect 30708 16600 30714 16652
rect 31726 16640 31754 16680
rect 44082 16668 44088 16720
rect 44140 16708 44146 16720
rect 46566 16708 46572 16720
rect 44140 16680 46572 16708
rect 44140 16668 44146 16680
rect 32309 16643 32367 16649
rect 32309 16640 32321 16643
rect 31726 16612 32321 16640
rect 32309 16609 32321 16612
rect 32355 16609 32367 16643
rect 32309 16603 32367 16609
rect 27617 16575 27675 16581
rect 27617 16541 27629 16575
rect 27663 16541 27675 16575
rect 27617 16535 27675 16541
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 28350 16532 28356 16584
rect 28408 16572 28414 16584
rect 29638 16572 29644 16584
rect 28408 16544 28672 16572
rect 29599 16544 29644 16572
rect 28408 16532 28414 16544
rect 28644 16516 28672 16544
rect 29638 16532 29644 16544
rect 29696 16532 29702 16584
rect 29822 16572 29828 16584
rect 29783 16544 29828 16572
rect 29822 16532 29828 16544
rect 29880 16532 29886 16584
rect 45572 16581 45600 16680
rect 46566 16668 46572 16680
rect 46624 16668 46630 16720
rect 45646 16600 45652 16652
rect 45704 16640 45710 16652
rect 46293 16643 46351 16649
rect 45704 16612 45784 16640
rect 45704 16600 45710 16612
rect 45756 16581 45784 16612
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47762 16640 47768 16652
rect 46339 16612 47768 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47762 16600 47768 16612
rect 47820 16600 47826 16652
rect 48130 16640 48136 16652
rect 48091 16612 48136 16640
rect 48130 16600 48136 16612
rect 48188 16600 48194 16652
rect 45557 16575 45615 16581
rect 45557 16541 45569 16575
rect 45603 16541 45615 16575
rect 45557 16535 45615 16541
rect 45741 16575 45799 16581
rect 45741 16541 45753 16575
rect 45787 16541 45799 16575
rect 45741 16535 45799 16541
rect 24673 16507 24731 16513
rect 24673 16504 24685 16507
rect 23624 16476 24685 16504
rect 23624 16464 23630 16476
rect 24673 16473 24685 16476
rect 24719 16473 24731 16507
rect 24673 16467 24731 16473
rect 25501 16507 25559 16513
rect 25501 16473 25513 16507
rect 25547 16504 25559 16507
rect 25866 16504 25872 16516
rect 25547 16476 25872 16504
rect 25547 16473 25559 16476
rect 25501 16467 25559 16473
rect 25866 16464 25872 16476
rect 25924 16464 25930 16516
rect 28445 16507 28503 16513
rect 28445 16473 28457 16507
rect 28491 16504 28503 16507
rect 28534 16504 28540 16516
rect 28491 16476 28540 16504
rect 28491 16473 28503 16476
rect 28445 16467 28503 16473
rect 28534 16464 28540 16476
rect 28592 16464 28598 16516
rect 28626 16464 28632 16516
rect 28684 16504 28690 16516
rect 32490 16504 32496 16516
rect 28684 16476 28729 16504
rect 32451 16476 32496 16504
rect 28684 16464 28690 16476
rect 32490 16464 32496 16476
rect 32548 16464 32554 16516
rect 34149 16507 34207 16513
rect 34149 16473 34161 16507
rect 34195 16504 34207 16507
rect 42794 16504 42800 16516
rect 34195 16476 42800 16504
rect 34195 16473 34207 16476
rect 34149 16467 34207 16473
rect 42794 16464 42800 16476
rect 42852 16464 42858 16516
rect 45370 16464 45376 16516
rect 45428 16504 45434 16516
rect 45649 16507 45707 16513
rect 45649 16504 45661 16507
rect 45428 16476 45661 16504
rect 45428 16464 45434 16476
rect 45649 16473 45661 16476
rect 45695 16473 45707 16507
rect 45649 16467 45707 16473
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 16298 16436 16304 16448
rect 16259 16408 16304 16436
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 20070 16396 20076 16448
rect 20128 16436 20134 16448
rect 20355 16439 20413 16445
rect 20355 16436 20367 16439
rect 20128 16408 20367 16436
rect 20128 16396 20134 16408
rect 20355 16405 20367 16408
rect 20401 16405 20413 16439
rect 20355 16399 20413 16405
rect 20441 16439 20499 16445
rect 20441 16405 20453 16439
rect 20487 16436 20499 16439
rect 20898 16436 20904 16448
rect 20487 16408 20904 16436
rect 20487 16405 20499 16408
rect 20441 16399 20499 16405
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 23753 16439 23811 16445
rect 23753 16405 23765 16439
rect 23799 16436 23811 16439
rect 23842 16436 23848 16448
rect 23799 16408 23848 16436
rect 23799 16405 23811 16408
rect 23753 16399 23811 16405
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 24883 16439 24941 16445
rect 24883 16405 24895 16439
rect 24929 16436 24941 16439
rect 25590 16436 25596 16448
rect 24929 16408 25596 16436
rect 24929 16405 24941 16408
rect 24883 16399 24941 16405
rect 25590 16396 25596 16408
rect 25648 16396 25654 16448
rect 25711 16439 25769 16445
rect 25711 16405 25723 16439
rect 25757 16436 25769 16439
rect 25958 16436 25964 16448
rect 25757 16408 25964 16436
rect 25757 16405 25769 16408
rect 25711 16399 25769 16405
rect 25958 16396 25964 16408
rect 26016 16396 26022 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 19978 16232 19984 16244
rect 19939 16204 19984 16232
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 22738 16232 22744 16244
rect 20364 16204 22744 16232
rect 16025 16167 16083 16173
rect 16025 16133 16037 16167
rect 16071 16164 16083 16167
rect 16853 16167 16911 16173
rect 16853 16164 16865 16167
rect 16071 16136 16865 16164
rect 16071 16133 16083 16136
rect 16025 16127 16083 16133
rect 16853 16133 16865 16136
rect 16899 16133 16911 16167
rect 16853 16127 16911 16133
rect 19337 16167 19395 16173
rect 19337 16133 19349 16167
rect 19383 16164 19395 16167
rect 20162 16164 20168 16176
rect 19383 16136 20168 16164
rect 19383 16133 19395 16136
rect 19337 16127 19395 16133
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16096 2102 16108
rect 15933 16099 15991 16105
rect 2096 16068 2774 16096
rect 2096 16056 2102 16068
rect 2746 15892 2774 16068
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16206 16096 16212 16108
rect 15979 16068 16212 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16096 19303 16099
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19291 16068 19901 16096
rect 19291 16065 19303 16068
rect 19245 16059 19303 16065
rect 19889 16065 19901 16068
rect 19935 16096 19947 16099
rect 20364 16096 20392 16204
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 23566 16232 23572 16244
rect 23527 16204 23572 16232
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 25866 16232 25872 16244
rect 25827 16204 25872 16232
rect 25866 16192 25872 16204
rect 25924 16192 25930 16244
rect 28629 16235 28687 16241
rect 28629 16201 28641 16235
rect 28675 16232 28687 16235
rect 28718 16232 28724 16244
rect 28675 16204 28724 16232
rect 28675 16201 28687 16204
rect 28629 16195 28687 16201
rect 28718 16192 28724 16204
rect 28776 16192 28782 16244
rect 29181 16235 29239 16241
rect 29181 16201 29193 16235
rect 29227 16232 29239 16235
rect 29638 16232 29644 16244
rect 29227 16204 29644 16232
rect 29227 16201 29239 16204
rect 29181 16195 29239 16201
rect 29638 16192 29644 16204
rect 29696 16192 29702 16244
rect 32401 16235 32459 16241
rect 32401 16201 32413 16235
rect 32447 16232 32459 16235
rect 32490 16232 32496 16244
rect 32447 16204 32496 16232
rect 32447 16201 32459 16204
rect 32401 16195 32459 16201
rect 32490 16192 32496 16204
rect 32548 16192 32554 16244
rect 22186 16164 22192 16176
rect 19935 16068 20392 16096
rect 20456 16136 22192 16164
rect 19935 16065 19947 16068
rect 19889 16059 19947 16065
rect 16669 16031 16727 16037
rect 16669 15997 16681 16031
rect 16715 15997 16727 16031
rect 18506 16028 18512 16040
rect 18467 16000 18512 16028
rect 16669 15991 16727 15997
rect 16684 15960 16712 15991
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 20456 15960 20484 16136
rect 22186 16124 22192 16136
rect 22244 16124 22250 16176
rect 23106 16124 23112 16176
rect 23164 16124 23170 16176
rect 25958 16164 25964 16176
rect 25622 16136 25964 16164
rect 25958 16124 25964 16136
rect 26016 16124 26022 16176
rect 44266 16164 44272 16176
rect 44008 16136 44272 16164
rect 21174 16096 21180 16108
rect 21135 16068 21180 16096
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 26142 16056 26148 16108
rect 26200 16096 26206 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26200 16068 26985 16096
rect 26200 16056 26206 16068
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 28445 16099 28503 16105
rect 28445 16065 28457 16099
rect 28491 16096 28503 16099
rect 28534 16096 28540 16108
rect 28491 16068 28540 16096
rect 28491 16065 28503 16068
rect 28445 16059 28503 16065
rect 28534 16056 28540 16068
rect 28592 16056 28598 16108
rect 28626 16056 28632 16108
rect 28684 16096 28690 16108
rect 29086 16096 29092 16108
rect 28684 16068 28729 16096
rect 29047 16068 29092 16096
rect 28684 16056 28690 16068
rect 29086 16056 29092 16068
rect 29144 16056 29150 16108
rect 29273 16099 29331 16105
rect 29273 16065 29285 16099
rect 29319 16096 29331 16099
rect 30374 16096 30380 16108
rect 29319 16068 30380 16096
rect 29319 16065 29331 16068
rect 29273 16059 29331 16065
rect 30374 16056 30380 16068
rect 30432 16056 30438 16108
rect 31389 16099 31447 16105
rect 31389 16065 31401 16099
rect 31435 16096 31447 16099
rect 32309 16099 32367 16105
rect 32309 16096 32321 16099
rect 31435 16068 32321 16096
rect 31435 16065 31447 16068
rect 31389 16059 31447 16065
rect 32309 16065 32321 16068
rect 32355 16096 32367 16099
rect 32766 16096 32772 16108
rect 32355 16068 32772 16096
rect 32355 16065 32367 16068
rect 32309 16059 32367 16065
rect 32766 16056 32772 16068
rect 32824 16056 32830 16108
rect 44008 16105 44036 16136
rect 44266 16124 44272 16136
rect 44324 16124 44330 16176
rect 43993 16099 44051 16105
rect 43993 16065 44005 16099
rect 44039 16065 44051 16099
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 43993 16059 44051 16065
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 21269 16031 21327 16037
rect 21269 15997 21281 16031
rect 21315 16028 21327 16031
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21315 16000 21833 16028
rect 21315 15997 21327 16000
rect 21269 15991 21327 15997
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 24118 16028 24124 16040
rect 22152 16000 22197 16028
rect 24079 16000 24124 16028
rect 22152 15988 22158 16000
rect 24118 15988 24124 16000
rect 24176 15988 24182 16040
rect 24397 16031 24455 16037
rect 24397 15997 24409 16031
rect 24443 16028 24455 16031
rect 24854 16028 24860 16040
rect 24443 16000 24860 16028
rect 24443 15997 24455 16000
rect 24397 15991 24455 15997
rect 24854 15988 24860 16000
rect 24912 15988 24918 16040
rect 44174 16028 44180 16040
rect 44135 16000 44180 16028
rect 44174 15988 44180 16000
rect 44232 15988 44238 16040
rect 45830 16028 45836 16040
rect 45791 16000 45836 16028
rect 45830 15988 45836 16000
rect 45888 15988 45894 16040
rect 16684 15932 20484 15960
rect 21266 15892 21272 15904
rect 2746 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 26786 15892 26792 15904
rect 22244 15864 26792 15892
rect 22244 15852 22250 15864
rect 26786 15852 26792 15864
rect 26844 15852 26850 15904
rect 27065 15895 27123 15901
rect 27065 15861 27077 15895
rect 27111 15892 27123 15895
rect 27154 15892 27160 15904
rect 27111 15864 27160 15892
rect 27111 15861 27123 15864
rect 27065 15855 27123 15861
rect 27154 15852 27160 15864
rect 27212 15852 27218 15904
rect 30558 15852 30564 15904
rect 30616 15892 30622 15904
rect 31481 15895 31539 15901
rect 31481 15892 31493 15895
rect 30616 15864 31493 15892
rect 30616 15852 30622 15864
rect 31481 15861 31493 15864
rect 31527 15861 31539 15895
rect 31481 15855 31539 15861
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19613 15691 19671 15697
rect 19613 15688 19625 15691
rect 19392 15660 19625 15688
rect 19392 15648 19398 15660
rect 19613 15657 19625 15660
rect 19659 15657 19671 15691
rect 19613 15651 19671 15657
rect 21821 15691 21879 15697
rect 21821 15657 21833 15691
rect 21867 15688 21879 15691
rect 22094 15688 22100 15700
rect 21867 15660 22100 15688
rect 21867 15657 21879 15660
rect 21821 15651 21879 15657
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 23017 15691 23075 15697
rect 23017 15657 23029 15691
rect 23063 15688 23075 15691
rect 23106 15688 23112 15700
rect 23063 15660 23112 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 24854 15688 24860 15700
rect 23440 15660 23704 15688
rect 24815 15660 24860 15688
rect 23440 15648 23446 15660
rect 3510 15580 3516 15632
rect 3568 15620 3574 15632
rect 3568 15592 16620 15620
rect 3568 15580 3574 15592
rect 16298 15552 16304 15564
rect 16259 15524 16304 15552
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 16592 15561 16620 15592
rect 19076 15592 22094 15620
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15521 16635 15555
rect 16577 15515 16635 15521
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 16132 15416 16160 15447
rect 19076 15416 19104 15592
rect 20070 15552 20076 15564
rect 19628 15524 20076 15552
rect 19628 15493 19656 15524
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 22066 15552 22094 15592
rect 23566 15580 23572 15632
rect 23624 15580 23630 15632
rect 23676 15620 23704 15660
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 44085 15691 44143 15697
rect 26528 15660 31754 15688
rect 26528 15620 26556 15660
rect 23676 15592 26556 15620
rect 31726 15620 31754 15660
rect 44085 15657 44097 15691
rect 44131 15688 44143 15691
rect 44174 15688 44180 15700
rect 44131 15660 44180 15688
rect 44131 15657 44143 15660
rect 44085 15651 44143 15657
rect 44174 15648 44180 15660
rect 44232 15648 44238 15700
rect 45554 15620 45560 15632
rect 31726 15592 45560 15620
rect 45554 15580 45560 15592
rect 45612 15580 45618 15632
rect 23584 15552 23612 15580
rect 22066 15524 23612 15552
rect 23845 15555 23903 15561
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 20254 15484 20260 15496
rect 19843 15456 20260 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 22480 15493 22508 15524
rect 23845 15521 23857 15555
rect 23891 15552 23903 15555
rect 24118 15552 24124 15564
rect 23891 15524 24124 15552
rect 23891 15521 23903 15524
rect 23845 15515 23903 15521
rect 24118 15512 24124 15524
rect 24176 15512 24182 15564
rect 24670 15552 24676 15564
rect 24631 15524 24676 15552
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 25501 15555 25559 15561
rect 25501 15521 25513 15555
rect 25547 15521 25559 15555
rect 25501 15515 25559 15521
rect 25961 15555 26019 15561
rect 25961 15521 25973 15555
rect 26007 15552 26019 15555
rect 26697 15555 26755 15561
rect 26697 15552 26709 15555
rect 26007 15524 26709 15552
rect 26007 15521 26019 15524
rect 25961 15515 26019 15521
rect 26697 15521 26709 15524
rect 26743 15521 26755 15555
rect 26697 15515 26755 15521
rect 28169 15555 28227 15561
rect 28169 15521 28181 15555
rect 28215 15552 28227 15555
rect 30377 15555 30435 15561
rect 30377 15552 30389 15555
rect 28215 15524 30389 15552
rect 28215 15521 28227 15524
rect 28169 15515 28227 15521
rect 30377 15521 30389 15524
rect 30423 15521 30435 15555
rect 30558 15552 30564 15564
rect 30519 15524 30564 15552
rect 30377 15515 30435 15521
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 20772 15456 22017 15484
rect 20772 15444 20778 15456
rect 22005 15453 22017 15456
rect 22051 15453 22063 15487
rect 22005 15447 22063 15453
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 22465 15487 22523 15493
rect 22465 15453 22477 15487
rect 22511 15453 22523 15487
rect 22465 15447 22523 15453
rect 16132 15388 19104 15416
rect 22296 15416 22324 15447
rect 22738 15444 22744 15496
rect 22796 15484 22802 15496
rect 22925 15487 22983 15493
rect 22925 15484 22937 15487
rect 22796 15456 22937 15484
rect 22796 15444 22802 15456
rect 22925 15453 22937 15456
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 23658 15416 23664 15428
rect 22296 15388 23664 15416
rect 23658 15376 23664 15388
rect 23716 15376 23722 15428
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 23768 15348 23796 15447
rect 23934 15444 23940 15496
rect 23992 15484 23998 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 23992 15456 24593 15484
rect 23992 15444 23998 15456
rect 24581 15453 24593 15456
rect 24627 15484 24639 15487
rect 24762 15484 24768 15496
rect 24627 15456 24768 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 25222 15376 25228 15428
rect 25280 15416 25286 15428
rect 25516 15416 25544 15515
rect 25593 15487 25651 15493
rect 25593 15453 25605 15487
rect 25639 15484 25651 15487
rect 25774 15484 25780 15496
rect 25639 15456 25780 15484
rect 25639 15453 25651 15456
rect 25593 15447 25651 15453
rect 25774 15444 25780 15456
rect 25832 15484 25838 15496
rect 26421 15487 26479 15493
rect 25832 15456 26372 15484
rect 25832 15444 25838 15456
rect 26050 15416 26056 15428
rect 25280 15388 26056 15416
rect 25280 15376 25286 15388
rect 26050 15376 26056 15388
rect 26108 15376 26114 15428
rect 25682 15348 25688 15360
rect 21232 15320 25688 15348
rect 21232 15308 21238 15320
rect 25682 15308 25688 15320
rect 25740 15308 25746 15360
rect 26344 15348 26372 15456
rect 26421 15453 26433 15487
rect 26467 15453 26479 15487
rect 26421 15447 26479 15453
rect 26436 15416 26464 15447
rect 26602 15416 26608 15428
rect 26436 15388 26608 15416
rect 26602 15376 26608 15388
rect 26660 15376 26666 15428
rect 27154 15376 27160 15428
rect 27212 15376 27218 15428
rect 28184 15348 28212 15515
rect 30558 15512 30564 15524
rect 30616 15512 30622 15564
rect 30650 15512 30656 15564
rect 30708 15552 30714 15564
rect 30837 15555 30895 15561
rect 30837 15552 30849 15555
rect 30708 15524 30849 15552
rect 30708 15512 30714 15524
rect 30837 15521 30849 15524
rect 30883 15521 30895 15555
rect 30837 15515 30895 15521
rect 43806 15444 43812 15496
rect 43864 15484 43870 15496
rect 43990 15484 43996 15496
rect 43864 15456 43996 15484
rect 43864 15444 43870 15456
rect 43990 15444 43996 15456
rect 44048 15444 44054 15496
rect 26344 15320 28212 15348
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 25958 15144 25964 15156
rect 25919 15116 25964 15144
rect 25958 15104 25964 15116
rect 26016 15104 26022 15156
rect 26602 15104 26608 15156
rect 26660 15144 26666 15156
rect 27157 15147 27215 15153
rect 27157 15144 27169 15147
rect 26660 15116 27169 15144
rect 26660 15104 26666 15116
rect 27157 15113 27169 15116
rect 27203 15113 27215 15147
rect 27157 15107 27215 15113
rect 23753 15079 23811 15085
rect 23753 15045 23765 15079
rect 23799 15076 23811 15079
rect 23842 15076 23848 15088
rect 23799 15048 23848 15076
rect 23799 15045 23811 15048
rect 23753 15039 23811 15045
rect 23842 15036 23848 15048
rect 23900 15036 23906 15088
rect 25682 15036 25688 15088
rect 25740 15076 25746 15088
rect 25740 15048 27016 15076
rect 25740 15036 25746 15048
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 25869 15011 25927 15017
rect 25869 14977 25881 15011
rect 25915 15008 25927 15011
rect 26142 15008 26148 15020
rect 25915 14980 26148 15008
rect 25915 14977 25927 14980
rect 25869 14971 25927 14977
rect 26142 14968 26148 14980
rect 26200 14968 26206 15020
rect 26988 15017 27016 15048
rect 26973 15011 27031 15017
rect 26973 14977 26985 15011
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 42518 14968 42524 15020
rect 42576 15008 42582 15020
rect 43625 15011 43683 15017
rect 43625 15008 43637 15011
rect 42576 14980 43637 15008
rect 42576 14968 42582 14980
rect 43625 14977 43637 14980
rect 43671 14977 43683 15011
rect 43625 14971 43683 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2314 14940 2320 14952
rect 1995 14912 2320 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 23569 14943 23627 14949
rect 2832 14912 2877 14940
rect 2832 14900 2838 14912
rect 23569 14909 23581 14943
rect 23615 14940 23627 14943
rect 23934 14940 23940 14952
rect 23615 14912 23940 14940
rect 23615 14909 23627 14912
rect 23569 14903 23627 14909
rect 23934 14900 23940 14912
rect 23992 14900 23998 14952
rect 24029 14943 24087 14949
rect 24029 14909 24041 14943
rect 24075 14909 24087 14943
rect 43806 14940 43812 14952
rect 43767 14912 43812 14940
rect 24029 14903 24087 14909
rect 14734 14832 14740 14884
rect 14792 14872 14798 14884
rect 24044 14872 24072 14903
rect 43806 14900 43812 14912
rect 43864 14900 43870 14952
rect 45094 14940 45100 14952
rect 45055 14912 45100 14940
rect 45094 14900 45100 14912
rect 45152 14900 45158 14952
rect 14792 14844 24072 14872
rect 14792 14832 14798 14844
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2314 14600 2320 14612
rect 2275 14572 2320 14600
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 24670 14560 24676 14612
rect 24728 14600 24734 14612
rect 24765 14603 24823 14609
rect 24765 14600 24777 14603
rect 24728 14572 24777 14600
rect 24728 14560 24734 14572
rect 24765 14569 24777 14572
rect 24811 14569 24823 14603
rect 43806 14600 43812 14612
rect 43767 14572 43812 14600
rect 24765 14563 24823 14569
rect 43806 14560 43812 14572
rect 43864 14560 43870 14612
rect 25222 14464 25228 14476
rect 24688 14436 25228 14464
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2682 14396 2688 14408
rect 2271 14368 2688 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 24688 14405 24716 14436
rect 25222 14424 25228 14436
rect 25280 14424 25286 14476
rect 24673 14399 24731 14405
rect 2740 14356 2774 14396
rect 24673 14365 24685 14399
rect 24719 14365 24731 14399
rect 24673 14359 24731 14365
rect 24857 14399 24915 14405
rect 24857 14365 24869 14399
rect 24903 14396 24915 14399
rect 25774 14396 25780 14408
rect 24903 14368 25780 14396
rect 24903 14365 24915 14368
rect 24857 14359 24915 14365
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 43717 14399 43775 14405
rect 43717 14365 43729 14399
rect 43763 14396 43775 14399
rect 43990 14396 43996 14408
rect 43763 14368 43996 14396
rect 43763 14365 43775 14368
rect 43717 14359 43775 14365
rect 43990 14356 43996 14368
rect 44048 14356 44054 14408
rect 2746 14328 2774 14356
rect 33870 14328 33876 14340
rect 2746 14300 33876 14328
rect 33870 14288 33876 14300
rect 33928 14288 33934 14340
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 43990 13880 43996 13932
rect 44048 13920 44054 13932
rect 47581 13923 47639 13929
rect 47581 13920 47593 13923
rect 44048 13892 47593 13920
rect 44048 13880 44054 13892
rect 47581 13889 47593 13892
rect 47627 13889 47639 13923
rect 47581 13883 47639 13889
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 15286 13784 15292 13796
rect 4028 13756 15292 13784
rect 4028 13744 4034 13756
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 47670 13716 47676 13728
rect 47631 13688 47676 13716
rect 47670 13676 47676 13688
rect 47728 13676 47734 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 46477 13379 46535 13385
rect 46477 13345 46489 13379
rect 46523 13376 46535 13379
rect 47670 13376 47676 13388
rect 46523 13348 47676 13376
rect 46523 13345 46535 13348
rect 46477 13339 46535 13345
rect 47670 13336 47676 13348
rect 47728 13336 47734 13388
rect 46290 13308 46296 13320
rect 46251 13280 46296 13308
rect 46290 13268 46296 13280
rect 46348 13268 46354 13320
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 46290 12792 46296 12844
rect 46348 12832 46354 12844
rect 47765 12835 47823 12841
rect 47765 12832 47777 12835
rect 46348 12804 47777 12832
rect 46348 12792 46354 12804
rect 47765 12801 47777 12804
rect 47811 12801 47823 12835
rect 47765 12795 47823 12801
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 29362 12628 29368 12640
rect 1627 12600 29368 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 29362 12588 29368 12600
rect 29420 12588 29426 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 47670 11132 47676 11144
rect 47631 11104 47676 11132
rect 47670 11092 47676 11104
rect 47728 11092 47734 11144
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 12434 10996 12440 11008
rect 4120 10968 12440 10996
rect 4120 10956 4126 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 27614 10684 27620 10736
rect 27672 10724 27678 10736
rect 27798 10724 27804 10736
rect 27672 10696 27804 10724
rect 27672 10684 27678 10696
rect 27798 10684 27804 10696
rect 27856 10684 27862 10736
rect 47486 10616 47492 10668
rect 47544 10656 47550 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 47544 10628 47593 10656
rect 47544 10616 47550 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 46474 10412 46480 10464
rect 46532 10452 46538 10464
rect 47673 10455 47731 10461
rect 47673 10452 47685 10455
rect 46532 10424 47685 10452
rect 46532 10412 46538 10424
rect 47673 10421 47685 10424
rect 47719 10421 47731 10455
rect 47673 10415 47731 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 47670 10180 47676 10192
rect 46308 10152 47676 10180
rect 24397 10115 24455 10121
rect 24397 10081 24409 10115
rect 24443 10112 24455 10115
rect 25498 10112 25504 10124
rect 24443 10084 25504 10112
rect 24443 10081 24455 10084
rect 24397 10075 24455 10081
rect 25498 10072 25504 10084
rect 25556 10072 25562 10124
rect 26142 10112 26148 10124
rect 26103 10084 26148 10112
rect 26142 10072 26148 10084
rect 26200 10072 26206 10124
rect 46308 10121 46336 10152
rect 47670 10140 47676 10152
rect 47728 10140 47734 10192
rect 46293 10115 46351 10121
rect 46293 10081 46305 10115
rect 46339 10081 46351 10115
rect 46474 10112 46480 10124
rect 46435 10084 46480 10112
rect 46293 10075 46351 10081
rect 46474 10072 46480 10084
rect 46532 10072 46538 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 24578 9976 24584 9988
rect 24539 9948 24584 9976
rect 24578 9936 24584 9948
rect 24636 9936 24642 9988
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 24578 9704 24584 9716
rect 24539 9676 24584 9704
rect 24578 9664 24584 9676
rect 24636 9664 24642 9716
rect 24394 9528 24400 9580
rect 24452 9568 24458 9580
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 24452 9540 24501 9568
rect 24452 9528 24458 9540
rect 24489 9537 24501 9540
rect 24535 9568 24547 9571
rect 38930 9568 38936 9580
rect 24535 9540 38936 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 38930 9528 38936 9540
rect 38988 9528 38994 9580
rect 47854 9568 47860 9580
rect 47815 9540 47860 9568
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 46658 9392 46664 9444
rect 46716 9432 46722 9444
rect 48041 9435 48099 9441
rect 48041 9432 48053 9435
rect 46716 9404 48053 9432
rect 46716 9392 46722 9404
rect 48041 9401 48053 9404
rect 48087 9401 48099 9435
rect 48041 9395 48099 9401
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47762 8888 47768 8900
rect 47723 8860 47768 8888
rect 47762 8848 47768 8860
rect 47820 8848 47826 8900
rect 27338 8780 27344 8832
rect 27396 8820 27402 8832
rect 47857 8823 47915 8829
rect 47857 8820 47869 8823
rect 27396 8792 47869 8820
rect 27396 8780 27402 8792
rect 47857 8789 47869 8792
rect 47903 8789 47915 8823
rect 47857 8783 47915 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 44818 8616 44824 8628
rect 44779 8588 44824 8616
rect 44818 8576 44824 8588
rect 44876 8576 44882 8628
rect 45189 8483 45247 8489
rect 45189 8449 45201 8483
rect 45235 8480 45247 8483
rect 45554 8480 45560 8492
rect 45235 8452 45560 8480
rect 45235 8449 45247 8452
rect 45189 8443 45247 8449
rect 45554 8440 45560 8452
rect 45612 8440 45618 8492
rect 44818 8236 44824 8288
rect 44876 8276 44882 8288
rect 45281 8279 45339 8285
rect 45281 8276 45293 8279
rect 44876 8248 45293 8276
rect 44876 8236 44882 8248
rect 45281 8245 45293 8248
rect 45327 8245 45339 8279
rect 45646 8276 45652 8288
rect 45607 8248 45652 8276
rect 45281 8239 45339 8245
rect 45646 8236 45652 8248
rect 45704 8236 45710 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 42794 8032 42800 8084
rect 42852 8072 42858 8084
rect 46842 8072 46848 8084
rect 42852 8044 46848 8072
rect 42852 8032 42858 8044
rect 46842 8032 46848 8044
rect 46900 8032 46906 8084
rect 46566 7936 46572 7948
rect 46527 7908 46572 7936
rect 46566 7896 46572 7908
rect 46624 7896 46630 7948
rect 45373 7871 45431 7877
rect 45373 7837 45385 7871
rect 45419 7868 45431 7871
rect 45646 7868 45652 7880
rect 45419 7840 45652 7868
rect 45419 7837 45431 7840
rect 45373 7831 45431 7837
rect 45646 7828 45652 7840
rect 45704 7828 45710 7880
rect 45922 7800 45928 7812
rect 45883 7772 45928 7800
rect 45922 7760 45928 7772
rect 45980 7760 45986 7812
rect 46017 7803 46075 7809
rect 46017 7769 46029 7803
rect 46063 7769 46075 7803
rect 46017 7763 46075 7769
rect 45189 7735 45247 7741
rect 45189 7701 45201 7735
rect 45235 7732 45247 7735
rect 46032 7732 46060 7763
rect 45235 7704 46060 7732
rect 45235 7701 45247 7704
rect 45189 7695 45247 7701
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 45922 7488 45928 7540
rect 45980 7528 45986 7540
rect 47949 7531 48007 7537
rect 47949 7528 47961 7531
rect 45980 7500 47961 7528
rect 45980 7488 45986 7500
rect 47949 7497 47961 7500
rect 47995 7497 48007 7531
rect 47949 7491 48007 7497
rect 45646 7460 45652 7472
rect 45607 7432 45652 7460
rect 45646 7420 45652 7432
rect 45704 7420 45710 7472
rect 46566 7460 46572 7472
rect 46527 7432 46572 7460
rect 46566 7420 46572 7432
rect 46624 7420 46630 7472
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 45554 7284 45560 7336
rect 45612 7324 45618 7336
rect 45612 7296 45657 7324
rect 45612 7284 45618 7296
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 18506 6848 18512 6860
rect 4120 6820 18512 6848
rect 4120 6808 4126 6820
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 42334 6848 42340 6860
rect 42295 6820 42340 6848
rect 42334 6808 42340 6820
rect 42392 6808 42398 6860
rect 47302 6848 47308 6860
rect 47263 6820 47308 6848
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 46014 6740 46020 6792
rect 46072 6780 46078 6792
rect 47581 6783 47639 6789
rect 47581 6780 47593 6783
rect 46072 6752 47593 6780
rect 46072 6740 46078 6752
rect 47581 6749 47593 6752
rect 47627 6749 47639 6783
rect 47581 6743 47639 6749
rect 41325 6715 41383 6721
rect 41325 6712 41337 6715
rect 40880 6684 41337 6712
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 40880 6653 40908 6684
rect 41325 6681 41337 6684
rect 41371 6681 41383 6715
rect 41325 6675 41383 6681
rect 41414 6672 41420 6724
rect 41472 6712 41478 6724
rect 41472 6684 41517 6712
rect 41472 6672 41478 6684
rect 40865 6647 40923 6653
rect 40865 6644 40877 6647
rect 4028 6616 40877 6644
rect 4028 6604 4034 6616
rect 40865 6613 40877 6616
rect 40911 6613 40923 6647
rect 40865 6607 40923 6613
rect 42610 6604 42616 6656
rect 42668 6644 42674 6656
rect 45554 6644 45560 6656
rect 42668 6616 45560 6644
rect 42668 6604 42674 6616
rect 45554 6604 45560 6616
rect 45612 6604 45618 6656
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 41233 6443 41291 6449
rect 41233 6409 41245 6443
rect 41279 6440 41291 6443
rect 41414 6440 41420 6452
rect 41279 6412 41420 6440
rect 41279 6409 41291 6412
rect 41233 6403 41291 6409
rect 41414 6400 41420 6412
rect 41472 6400 41478 6452
rect 43806 6400 43812 6452
rect 43864 6440 43870 6452
rect 48041 6443 48099 6449
rect 48041 6440 48053 6443
rect 43864 6412 48053 6440
rect 43864 6400 43870 6412
rect 48041 6409 48053 6412
rect 48087 6409 48099 6443
rect 48041 6403 48099 6409
rect 42613 6375 42671 6381
rect 42613 6341 42625 6375
rect 42659 6372 42671 6375
rect 44174 6372 44180 6384
rect 42659 6344 44180 6372
rect 42659 6341 42671 6344
rect 42613 6335 42671 6341
rect 44174 6332 44180 6344
rect 44232 6332 44238 6384
rect 41322 6264 41328 6316
rect 41380 6304 41386 6316
rect 41417 6307 41475 6313
rect 41417 6304 41429 6307
rect 41380 6276 41429 6304
rect 41380 6264 41386 6276
rect 41417 6273 41429 6276
rect 41463 6273 41475 6307
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 41417 6267 41475 6273
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 41598 6196 41604 6248
rect 41656 6236 41662 6248
rect 42521 6239 42579 6245
rect 42521 6236 42533 6239
rect 41656 6208 42533 6236
rect 41656 6196 41662 6208
rect 42521 6205 42533 6208
rect 42567 6236 42579 6239
rect 42610 6236 42616 6248
rect 42567 6208 42616 6236
rect 42567 6205 42579 6208
rect 42521 6199 42579 6205
rect 42610 6196 42616 6208
rect 42668 6196 42674 6248
rect 42797 6239 42855 6245
rect 42797 6205 42809 6239
rect 42843 6205 42855 6239
rect 42797 6199 42855 6205
rect 42334 6128 42340 6180
rect 42392 6168 42398 6180
rect 42812 6168 42840 6199
rect 42392 6140 42840 6168
rect 42392 6128 42398 6140
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 38470 5856 38476 5908
rect 38528 5896 38534 5908
rect 40957 5899 41015 5905
rect 40957 5896 40969 5899
rect 38528 5868 40969 5896
rect 38528 5856 38534 5868
rect 40957 5865 40969 5868
rect 41003 5865 41015 5899
rect 41322 5896 41328 5908
rect 41283 5868 41328 5896
rect 40957 5859 41015 5865
rect 41322 5856 41328 5868
rect 41380 5856 41386 5908
rect 40865 5695 40923 5701
rect 40865 5661 40877 5695
rect 40911 5692 40923 5695
rect 44174 5692 44180 5704
rect 40911 5664 44180 5692
rect 40911 5661 40923 5664
rect 40865 5655 40923 5661
rect 44174 5652 44180 5664
rect 44232 5652 44238 5704
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 38657 5355 38715 5361
rect 38657 5352 38669 5355
rect 37384 5324 38669 5352
rect 37384 5293 37412 5324
rect 38657 5321 38669 5324
rect 38703 5321 38715 5355
rect 38657 5315 38715 5321
rect 37369 5287 37427 5293
rect 37369 5284 37381 5287
rect 22066 5256 37381 5284
rect 6638 5108 6644 5160
rect 6696 5148 6702 5160
rect 22066 5148 22094 5256
rect 37369 5253 37381 5256
rect 37415 5253 37427 5287
rect 37369 5247 37427 5253
rect 37458 5244 37464 5296
rect 37516 5284 37522 5296
rect 37516 5256 37561 5284
rect 37516 5244 37522 5256
rect 39669 5219 39727 5225
rect 39669 5185 39681 5219
rect 39715 5216 39727 5219
rect 41322 5216 41328 5228
rect 39715 5188 41328 5216
rect 39715 5185 39727 5188
rect 39669 5179 39727 5185
rect 41322 5176 41328 5188
rect 41380 5176 41386 5228
rect 47762 5216 47768 5228
rect 47723 5188 47768 5216
rect 47762 5176 47768 5188
rect 47820 5176 47826 5228
rect 38378 5148 38384 5160
rect 6696 5120 22094 5148
rect 38339 5120 38384 5148
rect 6696 5108 6702 5120
rect 38378 5108 38384 5120
rect 38436 5108 38442 5160
rect 23474 5040 23480 5092
rect 23532 5080 23538 5092
rect 47949 5083 48007 5089
rect 47949 5080 47961 5083
rect 23532 5052 47961 5080
rect 23532 5040 23538 5052
rect 47949 5049 47961 5052
rect 47995 5049 48007 5083
rect 47949 5043 48007 5049
rect 39114 4972 39120 5024
rect 39172 5012 39178 5024
rect 39761 5015 39819 5021
rect 39761 5012 39773 5015
rect 39172 4984 39773 5012
rect 39172 4972 39178 4984
rect 39761 4981 39773 4984
rect 39807 4981 39819 5015
rect 39761 4975 39819 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 20438 4700 20444 4752
rect 20496 4740 20502 4752
rect 28626 4740 28632 4752
rect 20496 4712 28632 4740
rect 20496 4700 20502 4712
rect 28626 4700 28632 4712
rect 28684 4700 28690 4752
rect 45646 4700 45652 4752
rect 45704 4740 45710 4752
rect 45704 4712 47624 4740
rect 45704 4700 45710 4712
rect 31110 4672 31116 4684
rect 12406 4644 31116 4672
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7708 4576 7941 4604
rect 7708 4564 7714 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 12406 4604 12434 4644
rect 31110 4632 31116 4644
rect 31168 4632 31174 4684
rect 47486 4672 47492 4684
rect 46676 4644 47492 4672
rect 15654 4604 15660 4616
rect 8987 4576 12434 4604
rect 15615 4576 15660 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 15654 4564 15660 4576
rect 15712 4564 15718 4616
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 16666 4604 16672 4616
rect 16347 4576 16672 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 20254 4564 20260 4616
rect 20312 4604 20318 4616
rect 20441 4607 20499 4613
rect 20441 4604 20453 4607
rect 20312 4576 20453 4604
rect 20312 4564 20318 4576
rect 20441 4573 20453 4576
rect 20487 4573 20499 4607
rect 21082 4604 21088 4616
rect 21043 4576 21088 4604
rect 20441 4567 20499 4573
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 21177 4607 21235 4613
rect 21177 4573 21189 4607
rect 21223 4604 21235 4607
rect 21729 4607 21787 4613
rect 21729 4604 21741 4607
rect 21223 4576 21741 4604
rect 21223 4573 21235 4576
rect 21177 4567 21235 4573
rect 21729 4573 21741 4576
rect 21775 4573 21787 4607
rect 22462 4604 22468 4616
rect 22423 4576 22468 4604
rect 21729 4567 21787 4573
rect 22462 4564 22468 4576
rect 22520 4564 22526 4616
rect 39114 4604 39120 4616
rect 39075 4576 39120 4604
rect 39114 4564 39120 4576
rect 39172 4564 39178 4616
rect 46676 4613 46704 4644
rect 47486 4632 47492 4644
rect 47544 4632 47550 4684
rect 47596 4681 47624 4712
rect 47581 4675 47639 4681
rect 47581 4641 47593 4675
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 39209 4607 39267 4613
rect 39209 4573 39221 4607
rect 39255 4604 39267 4607
rect 39853 4607 39911 4613
rect 39853 4604 39865 4607
rect 39255 4576 39865 4604
rect 39255 4573 39267 4576
rect 39209 4567 39267 4573
rect 39853 4573 39865 4576
rect 39899 4573 39911 4607
rect 39853 4567 39911 4573
rect 46661 4607 46719 4613
rect 46661 4573 46673 4607
rect 46707 4573 46719 4607
rect 46661 4567 46719 4573
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47305 4607 47363 4613
rect 47305 4604 47317 4607
rect 46900 4576 47317 4604
rect 46900 4564 46906 4576
rect 47305 4573 47317 4576
rect 47351 4573 47363 4607
rect 47305 4567 47363 4573
rect 15749 4539 15807 4545
rect 15749 4505 15761 4539
rect 15795 4536 15807 4539
rect 16850 4536 16856 4548
rect 15795 4508 16856 4536
rect 15795 4505 15807 4508
rect 15749 4499 15807 4505
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 40034 4536 40040 4548
rect 39995 4508 40040 4536
rect 40034 4496 40040 4508
rect 40092 4496 40098 4548
rect 41690 4536 41696 4548
rect 41603 4508 41696 4536
rect 41690 4496 41696 4508
rect 41748 4536 41754 4548
rect 42242 4536 42248 4548
rect 41748 4508 42248 4536
rect 41748 4496 41754 4508
rect 42242 4496 42248 4508
rect 42300 4496 42306 4548
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8352 4440 9045 4468
rect 8352 4428 8358 4440
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 9033 4431 9091 4437
rect 16393 4471 16451 4477
rect 16393 4437 16405 4471
rect 16439 4468 16451 4471
rect 17310 4468 17316 4480
rect 16439 4440 17316 4468
rect 16439 4437 16451 4440
rect 16393 4431 16451 4437
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 20533 4471 20591 4477
rect 20533 4437 20545 4471
rect 20579 4468 20591 4471
rect 21726 4468 21732 4480
rect 20579 4440 21732 4468
rect 20579 4437 20591 4440
rect 20533 4431 20591 4437
rect 21726 4428 21732 4440
rect 21784 4428 21790 4480
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4468 21879 4471
rect 22278 4468 22284 4480
rect 21867 4440 22284 4468
rect 21867 4437 21879 4440
rect 21821 4431 21879 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 22557 4471 22615 4477
rect 22557 4437 22569 4471
rect 22603 4468 22615 4471
rect 22646 4468 22652 4480
rect 22603 4440 22652 4468
rect 22603 4437 22615 4440
rect 22557 4431 22615 4437
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 45738 4428 45744 4480
rect 45796 4468 45802 4480
rect 46753 4471 46811 4477
rect 46753 4468 46765 4471
rect 45796 4440 46765 4468
rect 45796 4428 45802 4440
rect 46753 4437 46765 4440
rect 46799 4437 46811 4471
rect 46753 4431 46811 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 21082 4224 21088 4276
rect 21140 4264 21146 4276
rect 21913 4267 21971 4273
rect 21913 4264 21925 4267
rect 21140 4236 21925 4264
rect 21140 4224 21146 4236
rect 21913 4233 21925 4236
rect 21959 4233 21971 4267
rect 21913 4227 21971 4233
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 22833 4267 22891 4273
rect 22833 4264 22845 4267
rect 22520 4236 22845 4264
rect 22520 4224 22526 4236
rect 22833 4233 22845 4236
rect 22879 4233 22891 4267
rect 22833 4227 22891 4233
rect 40034 4224 40040 4276
rect 40092 4264 40098 4276
rect 40589 4267 40647 4273
rect 40589 4264 40601 4267
rect 40092 4236 40601 4264
rect 40092 4224 40098 4236
rect 40589 4233 40601 4236
rect 40635 4233 40647 4267
rect 40589 4227 40647 4233
rect 16942 4196 16948 4208
rect 16684 4168 16948 4196
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 7650 4128 7656 4140
rect 7611 4100 7656 4128
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 12069 4131 12127 4137
rect 9048 4100 9260 4128
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 8294 4060 8300 4072
rect 7883 4032 8300 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 4062 3952 4068 4004
rect 4120 3992 4126 4004
rect 9048 3992 9076 4100
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 4120 3964 9076 3992
rect 4120 3952 4126 3964
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1636 3896 2145 3924
rect 1636 3884 1642 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2832 3896 2881 3924
rect 2832 3884 2838 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 2869 3887 2927 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 9140 3924 9168 4023
rect 9232 3992 9260 4100
rect 12069 4097 12081 4131
rect 12115 4128 12127 4131
rect 12115 4100 12434 4128
rect 12115 4097 12127 4100
rect 12069 4091 12127 4097
rect 12406 4060 12434 4100
rect 13630 4088 13636 4140
rect 13688 4128 13694 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13688 4100 13737 4128
rect 13688 4088 13694 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 14366 4128 14372 4140
rect 14327 4100 14372 4128
rect 13725 4091 13783 4097
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14976 4100 15025 4128
rect 14976 4088 14982 4100
rect 15013 4097 15025 4100
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 16684 4137 16712 4168
rect 16942 4156 16948 4168
rect 17000 4156 17006 4208
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17184 4168 17448 4196
rect 17184 4156 17190 4168
rect 15657 4131 15715 4137
rect 15657 4128 15669 4131
rect 15252 4100 15669 4128
rect 15252 4088 15258 4100
rect 15657 4097 15669 4100
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 16816 4100 17325 4128
rect 16816 4088 16822 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 17420 4128 17448 4168
rect 19150 4156 19156 4208
rect 19208 4196 19214 4208
rect 21450 4196 21456 4208
rect 19208 4168 21456 4196
rect 19208 4156 19214 4168
rect 21450 4156 21456 4168
rect 21508 4156 21514 4208
rect 27614 4196 27620 4208
rect 27575 4168 27620 4196
rect 27614 4156 27620 4168
rect 27672 4156 27678 4208
rect 37366 4196 37372 4208
rect 37327 4168 37372 4196
rect 37366 4156 37372 4168
rect 37424 4156 37430 4208
rect 37461 4199 37519 4205
rect 37461 4165 37473 4199
rect 37507 4196 37519 4199
rect 37550 4196 37556 4208
rect 37507 4168 37556 4196
rect 37507 4165 37519 4168
rect 37461 4159 37519 4165
rect 37550 4156 37556 4168
rect 37608 4156 37614 4208
rect 38378 4196 38384 4208
rect 38339 4168 38384 4196
rect 38378 4156 38384 4168
rect 38436 4156 38442 4208
rect 39761 4199 39819 4205
rect 39761 4165 39773 4199
rect 39807 4196 39819 4199
rect 40218 4196 40224 4208
rect 39807 4168 40224 4196
rect 39807 4165 39819 4168
rect 39761 4159 39819 4165
rect 40218 4156 40224 4168
rect 40276 4156 40282 4208
rect 46382 4156 46388 4208
rect 46440 4196 46446 4208
rect 46569 4199 46627 4205
rect 46569 4196 46581 4199
rect 46440 4168 46581 4196
rect 46440 4156 46446 4168
rect 46569 4165 46581 4168
rect 46615 4165 46627 4199
rect 46569 4159 46627 4165
rect 46750 4156 46756 4208
rect 46808 4196 46814 4208
rect 47765 4199 47823 4205
rect 47765 4196 47777 4199
rect 46808 4168 47777 4196
rect 46808 4156 46814 4168
rect 47765 4165 47777 4168
rect 47811 4165 47823 4199
rect 47765 4159 47823 4165
rect 17954 4128 17960 4140
rect 17420 4100 17540 4128
rect 17915 4100 17960 4128
rect 17313 4091 17371 4097
rect 17512 4060 17540 4100
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18598 4128 18604 4140
rect 18559 4100 18604 4128
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 19242 4128 19248 4140
rect 19203 4100 19248 4128
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 19392 4100 19901 4128
rect 19392 4088 19398 4100
rect 19889 4097 19901 4100
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 20806 4128 20812 4140
rect 20579 4100 20812 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 21821 4131 21879 4137
rect 21821 4097 21833 4131
rect 21867 4128 21879 4131
rect 21910 4128 21916 4140
rect 21867 4100 21916 4128
rect 21867 4097 21879 4100
rect 21821 4091 21879 4097
rect 21910 4088 21916 4100
rect 21968 4088 21974 4140
rect 22278 4088 22284 4140
rect 22336 4128 22342 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22336 4100 22753 4128
rect 22336 4088 22342 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 23569 4131 23627 4137
rect 23569 4097 23581 4131
rect 23615 4128 23627 4131
rect 25130 4128 25136 4140
rect 23615 4100 25136 4128
rect 23615 4097 23627 4100
rect 23569 4091 23627 4097
rect 25130 4088 25136 4100
rect 25188 4088 25194 4140
rect 25222 4088 25228 4140
rect 25280 4128 25286 4140
rect 31386 4128 31392 4140
rect 25280 4100 25452 4128
rect 25280 4088 25286 4100
rect 25314 4060 25320 4072
rect 12406 4032 17356 4060
rect 17512 4032 25320 4060
rect 17126 3992 17132 4004
rect 9232 3964 17132 3992
rect 17126 3952 17132 3964
rect 17184 3952 17190 4004
rect 17328 3992 17356 4032
rect 25314 4020 25320 4032
rect 25372 4020 25378 4072
rect 25424 4060 25452 4100
rect 28368 4100 31392 4128
rect 27525 4063 27583 4069
rect 27525 4060 27537 4063
rect 25424 4032 27537 4060
rect 27525 4029 27537 4032
rect 27571 4060 27583 4063
rect 28368 4060 28396 4100
rect 31386 4088 31392 4100
rect 31444 4088 31450 4140
rect 36722 4128 36728 4140
rect 36683 4100 36728 4128
rect 36722 4088 36728 4100
rect 36780 4088 36786 4140
rect 39114 4128 39120 4140
rect 39075 4100 39120 4128
rect 39114 4088 39120 4100
rect 39172 4088 39178 4140
rect 39850 4088 39856 4140
rect 39908 4128 39914 4140
rect 39945 4131 40003 4137
rect 39945 4128 39957 4131
rect 39908 4100 39957 4128
rect 39908 4088 39914 4100
rect 39945 4097 39957 4100
rect 39991 4097 40003 4131
rect 39945 4091 40003 4097
rect 40129 4131 40187 4137
rect 40129 4097 40141 4131
rect 40175 4128 40187 4131
rect 40773 4131 40831 4137
rect 40773 4128 40785 4131
rect 40175 4100 40785 4128
rect 40175 4097 40187 4100
rect 40129 4091 40187 4097
rect 40773 4097 40785 4100
rect 40819 4097 40831 4131
rect 40773 4091 40831 4097
rect 41233 4131 41291 4137
rect 41233 4097 41245 4131
rect 41279 4097 41291 4131
rect 41233 4091 41291 4097
rect 28534 4060 28540 4072
rect 27571 4032 28396 4060
rect 28495 4032 28540 4060
rect 27571 4029 27583 4032
rect 27525 4023 27583 4029
rect 28534 4020 28540 4032
rect 28592 4020 28598 4072
rect 38010 4060 38016 4072
rect 28644 4032 38016 4060
rect 28644 3992 28672 4032
rect 38010 4020 38016 4032
rect 38068 4020 38074 4072
rect 39209 4063 39267 4069
rect 39209 4029 39221 4063
rect 39255 4060 39267 4063
rect 41248 4060 41276 4091
rect 41322 4088 41328 4140
rect 41380 4128 41386 4140
rect 42426 4128 42432 4140
rect 41380 4100 41425 4128
rect 42387 4100 42432 4128
rect 41380 4088 41386 4100
rect 42426 4088 42432 4100
rect 42484 4088 42490 4140
rect 39255 4032 41276 4060
rect 39255 4029 39267 4032
rect 39209 4023 39267 4029
rect 47949 3995 48007 4001
rect 47949 3992 47961 3995
rect 17328 3964 25360 3992
rect 7156 3896 9168 3924
rect 7156 3884 7162 3896
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 10137 3927 10195 3933
rect 10137 3924 10149 3927
rect 9272 3896 10149 3924
rect 9272 3884 9278 3896
rect 10137 3893 10149 3896
rect 10183 3893 10195 3927
rect 10137 3887 10195 3893
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11756 3896 12173 3924
rect 11756 3884 11762 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 14274 3924 14280 3936
rect 13863 3896 14280 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14826 3924 14832 3936
rect 14507 3896 14832 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15102 3924 15108 3936
rect 15063 3896 15108 3924
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15528 3896 15761 3924
rect 15528 3884 15534 3896
rect 15749 3893 15761 3896
rect 15795 3893 15807 3927
rect 15749 3887 15807 3893
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 16761 3927 16819 3933
rect 16761 3924 16773 3927
rect 16632 3896 16773 3924
rect 16632 3884 16638 3896
rect 16761 3893 16773 3896
rect 16807 3893 16819 3927
rect 16761 3887 16819 3893
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17276 3896 17417 3924
rect 17276 3884 17282 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17405 3887 17463 3893
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17920 3896 18061 3924
rect 17920 3884 17926 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 18693 3927 18751 3933
rect 18693 3924 18705 3927
rect 18564 3896 18705 3924
rect 18564 3884 18570 3896
rect 18693 3893 18705 3896
rect 18739 3893 18751 3927
rect 18693 3887 18751 3893
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19337 3927 19395 3933
rect 19337 3924 19349 3927
rect 18840 3896 19349 3924
rect 18840 3884 18846 3896
rect 19337 3893 19349 3896
rect 19383 3893 19395 3927
rect 19337 3887 19395 3893
rect 19981 3927 20039 3933
rect 19981 3893 19993 3927
rect 20027 3924 20039 3927
rect 20530 3924 20536 3936
rect 20027 3896 20536 3924
rect 20027 3893 20039 3896
rect 19981 3887 20039 3893
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 20680 3896 20725 3924
rect 20680 3884 20686 3896
rect 20898 3884 20904 3936
rect 20956 3924 20962 3936
rect 22830 3924 22836 3936
rect 20956 3896 22836 3924
rect 20956 3884 20962 3896
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 22922 3884 22928 3936
rect 22980 3924 22986 3936
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 22980 3896 23673 3924
rect 22980 3884 22986 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 23661 3887 23719 3893
rect 23842 3884 23848 3936
rect 23900 3924 23906 3936
rect 25222 3924 25228 3936
rect 23900 3896 25228 3924
rect 23900 3884 23906 3896
rect 25222 3884 25228 3896
rect 25280 3884 25286 3936
rect 25332 3924 25360 3964
rect 25516 3964 28672 3992
rect 31726 3964 47961 3992
rect 25516 3924 25544 3964
rect 25332 3896 25544 3924
rect 26418 3884 26424 3936
rect 26476 3924 26482 3936
rect 31726 3924 31754 3964
rect 47949 3961 47961 3964
rect 47995 3961 48007 3995
rect 47949 3955 48007 3961
rect 26476 3896 31754 3924
rect 36541 3927 36599 3933
rect 26476 3884 26482 3896
rect 36541 3893 36553 3927
rect 36587 3924 36599 3927
rect 37458 3924 37464 3936
rect 36587 3896 37464 3924
rect 36587 3893 36599 3896
rect 36541 3887 36599 3893
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 37550 3884 37556 3936
rect 37608 3924 37614 3936
rect 41782 3924 41788 3936
rect 37608 3896 41788 3924
rect 37608 3884 37614 3896
rect 41782 3884 41788 3896
rect 41840 3884 41846 3936
rect 42521 3927 42579 3933
rect 42521 3893 42533 3927
rect 42567 3924 42579 3927
rect 42610 3924 42616 3936
rect 42567 3896 42616 3924
rect 42567 3893 42579 3896
rect 42521 3887 42579 3893
rect 42610 3884 42616 3896
rect 42668 3884 42674 3936
rect 46017 3927 46075 3933
rect 46017 3893 46029 3927
rect 46063 3924 46075 3927
rect 46290 3924 46296 3936
rect 46063 3896 46296 3924
rect 46063 3893 46075 3896
rect 46017 3887 46075 3893
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 46658 3924 46664 3936
rect 46619 3896 46664 3924
rect 46658 3884 46664 3896
rect 46716 3884 46722 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 8018 3680 8024 3732
rect 8076 3720 8082 3732
rect 17313 3723 17371 3729
rect 8076 3692 17264 3720
rect 8076 3680 8082 3692
rect 9306 3612 9312 3664
rect 9364 3652 9370 3664
rect 16482 3652 16488 3664
rect 9364 3624 16488 3652
rect 9364 3612 9370 3624
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 16669 3655 16727 3661
rect 16669 3621 16681 3655
rect 16715 3652 16727 3655
rect 16758 3652 16764 3664
rect 16715 3624 16764 3652
rect 16715 3621 16727 3624
rect 16669 3615 16727 3621
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 17236 3652 17264 3692
rect 17313 3689 17325 3723
rect 17359 3720 17371 3723
rect 17954 3720 17960 3732
rect 17359 3692 17960 3720
rect 17359 3689 17371 3692
rect 17313 3683 17371 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 19242 3720 19248 3732
rect 18647 3692 19248 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 20806 3720 20812 3732
rect 20767 3692 20812 3720
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21450 3680 21456 3732
rect 21508 3720 21514 3732
rect 27893 3723 27951 3729
rect 21508 3692 27752 3720
rect 21508 3680 21514 3692
rect 20070 3652 20076 3664
rect 17236 3624 20076 3652
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 27724 3652 27752 3692
rect 27893 3689 27905 3723
rect 27939 3720 27951 3723
rect 35526 3720 35532 3732
rect 27939 3692 35532 3720
rect 27939 3689 27951 3692
rect 27893 3683 27951 3689
rect 35526 3680 35532 3692
rect 35584 3680 35590 3732
rect 37366 3720 37372 3732
rect 35866 3692 37372 3720
rect 29086 3652 29092 3664
rect 27724 3624 29092 3652
rect 29086 3612 29092 3624
rect 29144 3612 29150 3664
rect 31386 3612 31392 3664
rect 31444 3652 31450 3664
rect 35866 3652 35894 3692
rect 37366 3680 37372 3692
rect 37424 3680 37430 3732
rect 38562 3680 38568 3732
rect 38620 3720 38626 3732
rect 42426 3720 42432 3732
rect 38620 3692 42432 3720
rect 38620 3680 38626 3692
rect 42426 3680 42432 3692
rect 42484 3680 42490 3732
rect 31444 3624 35894 3652
rect 31444 3612 31450 3624
rect 39298 3612 39304 3664
rect 39356 3652 39362 3664
rect 42334 3652 42340 3664
rect 39356 3624 42340 3652
rect 39356 3612 39362 3624
rect 42334 3612 42340 3624
rect 42392 3612 42398 3664
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 1912 3556 3985 3584
rect 1912 3544 1918 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 8938 3584 8944 3596
rect 3973 3547 4031 3553
rect 7392 3556 8944 3584
rect 2682 3516 2688 3528
rect 2643 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3516 6975 3519
rect 7282 3516 7288 3528
rect 6963 3488 7288 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7392 3525 7420 3556
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9214 3584 9220 3596
rect 9175 3556 9220 3584
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9456 3556 9689 3584
rect 9456 3544 9462 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 14274 3584 14280 3596
rect 14235 3556 14280 3584
rect 9677 3547 9735 3553
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14516 3556 14565 3584
rect 14516 3544 14522 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3584 18015 3587
rect 18598 3584 18604 3596
rect 18003 3556 18604 3584
rect 18003 3553 18015 3556
rect 17957 3547 18015 3553
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 20438 3584 20444 3596
rect 18708 3556 20444 3584
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 8018 3516 8024 3528
rect 7979 3488 8024 3516
rect 7377 3479 7435 3485
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11572 3488 11713 3516
rect 11572 3476 11578 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13587 3488 14105 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 16574 3516 16580 3528
rect 16535 3488 16580 3516
rect 14093 3479 14151 3485
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 17218 3516 17224 3528
rect 17179 3488 17224 3516
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18506 3516 18512 3528
rect 18467 3488 18512 3516
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1360 3420 1869 3448
rect 1360 3408 1366 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 1857 3411 1915 3417
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 9401 3451 9459 3457
rect 2271 3420 8248 3448
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2777 3383 2835 3389
rect 2777 3380 2789 3383
rect 2096 3352 2789 3380
rect 2096 3340 2102 3352
rect 2777 3349 2789 3352
rect 2823 3349 2835 3383
rect 7466 3380 7472 3392
rect 7427 3352 7472 3380
rect 2777 3343 2835 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 8110 3380 8116 3392
rect 8071 3352 8116 3380
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 8220 3380 8248 3420
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 10042 3448 10048 3460
rect 9447 3420 10048 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 14642 3408 14648 3460
rect 14700 3448 14706 3460
rect 18598 3448 18604 3460
rect 14700 3420 18604 3448
rect 14700 3408 14706 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 18708 3380 18736 3556
rect 20438 3544 20444 3556
rect 20496 3544 20502 3596
rect 22462 3544 22468 3596
rect 22520 3584 22526 3596
rect 22925 3587 22983 3593
rect 22925 3584 22937 3587
rect 22520 3556 22937 3584
rect 22520 3544 22526 3556
rect 22925 3553 22937 3556
rect 22971 3584 22983 3587
rect 23842 3584 23848 3596
rect 22971 3556 23848 3584
rect 22971 3553 22983 3556
rect 22925 3547 22983 3553
rect 23842 3544 23848 3556
rect 23900 3544 23906 3596
rect 27890 3544 27896 3596
rect 27948 3584 27954 3596
rect 27948 3556 32260 3584
rect 27948 3544 27954 3556
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 19444 3448 19472 3479
rect 19978 3476 19984 3528
rect 20036 3516 20042 3528
rect 20257 3519 20315 3525
rect 20257 3516 20269 3519
rect 20036 3488 20269 3516
rect 20036 3476 20042 3488
rect 20257 3485 20269 3488
rect 20303 3485 20315 3519
rect 20257 3479 20315 3485
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 20588 3488 20729 3516
rect 20588 3476 20594 3488
rect 20717 3485 20729 3488
rect 20763 3485 20775 3519
rect 20717 3479 20775 3485
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22646 3516 22652 3528
rect 22336 3488 22381 3516
rect 22607 3488 22652 3516
rect 22336 3476 22342 3488
rect 22646 3476 22652 3488
rect 22704 3476 22710 3528
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 22796 3488 23765 3516
rect 22796 3476 22802 3488
rect 23753 3485 23765 3488
rect 23799 3485 23811 3519
rect 24670 3516 24676 3528
rect 24631 3488 24676 3516
rect 23753 3479 23811 3485
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 25498 3516 25504 3528
rect 25459 3488 25504 3516
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 27614 3516 27620 3528
rect 27575 3488 27620 3516
rect 27614 3476 27620 3488
rect 27672 3476 27678 3528
rect 32232 3516 32260 3556
rect 32858 3544 32864 3596
rect 32916 3584 32922 3596
rect 33781 3587 33839 3593
rect 33781 3584 33793 3587
rect 32916 3556 33793 3584
rect 32916 3544 32922 3556
rect 33781 3553 33793 3556
rect 33827 3553 33839 3587
rect 33781 3547 33839 3553
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 46290 3584 46296 3596
rect 33928 3556 45554 3584
rect 46251 3556 46296 3584
rect 33928 3544 33934 3556
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 32232 3488 32965 3516
rect 32953 3485 32965 3488
rect 32999 3516 33011 3519
rect 37918 3516 37924 3528
rect 32999 3488 37924 3516
rect 32999 3485 33011 3488
rect 32953 3479 33011 3485
rect 37918 3476 37924 3488
rect 37976 3516 37982 3528
rect 38562 3516 38568 3528
rect 37976 3488 38568 3516
rect 37976 3476 37982 3488
rect 38562 3476 38568 3488
rect 38620 3476 38626 3528
rect 40402 3516 40408 3528
rect 40363 3488 40408 3516
rect 40402 3476 40408 3488
rect 40460 3476 40466 3528
rect 40862 3516 40868 3528
rect 40823 3488 40868 3516
rect 40862 3476 40868 3488
rect 40920 3476 40926 3528
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 43349 3519 43407 3525
rect 43349 3516 43361 3519
rect 42484 3488 43361 3516
rect 42484 3476 42490 3488
rect 43349 3485 43361 3488
rect 43395 3485 43407 3519
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 43349 3479 43407 3485
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45526 3516 45554 3556
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 45649 3519 45707 3525
rect 45649 3516 45661 3519
rect 45526 3488 45661 3516
rect 45649 3485 45661 3488
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 24762 3448 24768 3460
rect 19444 3420 22232 3448
rect 24723 3420 24768 3448
rect 8220 3352 18736 3380
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 19484 3352 19533 3380
rect 19484 3340 19490 3352
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 19521 3343 19579 3349
rect 20162 3340 20168 3392
rect 20220 3380 20226 3392
rect 20622 3380 20628 3392
rect 20220 3352 20628 3380
rect 20220 3340 20226 3352
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 22094 3380 22100 3392
rect 20772 3352 22100 3380
rect 20772 3340 20778 3352
rect 22094 3340 22100 3352
rect 22152 3340 22158 3392
rect 22204 3380 22232 3420
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 25038 3408 25044 3460
rect 25096 3448 25102 3460
rect 40770 3448 40776 3460
rect 25096 3420 40776 3448
rect 25096 3408 25102 3420
rect 40770 3408 40776 3420
rect 40828 3408 40834 3460
rect 41049 3451 41107 3457
rect 41049 3448 41061 3451
rect 40880 3420 41061 3448
rect 27890 3380 27896 3392
rect 22204 3352 27896 3380
rect 27890 3340 27896 3352
rect 27948 3340 27954 3392
rect 28077 3383 28135 3389
rect 28077 3349 28089 3383
rect 28123 3380 28135 3383
rect 29178 3380 29184 3392
rect 28123 3352 29184 3380
rect 28123 3349 28135 3352
rect 28077 3343 28135 3349
rect 29178 3340 29184 3352
rect 29236 3340 29242 3392
rect 33042 3380 33048 3392
rect 33003 3352 33048 3380
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 40221 3383 40279 3389
rect 40221 3349 40233 3383
rect 40267 3380 40279 3383
rect 40880 3380 40908 3420
rect 41049 3417 41061 3420
rect 41095 3417 41107 3451
rect 41049 3411 41107 3417
rect 42242 3408 42248 3460
rect 42300 3448 42306 3460
rect 42705 3451 42763 3457
rect 42705 3448 42717 3451
rect 42300 3420 42717 3448
rect 42300 3408 42306 3420
rect 42705 3417 42717 3420
rect 42751 3417 42763 3451
rect 42705 3411 42763 3417
rect 45741 3451 45799 3457
rect 45741 3417 45753 3451
rect 45787 3448 45799 3451
rect 46477 3451 46535 3457
rect 46477 3448 46489 3451
rect 45787 3420 46489 3448
rect 45787 3417 45799 3420
rect 45741 3411 45799 3417
rect 46477 3417 46489 3420
rect 46523 3417 46535 3451
rect 46477 3411 46535 3417
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 40267 3352 40908 3380
rect 40267 3349 40279 3352
rect 40221 3343 40279 3349
rect 41138 3340 41144 3392
rect 41196 3380 41202 3392
rect 45462 3380 45468 3392
rect 41196 3352 45468 3380
rect 41196 3340 41202 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 14642 3176 14648 3188
rect 3844 3148 8708 3176
rect 3844 3136 3850 3148
rect 2038 3108 2044 3120
rect 1999 3080 2044 3108
rect 2038 3068 2044 3080
rect 2096 3068 2102 3120
rect 7466 3108 7472 3120
rect 7427 3080 7472 3108
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2317 2975 2375 2981
rect 2317 2972 2329 2975
rect 716 2944 2329 2972
rect 716 2932 722 2944
rect 2317 2941 2329 2944
rect 2363 2941 2375 2975
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 2317 2935 2375 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 8680 2972 8708 3148
rect 9968 3148 14648 3176
rect 9968 3049 9996 3148
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 14918 3176 14924 3188
rect 14879 3148 14924 3176
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15565 3179 15623 3185
rect 15565 3145 15577 3179
rect 15611 3176 15623 3179
rect 15654 3176 15660 3188
rect 15611 3148 15660 3176
rect 15611 3145 15623 3148
rect 15565 3139 15623 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 16761 3179 16819 3185
rect 16761 3176 16773 3179
rect 16724 3148 16773 3176
rect 16724 3136 16730 3148
rect 16761 3145 16773 3148
rect 16807 3145 16819 3179
rect 16761 3139 16819 3145
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17000 3148 17417 3176
rect 17000 3136 17006 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 18877 3179 18935 3185
rect 18877 3145 18889 3179
rect 18923 3176 18935 3179
rect 19242 3176 19248 3188
rect 18923 3148 19248 3176
rect 18923 3145 18935 3148
rect 18877 3139 18935 3145
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 36722 3176 36728 3188
rect 19352 3148 21772 3176
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 11698 3108 11704 3120
rect 10100 3080 10145 3108
rect 11659 3080 11704 3108
rect 10100 3068 10106 3080
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 19352 3108 19380 3148
rect 14016 3080 19380 3108
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 9953 3003 10011 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 14016 3049 14044 3080
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19613 3111 19671 3117
rect 19613 3108 19625 3111
rect 19484 3080 19625 3108
rect 19484 3068 19490 3080
rect 19613 3077 19625 3080
rect 19659 3077 19671 3111
rect 19613 3071 19671 3077
rect 19702 3068 19708 3120
rect 19760 3108 19766 3120
rect 21744 3108 21772 3148
rect 21928 3148 35894 3176
rect 36683 3148 36728 3176
rect 21928 3108 21956 3148
rect 22922 3108 22928 3120
rect 19760 3080 20852 3108
rect 21744 3080 21956 3108
rect 22883 3080 22928 3108
rect 19760 3068 19766 3080
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3009 14059 3043
rect 14826 3040 14832 3052
rect 14787 3012 14832 3040
rect 14001 3003 14059 3009
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 15470 3040 15476 3052
rect 15431 3012 15476 3040
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 16850 3040 16856 3052
rect 16715 3012 16856 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17310 3040 17316 3052
rect 17271 3012 17316 3040
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 11882 2972 11888 2984
rect 8680 2944 11888 2972
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 12308 2944 12353 2972
rect 12308 2932 12314 2944
rect 12388 2932 12394 2984
rect 12446 2972 12452 2984
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 12446 2944 13921 2972
rect 12446 2932 12452 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 14366 2972 14372 2984
rect 14327 2944 14372 2972
rect 13909 2935 13967 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 16482 2932 16488 2984
rect 16540 2972 16546 2984
rect 19334 2972 19340 2984
rect 16540 2944 19340 2972
rect 16540 2932 16546 2944
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 19978 2972 19984 2984
rect 19475 2944 19984 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20346 2972 20352 2984
rect 20307 2944 20352 2972
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 20824 2972 20852 3080
rect 22922 3068 22928 3080
rect 22980 3068 22986 3120
rect 23014 3068 23020 3120
rect 23072 3108 23078 3120
rect 24394 3108 24400 3120
rect 23072 3080 24400 3108
rect 23072 3068 23078 3080
rect 24394 3068 24400 3080
rect 24452 3068 24458 3120
rect 25317 3111 25375 3117
rect 25317 3077 25329 3111
rect 25363 3108 25375 3111
rect 25406 3108 25412 3120
rect 25363 3080 25412 3108
rect 25363 3077 25375 3080
rect 25317 3071 25375 3077
rect 25406 3068 25412 3080
rect 25464 3068 25470 3120
rect 27525 3111 27583 3117
rect 27525 3108 27537 3111
rect 25516 3080 27537 3108
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21784 3012 21833 3040
rect 21784 3000 21790 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 22738 3040 22744 3052
rect 21968 3012 22013 3040
rect 22699 3012 22744 3040
rect 21968 3000 21974 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 24486 3000 24492 3052
rect 24544 3040 24550 3052
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 24544 3012 25145 3040
rect 24544 3000 24550 3012
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 23014 2972 23020 2984
rect 20824 2944 23020 2972
rect 23014 2932 23020 2944
rect 23072 2932 23078 2984
rect 23106 2932 23112 2984
rect 23164 2972 23170 2984
rect 23201 2975 23259 2981
rect 23201 2972 23213 2975
rect 23164 2944 23213 2972
rect 23164 2932 23170 2944
rect 23201 2941 23213 2944
rect 23247 2941 23259 2975
rect 23201 2935 23259 2941
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 25516 2972 25544 3080
rect 27525 3077 27537 3080
rect 27571 3077 27583 3111
rect 27525 3071 27583 3077
rect 27617 3111 27675 3117
rect 27617 3077 27629 3111
rect 27663 3108 27675 3111
rect 27890 3108 27896 3120
rect 27663 3080 27896 3108
rect 27663 3077 27675 3080
rect 27617 3071 27675 3077
rect 27890 3068 27896 3080
rect 27948 3068 27954 3120
rect 28534 3108 28540 3120
rect 28495 3080 28540 3108
rect 28534 3068 28540 3080
rect 28592 3068 28598 3120
rect 33042 3108 33048 3120
rect 33003 3080 33048 3108
rect 33042 3068 33048 3080
rect 33100 3068 33106 3120
rect 35866 3108 35894 3148
rect 36722 3136 36728 3148
rect 36780 3136 36786 3188
rect 39114 3136 39120 3188
rect 39172 3176 39178 3188
rect 39853 3179 39911 3185
rect 39853 3176 39865 3179
rect 39172 3148 39865 3176
rect 39172 3136 39178 3148
rect 39853 3145 39865 3148
rect 39899 3145 39911 3179
rect 39853 3139 39911 3145
rect 40034 3136 40040 3188
rect 40092 3176 40098 3188
rect 40678 3176 40684 3188
rect 40092 3148 40684 3176
rect 40092 3136 40098 3148
rect 40678 3136 40684 3148
rect 40736 3136 40742 3188
rect 40862 3136 40868 3188
rect 40920 3176 40926 3188
rect 41049 3179 41107 3185
rect 41049 3176 41061 3179
rect 40920 3148 41061 3176
rect 40920 3136 40926 3148
rect 41049 3145 41061 3148
rect 41095 3145 41107 3179
rect 48038 3176 48044 3188
rect 47999 3148 48044 3176
rect 41049 3139 41107 3145
rect 48038 3136 48044 3148
rect 48096 3136 48102 3188
rect 42242 3108 42248 3120
rect 35866 3080 42248 3108
rect 42242 3068 42248 3080
rect 42300 3068 42306 3120
rect 42610 3108 42616 3120
rect 42571 3080 42616 3108
rect 42610 3068 42616 3080
rect 42668 3068 42674 3120
rect 45373 3111 45431 3117
rect 45373 3077 45385 3111
rect 45419 3108 45431 3111
rect 45738 3108 45744 3120
rect 45419 3080 45744 3108
rect 45419 3077 45431 3080
rect 45373 3071 45431 3077
rect 45738 3068 45744 3080
rect 45796 3068 45802 3120
rect 29178 3040 29184 3052
rect 29139 3012 29184 3040
rect 29178 3000 29184 3012
rect 29236 3000 29242 3052
rect 32858 3040 32864 3052
rect 32819 3012 32864 3040
rect 32858 3000 32864 3012
rect 32916 3000 32922 3052
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3040 36323 3043
rect 37550 3040 37556 3052
rect 36311 3012 37556 3040
rect 36311 3009 36323 3012
rect 36265 3003 36323 3009
rect 37550 3000 37556 3012
rect 37608 3000 37614 3052
rect 39209 3043 39267 3049
rect 39209 3009 39221 3043
rect 39255 3040 39267 3043
rect 39255 3012 39988 3040
rect 39255 3009 39267 3012
rect 39209 3003 39267 3009
rect 23532 2944 25544 2972
rect 23532 2932 23538 2944
rect 25590 2932 25596 2984
rect 25648 2972 25654 2984
rect 32766 2972 32772 2984
rect 25648 2944 32772 2972
rect 25648 2932 25654 2944
rect 32766 2932 32772 2944
rect 32824 2932 32830 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 37366 2932 37372 2984
rect 37424 2972 37430 2984
rect 39224 2972 39252 3003
rect 37424 2944 39252 2972
rect 39393 2975 39451 2981
rect 37424 2932 37430 2944
rect 39393 2941 39405 2975
rect 39439 2972 39451 2975
rect 39850 2972 39856 2984
rect 39439 2944 39856 2972
rect 39439 2941 39451 2944
rect 39393 2935 39451 2941
rect 39850 2932 39856 2944
rect 39908 2932 39914 2984
rect 39960 2972 39988 3012
rect 40126 3000 40132 3052
rect 40184 3040 40190 3052
rect 41693 3043 41751 3049
rect 41693 3040 41705 3043
rect 40184 3012 41705 3040
rect 40184 3000 40190 3012
rect 41693 3009 41705 3012
rect 41739 3009 41751 3043
rect 42426 3040 42432 3052
rect 42387 3012 42432 3040
rect 41693 3003 41751 3009
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3040 47823 3043
rect 48314 3040 48320 3052
rect 47811 3012 48320 3040
rect 47811 3009 47823 3012
rect 47765 3003 47823 3009
rect 48314 3000 48320 3012
rect 48372 3000 48378 3052
rect 40405 2975 40463 2981
rect 40405 2972 40417 2975
rect 39960 2944 40417 2972
rect 40405 2941 40417 2944
rect 40451 2941 40463 2975
rect 40586 2972 40592 2984
rect 40547 2944 40592 2972
rect 40405 2935 40463 2941
rect 3878 2864 3884 2916
rect 3936 2904 3942 2916
rect 3936 2876 6960 2904
rect 3936 2864 3942 2876
rect 6822 2836 6828 2848
rect 6783 2808 6828 2836
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 6932 2836 6960 2876
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11974 2904 11980 2916
rect 11020 2876 11980 2904
rect 11020 2864 11026 2876
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 24118 2904 24124 2916
rect 12084 2876 24124 2904
rect 12084 2836 12112 2876
rect 24118 2864 24124 2876
rect 24176 2864 24182 2916
rect 27614 2864 27620 2916
rect 27672 2904 27678 2916
rect 40034 2904 40040 2916
rect 27672 2876 40040 2904
rect 27672 2864 27678 2876
rect 40034 2864 40040 2876
rect 40092 2864 40098 2916
rect 40420 2904 40448 2935
rect 40586 2932 40592 2944
rect 40644 2932 40650 2984
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 43162 2972 43168 2984
rect 40736 2944 41736 2972
rect 43123 2944 43168 2972
rect 40736 2932 40742 2944
rect 41598 2904 41604 2916
rect 40420 2876 41604 2904
rect 41598 2864 41604 2876
rect 41656 2864 41662 2916
rect 41708 2904 41736 2944
rect 43162 2932 43168 2944
rect 43220 2932 43226 2984
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 43898 2904 43904 2916
rect 41708 2876 43904 2904
rect 43898 2864 43904 2876
rect 43956 2864 43962 2916
rect 6932 2808 12112 2836
rect 12158 2796 12164 2848
rect 12216 2836 12222 2848
rect 19242 2836 19248 2848
rect 12216 2808 19248 2836
rect 12216 2796 12222 2808
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 27890 2796 27896 2848
rect 27948 2836 27954 2848
rect 28997 2839 29055 2845
rect 28997 2836 29009 2839
rect 27948 2808 29009 2836
rect 27948 2796 27954 2808
rect 28997 2805 29009 2808
rect 29043 2805 29055 2839
rect 28997 2799 29055 2805
rect 29086 2796 29092 2848
rect 29144 2836 29150 2848
rect 32214 2836 32220 2848
rect 29144 2808 32220 2836
rect 29144 2796 29150 2808
rect 32214 2796 32220 2808
rect 32272 2796 32278 2848
rect 36354 2836 36360 2848
rect 36315 2808 36360 2836
rect 36354 2796 36360 2808
rect 36412 2796 36418 2848
rect 39850 2796 39856 2848
rect 39908 2836 39914 2848
rect 41509 2839 41567 2845
rect 41509 2836 41521 2839
rect 39908 2808 41521 2836
rect 39908 2796 39914 2808
rect 41509 2805 41521 2808
rect 41555 2805 41567 2839
rect 41509 2799 41567 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 12342 2632 12348 2644
rect 5307 2604 12348 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14645 2635 14703 2641
rect 14645 2601 14657 2635
rect 14691 2632 14703 2635
rect 15194 2632 15200 2644
rect 14691 2604 15200 2632
rect 14691 2601 14703 2604
rect 14645 2595 14703 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 19889 2635 19947 2641
rect 16546 2604 19840 2632
rect 2774 2564 2780 2576
rect 1412 2536 2780 2564
rect 1412 2505 1440 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 6454 2524 6460 2576
rect 6512 2564 6518 2576
rect 16546 2564 16574 2604
rect 6512 2536 7052 2564
rect 6512 2524 6518 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2866 2496 2872 2508
rect 2827 2468 2872 2496
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 6822 2496 6828 2508
rect 6595 2468 6828 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7024 2505 7052 2536
rect 9600 2536 16574 2564
rect 17313 2567 17371 2573
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2792 2400 3801 2428
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2792 2360 2820 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 2648 2332 2820 2360
rect 2648 2320 2654 2332
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 6733 2363 6791 2369
rect 3292 2332 5396 2360
rect 3292 2320 3298 2332
rect 3970 2292 3976 2304
rect 3931 2264 3976 2292
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 5368 2292 5396 2332
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 8110 2360 8116 2372
rect 6779 2332 8116 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8444 2332 9413 2360
rect 8444 2320 8450 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 9600 2292 9628 2536
rect 17313 2533 17325 2567
rect 17359 2564 17371 2567
rect 17678 2564 17684 2576
rect 17359 2536 17684 2564
rect 17359 2533 17371 2536
rect 17313 2527 17371 2533
rect 17678 2524 17684 2536
rect 17736 2524 17742 2576
rect 19812 2564 19840 2604
rect 19889 2601 19901 2635
rect 19935 2632 19947 2635
rect 20438 2632 20444 2644
rect 19935 2604 20444 2632
rect 19935 2601 19947 2604
rect 19889 2595 19947 2601
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20680 2604 20913 2632
rect 20680 2592 20686 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 20901 2595 20959 2601
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 22373 2635 22431 2641
rect 22373 2632 22385 2635
rect 22336 2604 22385 2632
rect 22336 2592 22342 2604
rect 22373 2601 22385 2604
rect 22419 2601 22431 2635
rect 22373 2595 22431 2601
rect 23385 2635 23443 2641
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 23474 2632 23480 2644
rect 23431 2604 23480 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 24946 2592 24952 2644
rect 25004 2632 25010 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 25004 2604 28641 2632
rect 25004 2592 25010 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 35526 2632 35532 2644
rect 35487 2604 35532 2632
rect 28629 2595 28687 2601
rect 35526 2592 35532 2604
rect 35584 2592 35590 2644
rect 35618 2592 35624 2644
rect 35676 2632 35682 2644
rect 36357 2635 36415 2641
rect 36357 2632 36369 2635
rect 35676 2604 36369 2632
rect 35676 2592 35682 2604
rect 36357 2601 36369 2604
rect 36403 2601 36415 2635
rect 40218 2632 40224 2644
rect 40179 2604 40224 2632
rect 36357 2595 36415 2601
rect 40218 2592 40224 2604
rect 40276 2592 40282 2644
rect 40402 2592 40408 2644
rect 40460 2632 40466 2644
rect 40497 2635 40555 2641
rect 40497 2632 40509 2635
rect 40460 2604 40509 2632
rect 40460 2592 40466 2604
rect 40497 2601 40509 2604
rect 40543 2601 40555 2635
rect 40497 2595 40555 2601
rect 41141 2635 41199 2641
rect 41141 2601 41153 2635
rect 41187 2632 41199 2635
rect 42518 2632 42524 2644
rect 41187 2604 42524 2632
rect 41187 2601 41199 2604
rect 41141 2595 41199 2601
rect 42518 2592 42524 2604
rect 42576 2592 42582 2644
rect 25498 2564 25504 2576
rect 19812 2536 24164 2564
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2496 9735 2499
rect 24026 2496 24032 2508
rect 9723 2468 24032 2496
rect 9723 2465 9735 2468
rect 9677 2459 9735 2465
rect 24026 2456 24032 2468
rect 24084 2456 24090 2508
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2428 14611 2431
rect 15102 2428 15108 2440
rect 14599 2400 15108 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15470 2428 15476 2440
rect 15335 2400 15476 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 19797 2431 19855 2437
rect 15620 2400 15665 2428
rect 15620 2388 15626 2400
rect 19797 2397 19809 2431
rect 19843 2428 19855 2431
rect 20162 2428 20168 2440
rect 19843 2400 20168 2428
rect 19843 2397 19855 2400
rect 19797 2391 19855 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23256 2400 23581 2428
rect 23256 2388 23262 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16172 2332 17141 2360
rect 16172 2320 16178 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 21910 2320 21916 2372
rect 21968 2360 21974 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21968 2332 22293 2360
rect 21968 2320 21974 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 24136 2360 24164 2536
rect 24596 2536 25504 2564
rect 24596 2505 24624 2536
rect 25498 2524 25504 2536
rect 25556 2524 25562 2576
rect 27798 2524 27804 2576
rect 27856 2564 27862 2576
rect 30193 2567 30251 2573
rect 30193 2564 30205 2567
rect 27856 2536 30205 2564
rect 27856 2524 27862 2536
rect 30193 2533 30205 2536
rect 30239 2533 30251 2567
rect 30193 2527 30251 2533
rect 32122 2524 32128 2576
rect 32180 2564 32186 2576
rect 38289 2567 38347 2573
rect 38289 2564 38301 2567
rect 32180 2536 38301 2564
rect 32180 2524 32186 2536
rect 38289 2533 38301 2536
rect 38335 2533 38347 2567
rect 38289 2527 38347 2533
rect 41693 2567 41751 2573
rect 41693 2533 41705 2567
rect 41739 2533 41751 2567
rect 41693 2527 41751 2533
rect 24581 2499 24639 2505
rect 24581 2465 24593 2499
rect 24627 2465 24639 2499
rect 24762 2496 24768 2508
rect 24723 2468 24768 2496
rect 24581 2459 24639 2465
rect 24762 2456 24768 2468
rect 24820 2456 24826 2508
rect 25130 2496 25136 2508
rect 25091 2468 25136 2496
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 27249 2499 27307 2505
rect 27249 2465 27261 2499
rect 27295 2496 27307 2499
rect 27706 2496 27712 2508
rect 27295 2468 27712 2496
rect 27295 2465 27307 2468
rect 27249 2459 27307 2465
rect 27706 2456 27712 2468
rect 27764 2456 27770 2508
rect 32490 2456 32496 2508
rect 32548 2496 32554 2508
rect 39301 2499 39359 2505
rect 39301 2496 39313 2499
rect 32548 2468 39313 2496
rect 32548 2456 32554 2468
rect 39301 2465 39313 2468
rect 39347 2465 39359 2499
rect 39301 2459 39359 2465
rect 40221 2499 40279 2505
rect 40221 2465 40233 2499
rect 40267 2496 40279 2499
rect 40586 2496 40592 2508
rect 40267 2468 40592 2496
rect 40267 2465 40279 2468
rect 40221 2459 40279 2465
rect 40586 2456 40592 2468
rect 40644 2496 40650 2508
rect 41708 2496 41736 2527
rect 40644 2468 41736 2496
rect 40644 2456 40650 2468
rect 41782 2456 41788 2508
rect 41840 2496 41846 2508
rect 43901 2499 43959 2505
rect 43901 2496 43913 2499
rect 41840 2468 43913 2496
rect 41840 2456 41846 2468
rect 43901 2465 43913 2468
rect 43947 2465 43959 2499
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 43901 2459 43959 2465
rect 45526 2468 46489 2496
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 30837 2431 30895 2437
rect 30837 2428 30849 2431
rect 29696 2400 30849 2428
rect 29696 2388 29702 2400
rect 30837 2397 30849 2400
rect 30883 2397 30895 2431
rect 30837 2391 30895 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 38068 2400 38117 2428
rect 38068 2388 38074 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39850 2388 39856 2440
rect 39908 2428 39914 2440
rect 39945 2431 40003 2437
rect 39945 2428 39957 2431
rect 39908 2400 39957 2428
rect 39908 2388 39914 2400
rect 39945 2397 39957 2400
rect 39991 2397 40003 2431
rect 39945 2391 40003 2397
rect 41230 2388 41236 2440
rect 41288 2428 41294 2440
rect 41877 2431 41935 2437
rect 41877 2428 41889 2431
rect 41288 2400 41889 2428
rect 41288 2388 41294 2400
rect 41877 2397 41889 2400
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 44174 2388 44180 2440
rect 44232 2428 44238 2440
rect 45526 2428 45554 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 46477 2459 46535 2465
rect 46566 2456 46572 2508
rect 46624 2496 46630 2508
rect 47857 2499 47915 2505
rect 47857 2496 47869 2499
rect 46624 2468 47869 2496
rect 46624 2456 46630 2468
rect 47857 2465 47869 2468
rect 47903 2465 47915 2499
rect 47857 2459 47915 2465
rect 44232 2400 45554 2428
rect 46201 2431 46259 2437
rect 44232 2388 44238 2400
rect 46201 2397 46213 2431
rect 46247 2428 46259 2431
rect 47026 2428 47032 2440
rect 46247 2400 47032 2428
rect 46247 2397 46259 2400
rect 46201 2391 46259 2397
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 47673 2431 47731 2437
rect 47673 2397 47685 2431
rect 47719 2428 47731 2431
rect 48038 2428 48044 2440
rect 47719 2400 48044 2428
rect 47719 2397 47731 2400
rect 47673 2391 47731 2397
rect 48038 2388 48044 2400
rect 48096 2388 48102 2440
rect 26142 2360 26148 2372
rect 24136 2332 26148 2360
rect 22281 2323 22339 2329
rect 26142 2320 26148 2332
rect 26200 2320 26206 2372
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 30009 2363 30067 2369
rect 30009 2360 30021 2363
rect 27120 2332 30021 2360
rect 27120 2320 27126 2332
rect 30009 2329 30021 2332
rect 30055 2329 30067 2363
rect 30009 2323 30067 2329
rect 30668 2332 35894 2360
rect 30668 2301 30696 2332
rect 5368 2264 9628 2292
rect 30653 2295 30711 2301
rect 30653 2261 30665 2295
rect 30699 2261 30711 2295
rect 35866 2292 35894 2332
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 39117 2363 39175 2369
rect 39117 2329 39129 2363
rect 39163 2360 39175 2363
rect 39298 2360 39304 2372
rect 39163 2332 39304 2360
rect 39163 2329 39175 2332
rect 39117 2323 39175 2329
rect 39298 2320 39304 2332
rect 39356 2320 39362 2372
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41049 2363 41107 2369
rect 41049 2360 41061 2363
rect 40644 2332 41061 2360
rect 40644 2320 40650 2332
rect 41049 2329 41061 2332
rect 41095 2329 41107 2363
rect 41049 2323 41107 2329
rect 45373 2363 45431 2369
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46842 2360 46848 2372
rect 45419 2332 46848 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46842 2320 46848 2332
rect 46900 2320 46906 2372
rect 38470 2292 38476 2304
rect 35866 2264 38476 2292
rect 30653 2255 30711 2261
rect 38470 2252 38476 2264
rect 38528 2252 38534 2304
rect 45462 2292 45468 2304
rect 45423 2264 45468 2292
rect 45462 2252 45468 2264
rect 45520 2252 45526 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 15562 1980 15568 2032
rect 15620 2020 15626 2032
rect 36354 2020 36360 2032
rect 15620 1992 36360 2020
rect 15620 1980 15626 1992
rect 36354 1980 36360 1992
rect 36412 1980 36418 2032
rect 3970 1912 3976 1964
rect 4028 1952 4034 1964
rect 16022 1952 16028 1964
rect 4028 1924 16028 1952
rect 4028 1912 4034 1924
rect 16022 1912 16028 1924
rect 16080 1912 16086 1964
rect 29270 1912 29276 1964
rect 29328 1952 29334 1964
rect 45462 1952 45468 1964
rect 29328 1924 45468 1952
rect 29328 1912 29334 1924
rect 45462 1912 45468 1924
rect 45520 1912 45526 1964
rect 19334 1504 19340 1556
rect 19392 1544 19398 1556
rect 25590 1544 25596 1556
rect 19392 1516 25596 1544
rect 19392 1504 19398 1516
rect 25590 1504 25596 1516
rect 25648 1504 25654 1556
<< via1 >>
rect 12624 47404 12676 47456
rect 15844 47404 15896 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 40592 47200 40644 47252
rect 12256 47064 12308 47116
rect 12624 47107 12676 47116
rect 12624 47073 12633 47107
rect 12633 47073 12667 47107
rect 12667 47073 12676 47107
rect 12624 47064 12676 47073
rect 13820 47064 13872 47116
rect 1952 46996 2004 47048
rect 3240 46996 3292 47048
rect 4804 47039 4856 47048
rect 4804 47005 4813 47039
rect 4813 47005 4847 47039
rect 4847 47005 4856 47039
rect 4804 46996 4856 47005
rect 5816 46996 5868 47048
rect 7288 47039 7340 47048
rect 7288 47005 7297 47039
rect 7297 47005 7331 47039
rect 7331 47005 7340 47039
rect 7288 46996 7340 47005
rect 9036 46996 9088 47048
rect 4068 46971 4120 46980
rect 2596 46860 2648 46912
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 6644 46971 6696 46980
rect 6644 46937 6653 46971
rect 6653 46937 6687 46971
rect 6687 46937 6696 46971
rect 6644 46928 6696 46937
rect 9496 46928 9548 46980
rect 4896 46903 4948 46912
rect 4896 46869 4905 46903
rect 4905 46869 4939 46903
rect 4939 46869 4948 46903
rect 4896 46860 4948 46869
rect 7472 46903 7524 46912
rect 7472 46869 7481 46903
rect 7481 46869 7515 46903
rect 7515 46869 7524 46903
rect 7472 46860 7524 46869
rect 12900 46860 12952 46912
rect 15016 46928 15068 46980
rect 16488 46996 16540 47048
rect 21180 47064 21232 47116
rect 29092 47132 29144 47184
rect 30380 47132 30432 47184
rect 48044 47132 48096 47184
rect 35440 47064 35492 47116
rect 43168 47107 43220 47116
rect 43168 47073 43177 47107
rect 43177 47073 43211 47107
rect 43211 47073 43220 47107
rect 43168 47064 43220 47073
rect 48320 47064 48372 47116
rect 18696 46996 18748 47048
rect 20352 46996 20404 47048
rect 20904 47039 20956 47048
rect 20904 47005 20913 47039
rect 20913 47005 20947 47039
rect 20947 47005 20956 47039
rect 20904 46996 20956 47005
rect 19524 46971 19576 46980
rect 19524 46937 19533 46971
rect 19533 46937 19567 46971
rect 19567 46937 19576 46971
rect 19524 46928 19576 46937
rect 19984 46860 20036 46912
rect 24860 47039 24912 47048
rect 24860 47005 24869 47039
rect 24869 47005 24903 47039
rect 24903 47005 24912 47039
rect 24860 46996 24912 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 30932 46996 30984 47048
rect 38108 46996 38160 47048
rect 40224 46996 40276 47048
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 28816 46928 28868 46980
rect 21824 46903 21876 46912
rect 21824 46869 21833 46903
rect 21833 46869 21867 46903
rect 21867 46869 21876 46903
rect 21824 46860 21876 46869
rect 39304 46860 39356 46912
rect 43168 46928 43220 46980
rect 45376 46971 45428 46980
rect 45376 46937 45385 46971
rect 45385 46937 45419 46971
rect 45419 46937 45428 46971
rect 45376 46928 45428 46937
rect 41236 46860 41288 46912
rect 41788 46860 41840 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 3884 46588 3936 46640
rect 10968 46588 11020 46640
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 24860 46588 24912 46640
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 47952 46563 48004 46572
rect 47952 46529 47961 46563
rect 47961 46529 47995 46563
rect 47995 46529 48004 46563
rect 47952 46520 48004 46529
rect 3976 46495 4028 46504
rect 3976 46461 3985 46495
rect 3985 46461 4019 46495
rect 4019 46461 4028 46495
rect 3976 46452 4028 46461
rect 5356 46452 5408 46504
rect 13084 46452 13136 46504
rect 13820 46495 13872 46504
rect 13820 46461 13829 46495
rect 13829 46461 13863 46495
rect 13863 46461 13872 46495
rect 13820 46452 13872 46461
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 14280 46452 14332 46461
rect 20168 46452 20220 46504
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32312 46495 32364 46504
rect 32312 46461 32321 46495
rect 32321 46461 32355 46495
rect 32355 46461 32364 46495
rect 32312 46452 32364 46461
rect 38292 46495 38344 46504
rect 32220 46384 32272 46436
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 42524 46384 42576 46436
rect 46664 46452 46716 46504
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 45468 46384 45520 46436
rect 1492 46316 1544 46368
rect 41328 46316 41380 46368
rect 47768 46316 47820 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3976 46112 4028 46164
rect 5356 46155 5408 46164
rect 5356 46121 5365 46155
rect 5365 46121 5399 46155
rect 5399 46121 5408 46155
rect 5356 46112 5408 46121
rect 13084 46155 13136 46164
rect 13084 46121 13093 46155
rect 13093 46121 13127 46155
rect 13127 46121 13136 46155
rect 13084 46112 13136 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 20168 46155 20220 46164
rect 20168 46121 20177 46155
rect 20177 46121 20211 46155
rect 20211 46121 20220 46155
rect 20168 46112 20220 46121
rect 1768 45908 1820 45960
rect 11612 45976 11664 46028
rect 14096 46044 14148 46096
rect 20720 46112 20772 46164
rect 24768 46155 24820 46164
rect 24768 46121 24777 46155
rect 24777 46121 24811 46155
rect 24811 46121 24820 46155
rect 24768 46112 24820 46121
rect 32312 46112 32364 46164
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 20904 45976 20956 46028
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 13912 45908 13964 45960
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 26240 45976 26292 46028
rect 17316 45840 17368 45892
rect 20904 45883 20956 45892
rect 20904 45849 20913 45883
rect 20913 45849 20947 45883
rect 20947 45849 20956 45883
rect 20904 45840 20956 45849
rect 25504 45883 25556 45892
rect 25504 45849 25513 45883
rect 25513 45849 25547 45883
rect 25547 45849 25556 45883
rect 25504 45840 25556 45849
rect 14096 45772 14148 45824
rect 20076 45772 20128 45824
rect 25780 45772 25832 45824
rect 39396 46044 39448 46096
rect 42984 46044 43036 46096
rect 41328 46019 41380 46028
rect 41328 45985 41337 46019
rect 41337 45985 41371 46019
rect 41371 45985 41380 46019
rect 41328 45976 41380 45985
rect 41880 46019 41932 46028
rect 41880 45985 41889 46019
rect 41889 45985 41923 46019
rect 41923 45985 41932 46019
rect 41880 45976 41932 45985
rect 45836 45976 45888 46028
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 31760 45951 31812 45960
rect 31760 45917 31769 45951
rect 31769 45917 31803 45951
rect 31803 45917 31812 45951
rect 31760 45908 31812 45917
rect 38200 45951 38252 45960
rect 38200 45917 38209 45951
rect 38209 45917 38243 45951
rect 38243 45917 38252 45951
rect 38200 45908 38252 45917
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 41512 45883 41564 45892
rect 41512 45849 41521 45883
rect 41521 45849 41555 45883
rect 41555 45849 41564 45883
rect 41512 45840 41564 45849
rect 31024 45772 31076 45824
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 44088 45815 44140 45824
rect 44088 45781 44097 45815
rect 44097 45781 44131 45815
rect 44131 45781 44140 45815
rect 44088 45772 44140 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 20904 45568 20956 45620
rect 24768 45568 24820 45620
rect 25504 45611 25556 45620
rect 25504 45577 25513 45611
rect 25513 45577 25547 45611
rect 25547 45577 25556 45611
rect 25504 45568 25556 45577
rect 31024 45568 31076 45620
rect 31760 45568 31812 45620
rect 39396 45568 39448 45620
rect 41512 45568 41564 45620
rect 42616 45568 42668 45620
rect 45100 45568 45152 45620
rect 43168 45543 43220 45552
rect 43168 45509 43177 45543
rect 43177 45509 43211 45543
rect 43211 45509 43220 45543
rect 43168 45500 43220 45509
rect 44180 45500 44232 45552
rect 1768 45475 1820 45484
rect 1768 45441 1777 45475
rect 1777 45441 1811 45475
rect 1811 45441 1820 45475
rect 1768 45432 1820 45441
rect 13820 45432 13872 45484
rect 20720 45475 20772 45484
rect 20720 45441 20729 45475
rect 20729 45441 20763 45475
rect 20763 45441 20772 45475
rect 20720 45432 20772 45441
rect 38660 45432 38712 45484
rect 41328 45475 41380 45484
rect 41328 45441 41337 45475
rect 41337 45441 41371 45475
rect 41371 45441 41380 45475
rect 41328 45432 41380 45441
rect 43076 45475 43128 45484
rect 2228 45364 2280 45416
rect 2780 45407 2832 45416
rect 2780 45373 2789 45407
rect 2789 45373 2823 45407
rect 2823 45373 2832 45407
rect 2780 45364 2832 45373
rect 26240 45407 26292 45416
rect 26240 45373 26249 45407
rect 26249 45373 26283 45407
rect 26283 45373 26292 45407
rect 43076 45441 43085 45475
rect 43085 45441 43119 45475
rect 43119 45441 43128 45475
rect 43076 45432 43128 45441
rect 45652 45500 45704 45552
rect 44456 45407 44508 45416
rect 26240 45364 26292 45373
rect 44456 45373 44465 45407
rect 44465 45373 44499 45407
rect 44499 45373 44508 45407
rect 44456 45364 44508 45373
rect 45100 45364 45152 45416
rect 46664 45500 46716 45552
rect 46756 45475 46808 45484
rect 46756 45441 46765 45475
rect 46765 45441 46799 45475
rect 46799 45441 46808 45475
rect 46756 45432 46808 45441
rect 38200 45296 38252 45348
rect 43904 45271 43956 45280
rect 43904 45237 43913 45271
rect 43913 45237 43947 45271
rect 43947 45237 43956 45271
rect 43904 45228 43956 45237
rect 47308 45228 47360 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 2228 45067 2280 45076
rect 2228 45033 2237 45067
rect 2237 45033 2271 45067
rect 2271 45033 2280 45067
rect 2228 45024 2280 45033
rect 44456 45024 44508 45076
rect 45100 45067 45152 45076
rect 45100 45033 45109 45067
rect 45109 45033 45143 45067
rect 45143 45033 45152 45067
rect 45100 45024 45152 45033
rect 46480 45024 46532 45076
rect 43076 44956 43128 45008
rect 47492 44956 47544 45008
rect 45192 44888 45244 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 2044 44820 2096 44872
rect 45008 44863 45060 44872
rect 45008 44829 45017 44863
rect 45017 44829 45051 44863
rect 45051 44829 45060 44863
rect 45008 44820 45060 44829
rect 45652 44863 45704 44872
rect 45652 44829 45661 44863
rect 45661 44829 45695 44863
rect 45695 44829 45704 44863
rect 45652 44820 45704 44829
rect 46296 44863 46348 44872
rect 46296 44829 46305 44863
rect 46305 44829 46339 44863
rect 46339 44829 46348 44863
rect 46296 44820 46348 44829
rect 47676 44752 47728 44804
rect 46664 44684 46716 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 45376 44480 45428 44532
rect 47676 44523 47728 44532
rect 47676 44489 47685 44523
rect 47685 44489 47719 44523
rect 47719 44489 47728 44523
rect 47676 44480 47728 44489
rect 41328 44412 41380 44464
rect 45560 44412 45612 44464
rect 45744 44387 45796 44396
rect 45744 44353 45753 44387
rect 45753 44353 45787 44387
rect 45787 44353 45796 44387
rect 45744 44344 45796 44353
rect 46204 44387 46256 44396
rect 46204 44353 46213 44387
rect 46213 44353 46247 44387
rect 46247 44353 46256 44387
rect 46204 44344 46256 44353
rect 31760 44276 31812 44328
rect 38752 44319 38804 44328
rect 38752 44285 38761 44319
rect 38761 44285 38795 44319
rect 38795 44285 38804 44319
rect 38752 44276 38804 44285
rect 40040 44319 40092 44328
rect 40040 44285 40049 44319
rect 40049 44285 40083 44319
rect 40083 44285 40092 44319
rect 40040 44276 40092 44285
rect 45928 44140 45980 44192
rect 46940 44183 46992 44192
rect 46940 44149 46949 44183
rect 46949 44149 46983 44183
rect 46983 44149 46992 44183
rect 46940 44140 46992 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 31760 43936 31812 43988
rect 38752 43979 38804 43988
rect 38752 43945 38761 43979
rect 38761 43945 38795 43979
rect 38795 43945 38804 43979
rect 38752 43936 38804 43945
rect 46296 43936 46348 43988
rect 45928 43800 45980 43852
rect 46940 43800 46992 43852
rect 48228 43800 48280 43852
rect 25780 43732 25832 43784
rect 38660 43775 38712 43784
rect 38660 43741 38669 43775
rect 38669 43741 38703 43775
rect 38703 43741 38712 43775
rect 38660 43732 38712 43741
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 45468 43256 45520 43308
rect 35716 43188 35768 43240
rect 46940 43052 46992 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 46940 42712 46992 42764
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 47492 42168 47544 42220
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47676 41624 47728 41676
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46940 41488 46992 41540
rect 48136 41531 48188 41540
rect 48136 41497 48145 41531
rect 48145 41497 48179 41531
rect 48179 41497 48188 41531
rect 48136 41488 48188 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46940 41259 46992 41268
rect 46940 41225 46949 41259
rect 46949 41225 46983 41259
rect 46983 41225 46992 41259
rect 46940 41216 46992 41225
rect 14096 41080 14148 41132
rect 46664 41080 46716 41132
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 38936 40876 38988 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 1952 40375 2004 40384
rect 1952 40341 1961 40375
rect 1961 40341 1995 40375
rect 1995 40341 2004 40375
rect 1952 40332 2004 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 23572 39448 23624 39500
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 24768 39423 24820 39432
rect 22744 39244 22796 39296
rect 24768 39389 24777 39423
rect 24777 39389 24811 39423
rect 24811 39389 24820 39423
rect 24768 39380 24820 39389
rect 46848 39312 46900 39364
rect 24492 39244 24544 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 21824 38972 21876 39024
rect 23572 39040 23624 39092
rect 46848 39083 46900 39092
rect 46848 39049 46857 39083
rect 46857 39049 46891 39083
rect 46891 39049 46900 39083
rect 46848 39040 46900 39049
rect 22744 39015 22796 39024
rect 22744 38981 22753 39015
rect 22753 38981 22787 39015
rect 22787 38981 22796 39015
rect 22744 38972 22796 38981
rect 23480 38972 23532 39024
rect 44272 38947 44324 38956
rect 44272 38913 44281 38947
rect 44281 38913 44315 38947
rect 44315 38913 44324 38947
rect 44272 38904 44324 38913
rect 45836 38904 45888 38956
rect 47860 38947 47912 38956
rect 47860 38913 47869 38947
rect 47869 38913 47903 38947
rect 47903 38913 47912 38947
rect 47860 38904 47912 38913
rect 21916 38836 21968 38888
rect 44732 38836 44784 38888
rect 46664 38836 46716 38888
rect 20536 38700 20588 38752
rect 24216 38743 24268 38752
rect 24216 38709 24225 38743
rect 24225 38709 24259 38743
rect 24259 38709 24268 38743
rect 24216 38700 24268 38709
rect 44180 38700 44232 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 23480 38496 23532 38548
rect 38660 38496 38712 38548
rect 46756 38496 46808 38548
rect 21088 38428 21140 38480
rect 15844 38292 15896 38344
rect 17224 38292 17276 38344
rect 20352 38335 20404 38344
rect 20352 38301 20361 38335
rect 20361 38301 20395 38335
rect 20395 38301 20404 38335
rect 20352 38292 20404 38301
rect 20628 38292 20680 38344
rect 24492 38428 24544 38480
rect 23664 38360 23716 38412
rect 42984 38403 43036 38412
rect 42984 38369 42993 38403
rect 42993 38369 43027 38403
rect 43027 38369 43036 38403
rect 42984 38360 43036 38369
rect 45008 38360 45060 38412
rect 23572 38292 23624 38344
rect 24216 38292 24268 38344
rect 44272 38292 44324 38344
rect 46296 38335 46348 38344
rect 46296 38301 46305 38335
rect 46305 38301 46339 38335
rect 46339 38301 46348 38335
rect 46296 38292 46348 38301
rect 45468 38224 45520 38276
rect 45560 38224 45612 38276
rect 46848 38224 46900 38276
rect 48136 38267 48188 38276
rect 48136 38233 48145 38267
rect 48145 38233 48179 38267
rect 48179 38233 48188 38267
rect 48136 38224 48188 38233
rect 19248 38156 19300 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 23848 37884 23900 37936
rect 21824 37859 21876 37868
rect 21824 37825 21833 37859
rect 21833 37825 21867 37859
rect 21867 37825 21876 37859
rect 21824 37816 21876 37825
rect 23572 37859 23624 37868
rect 23572 37825 23581 37859
rect 23581 37825 23615 37859
rect 23615 37825 23624 37859
rect 23572 37816 23624 37825
rect 19524 37791 19576 37800
rect 19524 37757 19533 37791
rect 19533 37757 19567 37791
rect 19567 37757 19576 37791
rect 19524 37748 19576 37757
rect 19800 37791 19852 37800
rect 19800 37757 19809 37791
rect 19809 37757 19843 37791
rect 19843 37757 19852 37791
rect 19800 37748 19852 37757
rect 23756 37748 23808 37800
rect 46848 37995 46900 38004
rect 46848 37961 46857 37995
rect 46857 37961 46891 37995
rect 46891 37961 46900 37995
rect 46848 37952 46900 37961
rect 25964 37884 26016 37936
rect 46296 37884 46348 37936
rect 27804 37859 27856 37868
rect 27804 37825 27813 37859
rect 27813 37825 27847 37859
rect 27847 37825 27856 37859
rect 27804 37816 27856 37825
rect 44272 37859 44324 37868
rect 44272 37825 44281 37859
rect 44281 37825 44315 37859
rect 44315 37825 44324 37859
rect 44272 37816 44324 37825
rect 46756 37859 46808 37868
rect 46756 37825 46765 37859
rect 46765 37825 46799 37859
rect 46799 37825 46808 37859
rect 46756 37816 46808 37825
rect 24952 37791 25004 37800
rect 22100 37680 22152 37732
rect 23388 37612 23440 37664
rect 24952 37757 24961 37791
rect 24961 37757 24995 37791
rect 24995 37757 25004 37791
rect 24952 37748 25004 37757
rect 45560 37748 45612 37800
rect 46204 37748 46256 37800
rect 26332 37612 26384 37664
rect 27988 37612 28040 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19800 37408 19852 37460
rect 21824 37408 21876 37460
rect 24952 37408 25004 37460
rect 44272 37451 44324 37460
rect 44272 37417 44281 37451
rect 44281 37417 44315 37451
rect 44315 37417 44324 37451
rect 44272 37408 44324 37417
rect 1768 37204 1820 37256
rect 19248 37204 19300 37256
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 20260 37315 20312 37324
rect 20260 37281 20269 37315
rect 20269 37281 20303 37315
rect 20303 37281 20312 37315
rect 42984 37340 43036 37392
rect 47032 37340 47084 37392
rect 20260 37272 20312 37281
rect 20628 37204 20680 37256
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 17316 37136 17368 37188
rect 19524 37136 19576 37188
rect 19984 37136 20036 37188
rect 22192 37179 22244 37188
rect 22192 37145 22201 37179
rect 22201 37145 22235 37179
rect 22235 37145 22244 37179
rect 22192 37136 22244 37145
rect 25136 37204 25188 37256
rect 25964 37247 26016 37256
rect 25964 37213 25973 37247
rect 25973 37213 26007 37247
rect 26007 37213 26016 37247
rect 25964 37204 26016 37213
rect 26332 37204 26384 37256
rect 43628 37204 43680 37256
rect 44180 37247 44232 37256
rect 44180 37213 44189 37247
rect 44189 37213 44223 37247
rect 44223 37213 44232 37247
rect 44180 37204 44232 37213
rect 26976 37179 27028 37188
rect 23572 37068 23624 37120
rect 23848 37068 23900 37120
rect 26976 37145 26985 37179
rect 26985 37145 27019 37179
rect 27019 37145 27028 37179
rect 26976 37136 27028 37145
rect 27988 37136 28040 37188
rect 27804 37068 27856 37120
rect 28448 37111 28500 37120
rect 28448 37077 28457 37111
rect 28457 37077 28491 37111
rect 28491 37077 28500 37111
rect 28448 37068 28500 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 9496 36864 9548 36916
rect 18328 36796 18380 36848
rect 20076 36864 20128 36916
rect 23664 36864 23716 36916
rect 25780 36907 25832 36916
rect 25780 36873 25789 36907
rect 25789 36873 25823 36907
rect 25823 36873 25832 36907
rect 25780 36864 25832 36873
rect 26976 36907 27028 36916
rect 26976 36873 26985 36907
rect 26985 36873 27019 36907
rect 27019 36873 27028 36907
rect 26976 36864 27028 36873
rect 27804 36864 27856 36916
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 16028 36728 16080 36780
rect 17316 36771 17368 36780
rect 17316 36737 17325 36771
rect 17325 36737 17359 36771
rect 17359 36737 17368 36771
rect 17316 36728 17368 36737
rect 20444 36728 20496 36780
rect 20628 36728 20680 36780
rect 21824 36771 21876 36780
rect 21824 36737 21833 36771
rect 21833 36737 21867 36771
rect 21867 36737 21876 36771
rect 21824 36728 21876 36737
rect 23480 36728 23532 36780
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 18236 36660 18288 36712
rect 22100 36703 22152 36712
rect 22100 36669 22109 36703
rect 22109 36669 22143 36703
rect 22143 36669 22152 36703
rect 22100 36660 22152 36669
rect 23204 36592 23256 36644
rect 25228 36728 25280 36780
rect 27252 36771 27304 36780
rect 27252 36737 27261 36771
rect 27261 36737 27295 36771
rect 27295 36737 27304 36771
rect 27528 36771 27580 36780
rect 27252 36728 27304 36737
rect 27528 36737 27537 36771
rect 27537 36737 27571 36771
rect 27571 36737 27580 36771
rect 27528 36728 27580 36737
rect 27988 36703 28040 36712
rect 27988 36669 27997 36703
rect 27997 36669 28031 36703
rect 28031 36669 28040 36703
rect 27988 36660 28040 36669
rect 28448 36660 28500 36712
rect 27528 36592 27580 36644
rect 15752 36524 15804 36576
rect 19064 36567 19116 36576
rect 19064 36533 19073 36567
rect 19073 36533 19107 36567
rect 19107 36533 19116 36567
rect 19064 36524 19116 36533
rect 24860 36524 24912 36576
rect 29368 36524 29420 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 2320 36116 2372 36168
rect 45560 36320 45612 36372
rect 18236 36295 18288 36304
rect 18236 36261 18245 36295
rect 18245 36261 18279 36295
rect 18279 36261 18288 36295
rect 18236 36252 18288 36261
rect 17316 36184 17368 36236
rect 17408 36184 17460 36236
rect 15292 36048 15344 36100
rect 15752 36048 15804 36100
rect 16396 35980 16448 36032
rect 20076 36184 20128 36236
rect 22192 36252 22244 36304
rect 23480 36252 23532 36304
rect 24952 36295 25004 36304
rect 24952 36261 24961 36295
rect 24961 36261 24995 36295
rect 24995 36261 25004 36295
rect 24952 36252 25004 36261
rect 25136 36295 25188 36304
rect 25136 36261 25145 36295
rect 25145 36261 25179 36295
rect 25179 36261 25188 36295
rect 25136 36252 25188 36261
rect 22928 36184 22980 36236
rect 23020 36184 23072 36236
rect 19064 36116 19116 36168
rect 19248 36116 19300 36168
rect 22560 36116 22612 36168
rect 25228 36184 25280 36236
rect 18972 36048 19024 36100
rect 23848 36116 23900 36168
rect 27988 36116 28040 36168
rect 19340 35980 19392 36032
rect 23480 36048 23532 36100
rect 25136 36048 25188 36100
rect 27528 36048 27580 36100
rect 23020 36023 23072 36032
rect 23020 35989 23029 36023
rect 23029 35989 23063 36023
rect 23063 35989 23072 36023
rect 23020 35980 23072 35989
rect 24032 35980 24084 36032
rect 27804 36023 27856 36032
rect 27804 35989 27813 36023
rect 27813 35989 27847 36023
rect 27847 35989 27856 36023
rect 27804 35980 27856 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 18328 35819 18380 35828
rect 18328 35785 18337 35819
rect 18337 35785 18371 35819
rect 18371 35785 18380 35819
rect 18328 35776 18380 35785
rect 19340 35776 19392 35828
rect 23204 35819 23256 35828
rect 23204 35785 23213 35819
rect 23213 35785 23247 35819
rect 23247 35785 23256 35819
rect 23204 35776 23256 35785
rect 23756 35776 23808 35828
rect 25136 35819 25188 35828
rect 25136 35785 25145 35819
rect 25145 35785 25179 35819
rect 25179 35785 25188 35819
rect 25136 35776 25188 35785
rect 27252 35819 27304 35828
rect 27252 35785 27261 35819
rect 27261 35785 27295 35819
rect 27295 35785 27304 35819
rect 27252 35776 27304 35785
rect 27804 35776 27856 35828
rect 16028 35708 16080 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 16580 35640 16632 35692
rect 17224 35683 17276 35692
rect 15752 35572 15804 35624
rect 16120 35572 16172 35624
rect 16396 35572 16448 35624
rect 17224 35649 17233 35683
rect 17233 35649 17267 35683
rect 17267 35649 17276 35683
rect 17224 35640 17276 35649
rect 19248 35751 19300 35760
rect 19248 35717 19253 35751
rect 19253 35717 19287 35751
rect 19287 35717 19300 35751
rect 19248 35708 19300 35717
rect 20260 35708 20312 35760
rect 21916 35708 21968 35760
rect 18328 35640 18380 35692
rect 18972 35683 19024 35692
rect 18972 35649 18981 35683
rect 18981 35649 19015 35683
rect 19015 35649 19024 35683
rect 18972 35640 19024 35649
rect 17132 35615 17184 35624
rect 17132 35581 17141 35615
rect 17141 35581 17175 35615
rect 17175 35581 17184 35615
rect 17132 35572 17184 35581
rect 16948 35504 17000 35556
rect 21824 35640 21876 35692
rect 22652 35640 22704 35692
rect 23756 35640 23808 35692
rect 24584 35708 24636 35760
rect 26332 35708 26384 35760
rect 27528 35708 27580 35760
rect 20260 35504 20312 35556
rect 23572 35572 23624 35624
rect 24032 35615 24084 35624
rect 24032 35581 24041 35615
rect 24041 35581 24075 35615
rect 24075 35581 24084 35615
rect 24032 35572 24084 35581
rect 24124 35615 24176 35624
rect 24124 35581 24133 35615
rect 24133 35581 24167 35615
rect 24167 35581 24176 35615
rect 24124 35572 24176 35581
rect 24768 35572 24820 35624
rect 26976 35640 27028 35692
rect 26332 35572 26384 35624
rect 23112 35504 23164 35556
rect 24676 35504 24728 35556
rect 27988 35640 28040 35692
rect 29368 35708 29420 35760
rect 48136 35683 48188 35692
rect 48136 35649 48145 35683
rect 48145 35649 48179 35683
rect 48179 35649 48188 35683
rect 48136 35640 48188 35649
rect 29368 35572 29420 35624
rect 2228 35436 2280 35488
rect 15936 35436 15988 35488
rect 16672 35479 16724 35488
rect 16672 35445 16681 35479
rect 16681 35445 16715 35479
rect 16715 35445 16724 35479
rect 16672 35436 16724 35445
rect 23020 35479 23072 35488
rect 23020 35445 23029 35479
rect 23029 35445 23063 35479
rect 23063 35445 23072 35479
rect 23020 35436 23072 35445
rect 23204 35436 23256 35488
rect 26240 35479 26292 35488
rect 26240 35445 26249 35479
rect 26249 35445 26283 35479
rect 26283 35445 26292 35479
rect 26240 35436 26292 35445
rect 26424 35436 26476 35488
rect 28356 35436 28408 35488
rect 28908 35436 28960 35488
rect 47124 35436 47176 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 15292 35232 15344 35284
rect 15936 35275 15988 35284
rect 15936 35241 15945 35275
rect 15945 35241 15979 35275
rect 15979 35241 15988 35275
rect 15936 35232 15988 35241
rect 20812 35232 20864 35284
rect 22560 35232 22612 35284
rect 22652 35232 22704 35284
rect 23480 35232 23532 35284
rect 24952 35232 25004 35284
rect 25412 35232 25464 35284
rect 26424 35232 26476 35284
rect 27988 35232 28040 35284
rect 16672 35096 16724 35148
rect 15936 35028 15988 35080
rect 18328 35071 18380 35080
rect 18328 35037 18337 35071
rect 18337 35037 18371 35071
rect 18371 35037 18380 35071
rect 18328 35028 18380 35037
rect 21456 35096 21508 35148
rect 22744 35096 22796 35148
rect 21732 35071 21784 35080
rect 16580 34960 16632 35012
rect 21732 35037 21741 35071
rect 21741 35037 21775 35071
rect 21775 35037 21784 35071
rect 21732 35028 21784 35037
rect 22836 35028 22888 35080
rect 22100 34960 22152 35012
rect 18420 34935 18472 34944
rect 18420 34901 18429 34935
rect 18429 34901 18463 34935
rect 18463 34901 18472 34935
rect 18420 34892 18472 34901
rect 22284 34892 22336 34944
rect 24124 35164 24176 35216
rect 26332 35164 26384 35216
rect 24032 35096 24084 35148
rect 23940 35028 23992 35080
rect 23112 35003 23164 35012
rect 23112 34969 23121 35003
rect 23121 34969 23155 35003
rect 23155 34969 23164 35003
rect 23112 34960 23164 34969
rect 23296 35003 23348 35012
rect 23296 34969 23331 35003
rect 23331 34969 23348 35003
rect 24492 35028 24544 35080
rect 23296 34960 23348 34969
rect 24952 35096 25004 35148
rect 26240 35096 26292 35148
rect 25412 35071 25464 35080
rect 25412 35037 25421 35071
rect 25421 35037 25455 35071
rect 25455 35037 25464 35071
rect 25412 35028 25464 35037
rect 24768 34960 24820 35012
rect 25596 35028 25648 35080
rect 26424 35028 26476 35080
rect 27160 35071 27212 35080
rect 27160 35037 27169 35071
rect 27169 35037 27203 35071
rect 27203 35037 27212 35071
rect 27160 35028 27212 35037
rect 27068 34960 27120 35012
rect 27804 35028 27856 35080
rect 28448 35071 28500 35080
rect 28448 35037 28457 35071
rect 28457 35037 28491 35071
rect 28491 35037 28500 35071
rect 28448 35028 28500 35037
rect 29828 35028 29880 35080
rect 30380 35071 30432 35080
rect 30380 35037 30389 35071
rect 30389 35037 30423 35071
rect 30423 35037 30432 35071
rect 30380 35028 30432 35037
rect 48228 35028 48280 35080
rect 28908 34960 28960 35012
rect 29000 34960 29052 35012
rect 26148 34892 26200 34944
rect 28632 34892 28684 34944
rect 29460 34892 29512 34944
rect 30748 34892 30800 34944
rect 47860 34892 47912 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 18420 34620 18472 34672
rect 16028 34552 16080 34604
rect 17316 34552 17368 34604
rect 21272 34620 21324 34672
rect 22100 34688 22152 34740
rect 21916 34620 21968 34672
rect 20812 34552 20864 34604
rect 21456 34552 21508 34604
rect 17684 34527 17736 34536
rect 17684 34493 17693 34527
rect 17693 34493 17727 34527
rect 17727 34493 17736 34527
rect 17684 34484 17736 34493
rect 21180 34484 21232 34536
rect 22836 34484 22888 34536
rect 23388 34620 23440 34672
rect 23572 34620 23624 34672
rect 26332 34688 26384 34740
rect 25044 34620 25096 34672
rect 25596 34620 25648 34672
rect 27068 34688 27120 34740
rect 27436 34688 27488 34740
rect 29368 34731 29420 34740
rect 29368 34697 29377 34731
rect 29377 34697 29411 34731
rect 29411 34697 29420 34731
rect 29368 34688 29420 34697
rect 26516 34620 26568 34672
rect 29460 34620 29512 34672
rect 31392 34620 31444 34672
rect 26976 34595 27028 34604
rect 26976 34561 26985 34595
rect 26985 34561 27019 34595
rect 27019 34561 27028 34595
rect 26976 34552 27028 34561
rect 27160 34595 27212 34604
rect 27160 34561 27169 34595
rect 27169 34561 27203 34595
rect 27203 34561 27212 34595
rect 27160 34552 27212 34561
rect 28632 34595 28684 34604
rect 28632 34561 28641 34595
rect 28641 34561 28675 34595
rect 28675 34561 28684 34595
rect 28632 34552 28684 34561
rect 25412 34527 25464 34536
rect 21732 34416 21784 34468
rect 22100 34416 22152 34468
rect 25412 34493 25421 34527
rect 25421 34493 25455 34527
rect 25455 34493 25464 34527
rect 25412 34484 25464 34493
rect 26240 34484 26292 34536
rect 28540 34484 28592 34536
rect 28908 34595 28960 34604
rect 28908 34561 28917 34595
rect 28917 34561 28951 34595
rect 28951 34561 28960 34595
rect 29184 34595 29236 34604
rect 28908 34552 28960 34561
rect 29184 34561 29193 34595
rect 29193 34561 29227 34595
rect 29227 34561 29236 34595
rect 29184 34552 29236 34561
rect 30748 34595 30800 34604
rect 30748 34561 30757 34595
rect 30757 34561 30791 34595
rect 30791 34561 30800 34595
rect 30748 34552 30800 34561
rect 31024 34595 31076 34604
rect 31024 34561 31033 34595
rect 31033 34561 31067 34595
rect 31067 34561 31076 34595
rect 47768 34595 47820 34604
rect 31024 34552 31076 34561
rect 47768 34561 47777 34595
rect 47777 34561 47811 34595
rect 47811 34561 47820 34595
rect 47768 34552 47820 34561
rect 29276 34484 29328 34536
rect 15476 34348 15528 34400
rect 19064 34348 19116 34400
rect 20720 34348 20772 34400
rect 21824 34391 21876 34400
rect 21824 34357 21833 34391
rect 21833 34357 21867 34391
rect 21867 34357 21876 34391
rect 21824 34348 21876 34357
rect 22192 34348 22244 34400
rect 26516 34416 26568 34468
rect 26976 34416 27028 34468
rect 26884 34348 26936 34400
rect 27068 34391 27120 34400
rect 27068 34357 27077 34391
rect 27077 34357 27111 34391
rect 27111 34357 27120 34391
rect 27068 34348 27120 34357
rect 30564 34391 30616 34400
rect 30564 34357 30573 34391
rect 30573 34357 30607 34391
rect 30607 34357 30616 34391
rect 30564 34348 30616 34357
rect 47216 34348 47268 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 1952 34144 2004 34196
rect 17316 34076 17368 34128
rect 17684 34144 17736 34196
rect 21732 34187 21784 34196
rect 21732 34153 21741 34187
rect 21741 34153 21775 34187
rect 21775 34153 21784 34187
rect 21732 34144 21784 34153
rect 22284 34187 22336 34196
rect 22284 34153 22293 34187
rect 22293 34153 22327 34187
rect 22327 34153 22336 34187
rect 22284 34144 22336 34153
rect 23572 34187 23624 34196
rect 23572 34153 23581 34187
rect 23581 34153 23615 34187
rect 23615 34153 23624 34187
rect 23572 34144 23624 34153
rect 24492 34144 24544 34196
rect 24676 34144 24728 34196
rect 16856 34051 16908 34060
rect 16856 34017 16865 34051
rect 16865 34017 16899 34051
rect 16899 34017 16908 34051
rect 21272 34076 21324 34128
rect 30380 34144 30432 34196
rect 30564 34144 30616 34196
rect 16856 34008 16908 34017
rect 19984 34051 20036 34060
rect 19984 34017 19993 34051
rect 19993 34017 20027 34051
rect 20027 34017 20036 34051
rect 19984 34008 20036 34017
rect 20720 34008 20772 34060
rect 1584 33983 1636 33992
rect 1584 33949 1593 33983
rect 1593 33949 1627 33983
rect 1627 33949 1636 33983
rect 1584 33940 1636 33949
rect 16580 33983 16632 33992
rect 16580 33949 16589 33983
rect 16589 33949 16623 33983
rect 16623 33949 16632 33983
rect 16580 33940 16632 33949
rect 16948 33983 17000 33992
rect 14464 33915 14516 33924
rect 14464 33881 14473 33915
rect 14473 33881 14507 33915
rect 14507 33881 14516 33915
rect 14464 33872 14516 33881
rect 15476 33872 15528 33924
rect 1952 33804 2004 33856
rect 16304 33872 16356 33924
rect 16948 33949 16957 33983
rect 16957 33949 16991 33983
rect 16991 33949 17000 33983
rect 16948 33940 17000 33949
rect 17776 33983 17828 33992
rect 17776 33949 17785 33983
rect 17785 33949 17819 33983
rect 17819 33949 17828 33983
rect 17776 33940 17828 33949
rect 17960 33983 18012 33992
rect 17960 33949 17969 33983
rect 17969 33949 18003 33983
rect 18003 33949 18012 33983
rect 17960 33940 18012 33949
rect 18328 33983 18380 33992
rect 18328 33949 18337 33983
rect 18337 33949 18371 33983
rect 18371 33949 18380 33983
rect 18328 33940 18380 33949
rect 19064 33872 19116 33924
rect 20996 33872 21048 33924
rect 16396 33847 16448 33856
rect 16396 33813 16405 33847
rect 16405 33813 16439 33847
rect 16439 33813 16448 33847
rect 16396 33804 16448 33813
rect 20076 33804 20128 33856
rect 21824 34008 21876 34060
rect 27528 34076 27580 34128
rect 22008 33940 22060 33992
rect 22468 33983 22520 33992
rect 22468 33949 22477 33983
rect 22477 33949 22511 33983
rect 22511 33949 22520 33983
rect 22468 33940 22520 33949
rect 22100 33872 22152 33924
rect 27344 34008 27396 34060
rect 29920 34051 29972 34060
rect 29920 34017 29929 34051
rect 29929 34017 29963 34051
rect 29963 34017 29972 34051
rect 29920 34008 29972 34017
rect 32128 34008 32180 34060
rect 47124 34051 47176 34060
rect 47124 34017 47133 34051
rect 47133 34017 47167 34051
rect 47167 34017 47176 34051
rect 47124 34008 47176 34017
rect 47400 34051 47452 34060
rect 47400 34017 47409 34051
rect 47409 34017 47443 34051
rect 47443 34017 47452 34051
rect 47400 34008 47452 34017
rect 24584 33940 24636 33992
rect 26148 33983 26200 33992
rect 26148 33949 26157 33983
rect 26157 33949 26191 33983
rect 26191 33949 26200 33983
rect 26148 33940 26200 33949
rect 26240 33983 26292 33992
rect 26240 33949 26249 33983
rect 26249 33949 26283 33983
rect 26283 33949 26292 33983
rect 26240 33940 26292 33949
rect 25412 33872 25464 33924
rect 26884 33940 26936 33992
rect 27436 33940 27488 33992
rect 29828 33940 29880 33992
rect 25964 33847 26016 33856
rect 25964 33813 25973 33847
rect 25973 33813 26007 33847
rect 26007 33813 26016 33847
rect 25964 33804 26016 33813
rect 26148 33804 26200 33856
rect 31024 33804 31076 33856
rect 32864 33872 32916 33924
rect 47216 33915 47268 33924
rect 47216 33881 47225 33915
rect 47225 33881 47259 33915
rect 47259 33881 47268 33915
rect 47216 33872 47268 33881
rect 32588 33847 32640 33856
rect 32588 33813 32597 33847
rect 32597 33813 32631 33847
rect 32631 33813 32640 33847
rect 32588 33804 32640 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 14464 33600 14516 33652
rect 17776 33600 17828 33652
rect 19984 33600 20036 33652
rect 20628 33600 20680 33652
rect 14464 33507 14516 33516
rect 14464 33473 14473 33507
rect 14473 33473 14507 33507
rect 14507 33473 14516 33507
rect 14464 33464 14516 33473
rect 15752 33532 15804 33584
rect 16396 33464 16448 33516
rect 17868 33507 17920 33516
rect 17868 33473 17877 33507
rect 17877 33473 17911 33507
rect 17911 33473 17920 33507
rect 17868 33464 17920 33473
rect 19064 33507 19116 33516
rect 19064 33473 19073 33507
rect 19073 33473 19107 33507
rect 19107 33473 19116 33507
rect 19064 33464 19116 33473
rect 19248 33464 19300 33516
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 1860 33396 1912 33448
rect 15936 33396 15988 33448
rect 20352 33464 20404 33516
rect 21640 33464 21692 33516
rect 22192 33532 22244 33584
rect 27528 33600 27580 33652
rect 32864 33643 32916 33652
rect 32864 33609 32873 33643
rect 32873 33609 32907 33643
rect 32907 33609 32916 33643
rect 32864 33600 32916 33609
rect 47768 33600 47820 33652
rect 29368 33575 29420 33584
rect 29368 33541 29377 33575
rect 29377 33541 29411 33575
rect 29411 33541 29420 33575
rect 29368 33532 29420 33541
rect 22008 33464 22060 33516
rect 24584 33464 24636 33516
rect 25964 33507 26016 33516
rect 25964 33473 25973 33507
rect 25973 33473 26007 33507
rect 26007 33473 26016 33507
rect 25964 33464 26016 33473
rect 26148 33507 26200 33516
rect 26148 33473 26157 33507
rect 26157 33473 26191 33507
rect 26191 33473 26200 33507
rect 26148 33464 26200 33473
rect 27528 33464 27580 33516
rect 28356 33464 28408 33516
rect 30012 33464 30064 33516
rect 32312 33464 32364 33516
rect 32864 33464 32916 33516
rect 46848 33507 46900 33516
rect 46848 33473 46857 33507
rect 46857 33473 46891 33507
rect 46891 33473 46900 33507
rect 46848 33464 46900 33473
rect 19984 33396 20036 33448
rect 22468 33328 22520 33380
rect 23112 33328 23164 33380
rect 25596 33396 25648 33448
rect 26056 33396 26108 33448
rect 46664 33396 46716 33448
rect 18236 33303 18288 33312
rect 18236 33269 18245 33303
rect 18245 33269 18279 33303
rect 18279 33269 18288 33303
rect 18236 33260 18288 33269
rect 20076 33260 20128 33312
rect 21548 33260 21600 33312
rect 25596 33260 25648 33312
rect 25688 33260 25740 33312
rect 28632 33328 28684 33380
rect 31392 33328 31444 33380
rect 29552 33303 29604 33312
rect 29552 33269 29576 33303
rect 29576 33269 29604 33303
rect 29552 33260 29604 33269
rect 29920 33260 29972 33312
rect 32220 33303 32272 33312
rect 32220 33269 32229 33303
rect 32229 33269 32263 33303
rect 32263 33269 32272 33303
rect 32220 33260 32272 33269
rect 44180 33260 44232 33312
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1952 33099 2004 33108
rect 1952 33065 1961 33099
rect 1961 33065 1995 33099
rect 1995 33065 2004 33099
rect 1952 33056 2004 33065
rect 14464 33056 14516 33108
rect 1952 32852 2004 32904
rect 14464 32852 14516 32904
rect 15936 33056 15988 33108
rect 17132 33099 17184 33108
rect 17132 33065 17141 33099
rect 17141 33065 17175 33099
rect 17175 33065 17184 33099
rect 17132 33056 17184 33065
rect 17316 33056 17368 33108
rect 20996 33056 21048 33108
rect 21640 33056 21692 33108
rect 15752 33031 15804 33040
rect 15752 32997 15761 33031
rect 15761 32997 15795 33031
rect 15795 32997 15804 33031
rect 15752 32988 15804 32997
rect 16304 32988 16356 33040
rect 16396 32988 16448 33040
rect 15108 32852 15160 32904
rect 16120 32784 16172 32836
rect 16396 32827 16448 32836
rect 16396 32793 16405 32827
rect 16405 32793 16439 32827
rect 16439 32793 16448 32827
rect 17408 32895 17460 32904
rect 17408 32861 17417 32895
rect 17417 32861 17451 32895
rect 17451 32861 17460 32895
rect 17408 32852 17460 32861
rect 29368 33056 29420 33108
rect 22744 32988 22796 33040
rect 23204 32988 23256 33040
rect 24860 33031 24912 33040
rect 24860 32997 24869 33031
rect 24869 32997 24903 33031
rect 24903 32997 24912 33031
rect 24860 32988 24912 32997
rect 27160 33031 27212 33040
rect 27160 32997 27169 33031
rect 27169 32997 27203 33031
rect 27203 32997 27212 33031
rect 27160 32988 27212 32997
rect 29920 32988 29972 33040
rect 26976 32920 27028 32972
rect 27436 32920 27488 32972
rect 29552 32920 29604 32972
rect 30288 32988 30340 33040
rect 31668 33056 31720 33108
rect 48044 32988 48096 33040
rect 30380 32963 30432 32972
rect 19248 32895 19300 32904
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 21088 32852 21140 32904
rect 24400 32852 24452 32904
rect 24768 32895 24820 32904
rect 24768 32861 24777 32895
rect 24777 32861 24811 32895
rect 24811 32861 24820 32895
rect 24768 32852 24820 32861
rect 27344 32852 27396 32904
rect 28172 32895 28224 32904
rect 16396 32784 16448 32793
rect 2412 32716 2464 32768
rect 15844 32716 15896 32768
rect 19064 32784 19116 32836
rect 25596 32784 25648 32836
rect 25688 32827 25740 32836
rect 25688 32793 25697 32827
rect 25697 32793 25731 32827
rect 25731 32793 25740 32827
rect 25688 32784 25740 32793
rect 27436 32784 27488 32836
rect 28172 32861 28181 32895
rect 28181 32861 28215 32895
rect 28215 32861 28224 32895
rect 28172 32852 28224 32861
rect 30380 32929 30389 32963
rect 30389 32929 30423 32963
rect 30423 32929 30432 32963
rect 30380 32920 30432 32929
rect 30196 32895 30248 32904
rect 30196 32861 30205 32895
rect 30205 32861 30239 32895
rect 30239 32861 30248 32895
rect 30196 32852 30248 32861
rect 32220 32920 32272 32972
rect 31392 32895 31444 32904
rect 31392 32861 31401 32895
rect 31401 32861 31435 32895
rect 31435 32861 31444 32895
rect 31392 32852 31444 32861
rect 31484 32895 31536 32904
rect 31484 32861 31493 32895
rect 31493 32861 31527 32895
rect 31527 32861 31536 32895
rect 31484 32852 31536 32861
rect 32588 32852 32640 32904
rect 31668 32784 31720 32836
rect 32312 32784 32364 32836
rect 32772 32784 32824 32836
rect 46940 32784 46992 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 22100 32716 22152 32768
rect 22376 32716 22428 32768
rect 23204 32716 23256 32768
rect 27896 32716 27948 32768
rect 28264 32759 28316 32768
rect 28264 32725 28273 32759
rect 28273 32725 28307 32759
rect 28307 32725 28316 32759
rect 28264 32716 28316 32725
rect 29000 32716 29052 32768
rect 29460 32716 29512 32768
rect 30380 32716 30432 32768
rect 31484 32716 31536 32768
rect 31760 32716 31812 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 17408 32512 17460 32564
rect 23388 32512 23440 32564
rect 25596 32555 25648 32564
rect 25596 32521 25605 32555
rect 25605 32521 25639 32555
rect 25639 32521 25648 32555
rect 25596 32512 25648 32521
rect 26148 32512 26200 32564
rect 29920 32512 29972 32564
rect 2412 32487 2464 32496
rect 2412 32453 2421 32487
rect 2421 32453 2455 32487
rect 2455 32453 2464 32487
rect 2412 32444 2464 32453
rect 14740 32444 14792 32496
rect 15108 32444 15160 32496
rect 17868 32444 17920 32496
rect 20076 32444 20128 32496
rect 20628 32444 20680 32496
rect 22376 32487 22428 32496
rect 2228 32419 2280 32428
rect 2228 32385 2237 32419
rect 2237 32385 2271 32419
rect 2271 32385 2280 32419
rect 2228 32376 2280 32385
rect 15844 32419 15896 32428
rect 15844 32385 15853 32419
rect 15853 32385 15887 32419
rect 15887 32385 15896 32419
rect 15844 32376 15896 32385
rect 15936 32419 15988 32428
rect 15936 32385 15945 32419
rect 15945 32385 15979 32419
rect 15979 32385 15988 32419
rect 17224 32419 17276 32428
rect 15936 32376 15988 32385
rect 4620 32308 4672 32360
rect 17224 32385 17233 32419
rect 17233 32385 17267 32419
rect 17267 32385 17276 32419
rect 17224 32376 17276 32385
rect 22376 32453 22385 32487
rect 22385 32453 22419 32487
rect 22419 32453 22428 32487
rect 22376 32444 22428 32453
rect 22652 32444 22704 32496
rect 24768 32444 24820 32496
rect 44180 32512 44232 32564
rect 46940 32555 46992 32564
rect 46940 32521 46949 32555
rect 46949 32521 46983 32555
rect 46983 32521 46992 32555
rect 46940 32512 46992 32521
rect 48044 32555 48096 32564
rect 48044 32521 48053 32555
rect 48053 32521 48087 32555
rect 48087 32521 48096 32555
rect 48044 32512 48096 32521
rect 33048 32444 33100 32496
rect 24308 32419 24360 32428
rect 16212 32308 16264 32360
rect 1400 32172 1452 32224
rect 14464 32172 14516 32224
rect 18236 32240 18288 32292
rect 24308 32385 24317 32419
rect 24317 32385 24351 32419
rect 24351 32385 24360 32419
rect 24308 32376 24360 32385
rect 23664 32308 23716 32360
rect 24676 32308 24728 32360
rect 27804 32376 27856 32428
rect 29368 32376 29420 32428
rect 17592 32172 17644 32224
rect 18328 32172 18380 32224
rect 27344 32240 27396 32292
rect 27896 32308 27948 32360
rect 28816 32308 28868 32360
rect 30012 32376 30064 32428
rect 32128 32419 32180 32428
rect 32128 32385 32137 32419
rect 32137 32385 32171 32419
rect 32171 32385 32180 32419
rect 32128 32376 32180 32385
rect 45560 32376 45612 32428
rect 47952 32419 48004 32428
rect 47952 32385 47961 32419
rect 47961 32385 47995 32419
rect 47995 32385 48004 32419
rect 47952 32376 48004 32385
rect 28908 32240 28960 32292
rect 30196 32308 30248 32360
rect 32496 32308 32548 32360
rect 32772 32308 32824 32360
rect 30932 32240 30984 32292
rect 27252 32172 27304 32224
rect 27712 32172 27764 32224
rect 29000 32172 29052 32224
rect 29184 32172 29236 32224
rect 32220 32172 32272 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 16212 32011 16264 32020
rect 16212 31977 16221 32011
rect 16221 31977 16255 32011
rect 16255 31977 16264 32011
rect 16212 31968 16264 31977
rect 16304 31968 16356 32020
rect 19248 31968 19300 32020
rect 22652 32011 22704 32020
rect 16396 31900 16448 31952
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 1952 31832 2004 31884
rect 4620 31875 4672 31884
rect 4620 31841 4629 31875
rect 4629 31841 4663 31875
rect 4663 31841 4672 31875
rect 4620 31832 4672 31841
rect 5448 31832 5500 31884
rect 16120 31832 16172 31884
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 19340 31832 19392 31884
rect 20076 31875 20128 31884
rect 20076 31841 20085 31875
rect 20085 31841 20119 31875
rect 20119 31841 20128 31875
rect 20076 31832 20128 31841
rect 21088 31832 21140 31884
rect 22652 31977 22661 32011
rect 22661 31977 22695 32011
rect 22695 31977 22704 32011
rect 22652 31968 22704 31977
rect 24400 32011 24452 32020
rect 24400 31977 24409 32011
rect 24409 31977 24443 32011
rect 24443 31977 24452 32011
rect 24400 31968 24452 31977
rect 26332 31968 26384 32020
rect 23480 31875 23532 31884
rect 17592 31807 17644 31816
rect 17592 31773 17601 31807
rect 17601 31773 17635 31807
rect 17635 31773 17644 31807
rect 17592 31764 17644 31773
rect 16948 31628 17000 31680
rect 17132 31628 17184 31680
rect 17960 31628 18012 31680
rect 18328 31764 18380 31816
rect 22468 31764 22520 31816
rect 23480 31841 23489 31875
rect 23489 31841 23523 31875
rect 23523 31841 23532 31875
rect 23480 31832 23532 31841
rect 25044 31875 25096 31884
rect 25044 31841 25053 31875
rect 25053 31841 25087 31875
rect 25087 31841 25096 31875
rect 25044 31832 25096 31841
rect 23388 31807 23440 31816
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 23388 31764 23440 31773
rect 28816 31900 28868 31952
rect 29828 31968 29880 32020
rect 30288 31968 30340 32020
rect 32496 32011 32548 32020
rect 32496 31977 32505 32011
rect 32505 31977 32539 32011
rect 32539 31977 32548 32011
rect 32496 31968 32548 31977
rect 33048 32011 33100 32020
rect 33048 31977 33057 32011
rect 33057 31977 33091 32011
rect 33091 31977 33100 32011
rect 33048 31968 33100 31977
rect 48228 31968 48280 32020
rect 42708 31900 42760 31952
rect 26976 31875 27028 31884
rect 26976 31841 26985 31875
rect 26985 31841 27019 31875
rect 27019 31841 27028 31875
rect 26976 31832 27028 31841
rect 27252 31875 27304 31884
rect 27252 31841 27261 31875
rect 27261 31841 27295 31875
rect 27295 31841 27304 31875
rect 27252 31832 27304 31841
rect 27344 31832 27396 31884
rect 29000 31832 29052 31884
rect 25964 31764 26016 31816
rect 25688 31696 25740 31748
rect 28264 31764 28316 31816
rect 28632 31764 28684 31816
rect 32772 31832 32824 31884
rect 46756 31832 46808 31884
rect 47400 31875 47452 31884
rect 47400 31841 47409 31875
rect 47409 31841 47443 31875
rect 47443 31841 47452 31875
rect 47400 31832 47452 31841
rect 30012 31764 30064 31816
rect 30104 31807 30156 31816
rect 30104 31773 30113 31807
rect 30113 31773 30147 31807
rect 30147 31773 30156 31807
rect 30104 31764 30156 31773
rect 18144 31628 18196 31680
rect 18328 31671 18380 31680
rect 18328 31637 18337 31671
rect 18337 31637 18371 31671
rect 18371 31637 18380 31671
rect 18328 31628 18380 31637
rect 22008 31628 22060 31680
rect 25228 31628 25280 31680
rect 29368 31696 29420 31748
rect 26148 31628 26200 31680
rect 29000 31628 29052 31680
rect 30932 31807 30984 31816
rect 30932 31773 30941 31807
rect 30941 31773 30975 31807
rect 30975 31773 30984 31807
rect 30932 31764 30984 31773
rect 31760 31807 31812 31816
rect 31760 31773 31769 31807
rect 31769 31773 31803 31807
rect 31803 31773 31812 31807
rect 31760 31764 31812 31773
rect 31944 31807 31996 31816
rect 31944 31773 31953 31807
rect 31953 31773 31987 31807
rect 31987 31773 31996 31807
rect 31944 31764 31996 31773
rect 32128 31807 32180 31816
rect 32128 31773 32137 31807
rect 32137 31773 32171 31807
rect 32171 31773 32180 31807
rect 32128 31764 32180 31773
rect 32312 31807 32364 31816
rect 32312 31773 32321 31807
rect 32321 31773 32355 31807
rect 32355 31773 32364 31807
rect 32312 31764 32364 31773
rect 32864 31764 32916 31816
rect 46664 31739 46716 31748
rect 46664 31705 46673 31739
rect 46673 31705 46707 31739
rect 46707 31705 46716 31739
rect 46664 31696 46716 31705
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 17316 31424 17368 31476
rect 19340 31424 19392 31476
rect 21088 31424 21140 31476
rect 22468 31424 22520 31476
rect 18328 31356 18380 31408
rect 20352 31356 20404 31408
rect 21640 31356 21692 31408
rect 2044 31288 2096 31340
rect 2228 31288 2280 31340
rect 14464 31331 14516 31340
rect 14464 31297 14473 31331
rect 14473 31297 14507 31331
rect 14507 31297 14516 31331
rect 14464 31288 14516 31297
rect 14740 31220 14792 31272
rect 16856 31288 16908 31340
rect 17132 31331 17184 31340
rect 17132 31297 17141 31331
rect 17141 31297 17175 31331
rect 17175 31297 17184 31331
rect 17132 31288 17184 31297
rect 19340 31288 19392 31340
rect 20536 31331 20588 31340
rect 20536 31297 20545 31331
rect 20545 31297 20579 31331
rect 20579 31297 20588 31331
rect 20536 31288 20588 31297
rect 20720 31331 20772 31340
rect 20720 31297 20729 31331
rect 20729 31297 20763 31331
rect 20763 31297 20772 31331
rect 20720 31288 20772 31297
rect 21824 31288 21876 31340
rect 22560 31331 22612 31340
rect 17224 31220 17276 31272
rect 18052 31220 18104 31272
rect 20812 31263 20864 31272
rect 14924 31152 14976 31204
rect 20812 31229 20821 31263
rect 20821 31229 20855 31263
rect 20855 31229 20864 31263
rect 20812 31220 20864 31229
rect 21548 31220 21600 31272
rect 21180 31152 21232 31204
rect 22560 31297 22569 31331
rect 22569 31297 22603 31331
rect 22603 31297 22612 31331
rect 22560 31288 22612 31297
rect 22100 31195 22152 31204
rect 22100 31161 22109 31195
rect 22109 31161 22143 31195
rect 22143 31161 22152 31195
rect 22100 31152 22152 31161
rect 15292 31127 15344 31136
rect 15292 31093 15301 31127
rect 15301 31093 15335 31127
rect 15335 31093 15344 31127
rect 15292 31084 15344 31093
rect 17868 31084 17920 31136
rect 23756 31467 23808 31476
rect 23756 31433 23765 31467
rect 23765 31433 23799 31467
rect 23799 31433 23808 31467
rect 23756 31424 23808 31433
rect 24584 31467 24636 31476
rect 24584 31433 24593 31467
rect 24593 31433 24627 31467
rect 24627 31433 24636 31467
rect 24584 31424 24636 31433
rect 25044 31424 25096 31476
rect 27896 31467 27948 31476
rect 27896 31433 27905 31467
rect 27905 31433 27939 31467
rect 27939 31433 27948 31467
rect 27896 31424 27948 31433
rect 24216 31399 24268 31408
rect 24216 31365 24225 31399
rect 24225 31365 24259 31399
rect 24259 31365 24268 31399
rect 24216 31356 24268 31365
rect 25596 31356 25648 31408
rect 27528 31356 27580 31408
rect 25228 31288 25280 31340
rect 25964 31288 26016 31340
rect 27988 31288 28040 31340
rect 28448 31424 28500 31476
rect 28908 31424 28960 31476
rect 32312 31424 32364 31476
rect 30288 31356 30340 31408
rect 31944 31356 31996 31408
rect 28816 31288 28868 31340
rect 29000 31288 29052 31340
rect 29828 31288 29880 31340
rect 31116 31288 31168 31340
rect 23572 31127 23624 31136
rect 23572 31093 23581 31127
rect 23581 31093 23615 31127
rect 23615 31093 23624 31127
rect 23572 31084 23624 31093
rect 26332 31220 26384 31272
rect 28356 31263 28408 31272
rect 28356 31229 28365 31263
rect 28365 31229 28399 31263
rect 28399 31229 28408 31263
rect 28356 31220 28408 31229
rect 30104 31220 30156 31272
rect 30288 31220 30340 31272
rect 32404 31263 32456 31272
rect 32404 31229 32413 31263
rect 32413 31229 32447 31263
rect 32447 31229 32456 31263
rect 32404 31220 32456 31229
rect 40224 31220 40276 31272
rect 25228 31152 25280 31204
rect 30840 31152 30892 31204
rect 30012 31127 30064 31136
rect 30012 31093 30021 31127
rect 30021 31093 30055 31127
rect 30055 31093 30064 31127
rect 30012 31084 30064 31093
rect 30104 31127 30156 31136
rect 30104 31093 30113 31127
rect 30113 31093 30147 31127
rect 30147 31093 30156 31127
rect 30104 31084 30156 31093
rect 32220 31084 32272 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 17132 30880 17184 30932
rect 17868 30923 17920 30932
rect 17868 30889 17877 30923
rect 17877 30889 17911 30923
rect 17911 30889 17920 30923
rect 17868 30880 17920 30889
rect 19340 30923 19392 30932
rect 19340 30889 19349 30923
rect 19349 30889 19383 30923
rect 19383 30889 19392 30923
rect 19340 30880 19392 30889
rect 20812 30880 20864 30932
rect 23112 30880 23164 30932
rect 25228 30880 25280 30932
rect 17224 30812 17276 30864
rect 20720 30812 20772 30864
rect 25136 30812 25188 30864
rect 20996 30744 21048 30796
rect 23572 30744 23624 30796
rect 26240 30880 26292 30932
rect 27436 30923 27488 30932
rect 27436 30889 27445 30923
rect 27445 30889 27479 30923
rect 27479 30889 27488 30923
rect 27436 30880 27488 30889
rect 29552 30880 29604 30932
rect 30748 30923 30800 30932
rect 30748 30889 30757 30923
rect 30757 30889 30791 30923
rect 30791 30889 30800 30923
rect 30748 30880 30800 30889
rect 31116 30923 31168 30932
rect 31116 30889 31125 30923
rect 31125 30889 31159 30923
rect 31159 30889 31168 30923
rect 31116 30880 31168 30889
rect 29920 30812 29972 30864
rect 16948 30676 17000 30728
rect 15844 30608 15896 30660
rect 17316 30676 17368 30728
rect 19248 30719 19300 30728
rect 17776 30608 17828 30660
rect 19248 30685 19257 30719
rect 19257 30685 19291 30719
rect 19291 30685 19300 30719
rect 19248 30676 19300 30685
rect 22008 30676 22060 30728
rect 22284 30676 22336 30728
rect 25596 30676 25648 30728
rect 26608 30744 26660 30796
rect 30104 30744 30156 30796
rect 30840 30787 30892 30796
rect 30840 30753 30849 30787
rect 30849 30753 30883 30787
rect 30883 30753 30892 30787
rect 30840 30744 30892 30753
rect 32220 30787 32272 30796
rect 32220 30753 32229 30787
rect 32229 30753 32263 30787
rect 32263 30753 32272 30787
rect 32220 30744 32272 30753
rect 20076 30608 20128 30660
rect 23296 30608 23348 30660
rect 25688 30608 25740 30660
rect 26976 30608 27028 30660
rect 30012 30676 30064 30728
rect 30932 30676 30984 30728
rect 29184 30608 29236 30660
rect 33232 30608 33284 30660
rect 15476 30540 15528 30592
rect 17408 30583 17460 30592
rect 17408 30549 17417 30583
rect 17417 30549 17451 30583
rect 17451 30549 17460 30583
rect 17408 30540 17460 30549
rect 25136 30540 25188 30592
rect 26056 30540 26108 30592
rect 26608 30540 26660 30592
rect 26792 30583 26844 30592
rect 26792 30549 26801 30583
rect 26801 30549 26835 30583
rect 26835 30549 26844 30583
rect 26792 30540 26844 30549
rect 29000 30540 29052 30592
rect 32404 30540 32456 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 15292 30336 15344 30388
rect 15476 30379 15528 30388
rect 15476 30345 15485 30379
rect 15485 30345 15519 30379
rect 15519 30345 15528 30379
rect 15476 30336 15528 30345
rect 16856 30336 16908 30388
rect 19340 30336 19392 30388
rect 25136 30379 25188 30388
rect 15844 30268 15896 30320
rect 14924 30243 14976 30252
rect 14924 30209 14934 30243
rect 14934 30209 14968 30243
rect 14968 30209 14976 30243
rect 14924 30200 14976 30209
rect 15200 30243 15252 30252
rect 15200 30209 15209 30243
rect 15209 30209 15243 30243
rect 15243 30209 15252 30243
rect 15200 30200 15252 30209
rect 15936 30243 15988 30252
rect 15936 30209 15945 30243
rect 15945 30209 15979 30243
rect 15979 30209 15988 30243
rect 23756 30268 23808 30320
rect 15936 30200 15988 30209
rect 16120 30132 16172 30184
rect 17408 30200 17460 30252
rect 17868 30200 17920 30252
rect 19432 30200 19484 30252
rect 20812 30200 20864 30252
rect 20996 30200 21048 30252
rect 22284 30200 22336 30252
rect 24860 30268 24912 30320
rect 25136 30345 25145 30379
rect 25145 30345 25179 30379
rect 25179 30345 25188 30379
rect 25136 30336 25188 30345
rect 25688 30336 25740 30388
rect 29000 30336 29052 30388
rect 30288 30336 30340 30388
rect 24400 30200 24452 30252
rect 27528 30268 27580 30320
rect 30656 30268 30708 30320
rect 33232 30268 33284 30320
rect 25872 30200 25924 30252
rect 28632 30243 28684 30252
rect 28632 30209 28641 30243
rect 28641 30209 28675 30243
rect 28675 30209 28684 30243
rect 28632 30200 28684 30209
rect 32864 30243 32916 30252
rect 32864 30209 32873 30243
rect 32873 30209 32907 30243
rect 32907 30209 32916 30243
rect 32864 30200 32916 30209
rect 16856 30064 16908 30116
rect 18236 30064 18288 30116
rect 19340 30064 19392 30116
rect 21640 30064 21692 30116
rect 23756 30064 23808 30116
rect 24492 30132 24544 30184
rect 25136 30132 25188 30184
rect 28540 30132 28592 30184
rect 29000 30132 29052 30184
rect 34336 30175 34388 30184
rect 16672 29996 16724 30048
rect 20720 29996 20772 30048
rect 25964 30064 26016 30116
rect 27252 30107 27304 30116
rect 27252 30073 27261 30107
rect 27261 30073 27295 30107
rect 27295 30073 27304 30107
rect 34336 30141 34345 30175
rect 34345 30141 34379 30175
rect 34379 30141 34388 30175
rect 34336 30132 34388 30141
rect 34796 30132 34848 30184
rect 34888 30175 34940 30184
rect 34888 30141 34897 30175
rect 34897 30141 34931 30175
rect 34931 30141 34940 30175
rect 34888 30132 34940 30141
rect 27252 30064 27304 30073
rect 24492 30039 24544 30048
rect 24492 30005 24501 30039
rect 24501 30005 24535 30039
rect 24535 30005 24544 30039
rect 24492 29996 24544 30005
rect 28172 29996 28224 30048
rect 29828 29996 29880 30048
rect 30932 29996 30984 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 17776 29792 17828 29844
rect 20812 29792 20864 29844
rect 20996 29792 21048 29844
rect 21916 29835 21968 29844
rect 21916 29801 21925 29835
rect 21925 29801 21959 29835
rect 21959 29801 21968 29835
rect 21916 29792 21968 29801
rect 22652 29792 22704 29844
rect 22836 29792 22888 29844
rect 25136 29792 25188 29844
rect 21640 29724 21692 29776
rect 28632 29792 28684 29844
rect 30656 29835 30708 29844
rect 30656 29801 30665 29835
rect 30665 29801 30699 29835
rect 30699 29801 30708 29835
rect 30656 29792 30708 29801
rect 34796 29835 34848 29844
rect 34796 29801 34805 29835
rect 34805 29801 34839 29835
rect 34839 29801 34848 29835
rect 34796 29792 34848 29801
rect 27988 29724 28040 29776
rect 29000 29724 29052 29776
rect 29460 29724 29512 29776
rect 30012 29724 30064 29776
rect 17132 29656 17184 29708
rect 19248 29588 19300 29640
rect 21180 29656 21232 29708
rect 22652 29656 22704 29708
rect 27252 29656 27304 29708
rect 29552 29656 29604 29708
rect 16396 29563 16448 29572
rect 16396 29529 16405 29563
rect 16405 29529 16439 29563
rect 16439 29529 16448 29563
rect 16396 29520 16448 29529
rect 21272 29588 21324 29640
rect 21824 29588 21876 29640
rect 22008 29631 22060 29640
rect 22008 29597 22017 29631
rect 22017 29597 22051 29631
rect 22051 29597 22060 29631
rect 22008 29588 22060 29597
rect 22560 29588 22612 29640
rect 24492 29588 24544 29640
rect 29920 29656 29972 29708
rect 30012 29631 30064 29640
rect 21640 29520 21692 29572
rect 26332 29520 26384 29572
rect 27068 29520 27120 29572
rect 30012 29597 30021 29631
rect 30021 29597 30055 29631
rect 30055 29597 30064 29631
rect 30012 29588 30064 29597
rect 30564 29631 30616 29640
rect 30564 29597 30573 29631
rect 30573 29597 30607 29631
rect 30607 29597 30616 29631
rect 30564 29588 30616 29597
rect 32864 29588 32916 29640
rect 35348 29588 35400 29640
rect 47216 29656 47268 29708
rect 47400 29588 47452 29640
rect 43904 29520 43956 29572
rect 15200 29452 15252 29504
rect 17132 29452 17184 29504
rect 20076 29452 20128 29504
rect 20260 29495 20312 29504
rect 20260 29461 20269 29495
rect 20269 29461 20303 29495
rect 20303 29461 20312 29495
rect 20260 29452 20312 29461
rect 21732 29452 21784 29504
rect 23020 29495 23072 29504
rect 23020 29461 23029 29495
rect 23029 29461 23063 29495
rect 23063 29461 23072 29495
rect 23020 29452 23072 29461
rect 23112 29452 23164 29504
rect 23848 29452 23900 29504
rect 25688 29452 25740 29504
rect 26792 29452 26844 29504
rect 26884 29452 26936 29504
rect 28172 29452 28224 29504
rect 30564 29452 30616 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 16396 29248 16448 29300
rect 21272 29291 21324 29300
rect 21272 29257 21281 29291
rect 21281 29257 21315 29291
rect 21315 29257 21324 29291
rect 21272 29248 21324 29257
rect 21916 29248 21968 29300
rect 22928 29248 22980 29300
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 17776 29180 17828 29232
rect 20260 29180 20312 29232
rect 21640 29180 21692 29232
rect 23020 29180 23072 29232
rect 26332 29248 26384 29300
rect 27068 29291 27120 29300
rect 27068 29257 27077 29291
rect 27077 29257 27111 29291
rect 27111 29257 27120 29291
rect 27068 29248 27120 29257
rect 26516 29180 26568 29232
rect 16856 29112 16908 29164
rect 17500 29112 17552 29164
rect 21548 29112 21600 29164
rect 22652 29155 22704 29164
rect 22652 29121 22661 29155
rect 22661 29121 22695 29155
rect 22695 29121 22704 29155
rect 22652 29112 22704 29121
rect 25136 29112 25188 29164
rect 25688 29112 25740 29164
rect 19800 29087 19852 29096
rect 17132 28976 17184 29028
rect 17224 28976 17276 29028
rect 19800 29053 19809 29087
rect 19809 29053 19843 29087
rect 19843 29053 19852 29087
rect 19800 29044 19852 29053
rect 22928 29087 22980 29096
rect 22928 29053 22937 29087
rect 22937 29053 22971 29087
rect 22971 29053 22980 29087
rect 22928 29044 22980 29053
rect 23296 29044 23348 29096
rect 25596 29044 25648 29096
rect 26056 29155 26108 29164
rect 26056 29121 26065 29155
rect 26065 29121 26099 29155
rect 26099 29121 26108 29155
rect 26056 29112 26108 29121
rect 26424 29112 26476 29164
rect 26976 29155 27028 29164
rect 26976 29121 26985 29155
rect 26985 29121 27019 29155
rect 27019 29121 27028 29155
rect 26976 29112 27028 29121
rect 29184 29112 29236 29164
rect 26884 29044 26936 29096
rect 32680 29087 32732 29096
rect 32680 29053 32689 29087
rect 32689 29053 32723 29087
rect 32723 29053 32732 29087
rect 32680 29044 32732 29053
rect 32864 29087 32916 29096
rect 32864 29053 32873 29087
rect 32873 29053 32907 29087
rect 32907 29053 32916 29087
rect 32864 29044 32916 29053
rect 33140 29087 33192 29096
rect 33140 29053 33149 29087
rect 33149 29053 33183 29087
rect 33183 29053 33192 29087
rect 33140 29044 33192 29053
rect 25136 28908 25188 28960
rect 29552 28908 29604 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19800 28704 19852 28756
rect 21732 28747 21784 28756
rect 21732 28713 21741 28747
rect 21741 28713 21775 28747
rect 21775 28713 21784 28747
rect 21732 28704 21784 28713
rect 22652 28704 22704 28756
rect 22928 28704 22980 28756
rect 30196 28747 30248 28756
rect 15016 28568 15068 28620
rect 21272 28636 21324 28688
rect 18236 28568 18288 28620
rect 17960 28500 18012 28552
rect 20352 28543 20404 28552
rect 20352 28509 20361 28543
rect 20361 28509 20395 28543
rect 20395 28509 20404 28543
rect 20352 28500 20404 28509
rect 20536 28543 20588 28552
rect 20536 28509 20543 28543
rect 20543 28509 20588 28543
rect 20536 28500 20588 28509
rect 20076 28432 20128 28484
rect 26056 28636 26108 28688
rect 29552 28636 29604 28688
rect 30196 28713 30205 28747
rect 30205 28713 30239 28747
rect 30239 28713 30248 28747
rect 30196 28704 30248 28713
rect 30748 28704 30800 28756
rect 32864 28747 32916 28756
rect 32864 28713 32873 28747
rect 32873 28713 32907 28747
rect 32907 28713 32916 28747
rect 32864 28704 32916 28713
rect 34336 28704 34388 28756
rect 21824 28568 21876 28620
rect 23296 28568 23348 28620
rect 29460 28568 29512 28620
rect 30288 28568 30340 28620
rect 22652 28543 22704 28552
rect 17592 28364 17644 28416
rect 17776 28407 17828 28416
rect 17776 28373 17785 28407
rect 17785 28373 17819 28407
rect 17819 28373 17828 28407
rect 17776 28364 17828 28373
rect 19984 28364 20036 28416
rect 21640 28364 21692 28416
rect 22652 28509 22661 28543
rect 22661 28509 22695 28543
rect 22695 28509 22704 28543
rect 22652 28500 22704 28509
rect 22836 28543 22888 28552
rect 22836 28509 22845 28543
rect 22845 28509 22879 28543
rect 22879 28509 22888 28543
rect 22836 28500 22888 28509
rect 23020 28543 23072 28552
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 23204 28543 23256 28552
rect 23204 28509 23213 28543
rect 23213 28509 23247 28543
rect 23247 28509 23256 28543
rect 23204 28500 23256 28509
rect 29736 28475 29788 28484
rect 29736 28441 29745 28475
rect 29745 28441 29779 28475
rect 29779 28441 29788 28475
rect 29736 28432 29788 28441
rect 31668 28500 31720 28552
rect 36176 28568 36228 28620
rect 33692 28500 33744 28552
rect 46940 28500 46992 28552
rect 32404 28432 32456 28484
rect 34980 28475 35032 28484
rect 34980 28441 34989 28475
rect 34989 28441 35023 28475
rect 35023 28441 35032 28475
rect 34980 28432 35032 28441
rect 35440 28432 35492 28484
rect 23848 28364 23900 28416
rect 29000 28364 29052 28416
rect 29368 28364 29420 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1492 28160 1544 28212
rect 20352 28160 20404 28212
rect 17592 28067 17644 28076
rect 17592 28033 17601 28067
rect 17601 28033 17635 28067
rect 17635 28033 17644 28067
rect 17592 28024 17644 28033
rect 17776 28067 17828 28076
rect 17776 28033 17783 28067
rect 17783 28033 17828 28067
rect 17776 28024 17828 28033
rect 17960 28067 18012 28076
rect 17960 28033 17969 28067
rect 17969 28033 18003 28067
rect 18003 28033 18012 28067
rect 17960 28024 18012 28033
rect 18236 28024 18288 28076
rect 20076 28067 20128 28076
rect 20076 28033 20085 28067
rect 20085 28033 20119 28067
rect 20119 28033 20128 28067
rect 20076 28024 20128 28033
rect 20444 28024 20496 28076
rect 21640 28024 21692 28076
rect 21916 28067 21968 28076
rect 21916 28033 21925 28067
rect 21925 28033 21959 28067
rect 21959 28033 21968 28067
rect 21916 28024 21968 28033
rect 19984 27956 20036 28008
rect 24676 28160 24728 28212
rect 26516 28160 26568 28212
rect 25044 28092 25096 28144
rect 29000 28160 29052 28212
rect 29368 28160 29420 28212
rect 29644 28160 29696 28212
rect 33692 28203 33744 28212
rect 33692 28169 33701 28203
rect 33701 28169 33735 28203
rect 33735 28169 33744 28203
rect 33692 28160 33744 28169
rect 35440 28160 35492 28212
rect 42800 28160 42852 28212
rect 46848 28160 46900 28212
rect 23664 28024 23716 28076
rect 18236 27863 18288 27872
rect 18236 27829 18245 27863
rect 18245 27829 18279 27863
rect 18279 27829 18288 27863
rect 18236 27820 18288 27829
rect 21824 27863 21876 27872
rect 21824 27829 21833 27863
rect 21833 27829 21867 27863
rect 21867 27829 21876 27863
rect 21824 27820 21876 27829
rect 21916 27820 21968 27872
rect 23204 27888 23256 27940
rect 24584 27888 24636 27940
rect 26608 27956 26660 28008
rect 28080 27956 28132 28008
rect 29552 27956 29604 28008
rect 29368 27888 29420 27940
rect 31668 28024 31720 28076
rect 32496 28024 32548 28076
rect 34336 28024 34388 28076
rect 35532 28024 35584 28076
rect 47032 28024 47084 28076
rect 47400 28024 47452 28076
rect 30288 27956 30340 28008
rect 34704 27956 34756 28008
rect 34980 27956 35032 28008
rect 25136 27820 25188 27872
rect 26884 27820 26936 27872
rect 30380 27820 30432 27872
rect 30748 27863 30800 27872
rect 30748 27829 30757 27863
rect 30757 27829 30791 27863
rect 30791 27829 30800 27863
rect 30748 27820 30800 27829
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3516 27616 3568 27668
rect 31668 27659 31720 27668
rect 7472 27480 7524 27532
rect 31668 27625 31677 27659
rect 31677 27625 31711 27659
rect 31711 27625 31720 27659
rect 31668 27616 31720 27625
rect 15108 27548 15160 27600
rect 17868 27548 17920 27600
rect 15108 27455 15160 27464
rect 15108 27421 15117 27455
rect 15117 27421 15151 27455
rect 15151 27421 15160 27455
rect 15108 27412 15160 27421
rect 19984 27412 20036 27464
rect 22836 27548 22888 27600
rect 26056 27548 26108 27600
rect 15384 27344 15436 27396
rect 23204 27480 23256 27532
rect 21088 27455 21140 27464
rect 21088 27421 21097 27455
rect 21097 27421 21131 27455
rect 21131 27421 21140 27455
rect 21088 27412 21140 27421
rect 21272 27455 21324 27464
rect 21272 27421 21281 27455
rect 21281 27421 21315 27455
rect 21315 27421 21324 27455
rect 21272 27412 21324 27421
rect 20812 27344 20864 27396
rect 23848 27344 23900 27396
rect 25044 27412 25096 27464
rect 27896 27412 27948 27464
rect 28080 27455 28132 27464
rect 28080 27421 28089 27455
rect 28089 27421 28123 27455
rect 28123 27421 28132 27455
rect 28080 27412 28132 27421
rect 29460 27548 29512 27600
rect 29828 27480 29880 27532
rect 46940 27548 46992 27600
rect 47676 27480 47728 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 25228 27344 25280 27396
rect 26608 27344 26660 27396
rect 32496 27455 32548 27464
rect 32496 27421 32505 27455
rect 32505 27421 32539 27455
rect 32539 27421 32548 27455
rect 32496 27412 32548 27421
rect 35532 27412 35584 27464
rect 20628 27319 20680 27328
rect 20628 27285 20637 27319
rect 20637 27285 20671 27319
rect 20671 27285 20680 27319
rect 20628 27276 20680 27285
rect 21180 27319 21232 27328
rect 21180 27285 21189 27319
rect 21189 27285 21223 27319
rect 21223 27285 21232 27319
rect 21180 27276 21232 27285
rect 24768 27319 24820 27328
rect 24768 27285 24777 27319
rect 24777 27285 24811 27319
rect 24811 27285 24820 27319
rect 24768 27276 24820 27285
rect 27528 27319 27580 27328
rect 27528 27285 27537 27319
rect 27537 27285 27571 27319
rect 27571 27285 27580 27319
rect 27528 27276 27580 27285
rect 27988 27276 28040 27328
rect 30196 27387 30248 27396
rect 30196 27353 30205 27387
rect 30205 27353 30239 27387
rect 30239 27353 30248 27387
rect 30196 27344 30248 27353
rect 31208 27344 31260 27396
rect 28816 27319 28868 27328
rect 28816 27285 28831 27319
rect 28831 27285 28865 27319
rect 28865 27285 28868 27319
rect 28816 27276 28868 27285
rect 30288 27276 30340 27328
rect 32312 27276 32364 27328
rect 33324 27276 33376 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 15384 27115 15436 27124
rect 15384 27081 15393 27115
rect 15393 27081 15427 27115
rect 15427 27081 15436 27115
rect 15384 27072 15436 27081
rect 22008 27072 22060 27124
rect 28080 27072 28132 27124
rect 30196 27115 30248 27124
rect 15476 26936 15528 26988
rect 18604 26936 18656 26988
rect 21916 27004 21968 27056
rect 17224 26911 17276 26920
rect 17224 26877 17233 26911
rect 17233 26877 17267 26911
rect 17267 26877 17276 26911
rect 17224 26868 17276 26877
rect 18236 26868 18288 26920
rect 20076 26868 20128 26920
rect 20812 26979 20864 26988
rect 20812 26945 20821 26979
rect 20821 26945 20855 26979
rect 20855 26945 20864 26979
rect 20812 26936 20864 26945
rect 21548 26936 21600 26988
rect 21732 26936 21784 26988
rect 21088 26868 21140 26920
rect 21640 26868 21692 26920
rect 23756 26936 23808 26988
rect 23848 26979 23900 26988
rect 23848 26945 23857 26979
rect 23857 26945 23891 26979
rect 23891 26945 23900 26979
rect 27252 27004 27304 27056
rect 27528 27004 27580 27056
rect 30196 27081 30205 27115
rect 30205 27081 30239 27115
rect 30239 27081 30248 27115
rect 30196 27072 30248 27081
rect 31208 27115 31260 27124
rect 31208 27081 31217 27115
rect 31217 27081 31251 27115
rect 31251 27081 31260 27115
rect 31208 27072 31260 27081
rect 32680 27072 32732 27124
rect 34336 27072 34388 27124
rect 29736 27004 29788 27056
rect 31392 27004 31444 27056
rect 33324 27004 33376 27056
rect 33968 27004 34020 27056
rect 35808 27072 35860 27124
rect 34612 27004 34664 27056
rect 23848 26936 23900 26945
rect 29460 26979 29512 26988
rect 23388 26868 23440 26920
rect 29460 26945 29469 26979
rect 29469 26945 29503 26979
rect 29503 26945 29512 26979
rect 29460 26936 29512 26945
rect 30380 26979 30432 26988
rect 30380 26945 30389 26979
rect 30389 26945 30423 26979
rect 30423 26945 30432 26979
rect 30380 26936 30432 26945
rect 30748 26936 30800 26988
rect 32312 26979 32364 26988
rect 24860 26868 24912 26920
rect 26884 26868 26936 26920
rect 30288 26868 30340 26920
rect 15016 26732 15068 26784
rect 17960 26732 18012 26784
rect 21548 26800 21600 26852
rect 21272 26732 21324 26784
rect 22008 26732 22060 26784
rect 23480 26732 23532 26784
rect 24860 26775 24912 26784
rect 24860 26741 24869 26775
rect 24869 26741 24903 26775
rect 24903 26741 24912 26775
rect 24860 26732 24912 26741
rect 27896 26732 27948 26784
rect 32312 26945 32321 26979
rect 32321 26945 32355 26979
rect 32355 26945 32364 26979
rect 32312 26936 32364 26945
rect 33876 26936 33928 26988
rect 33140 26868 33192 26920
rect 34612 26800 34664 26852
rect 34796 26732 34848 26784
rect 35348 26775 35400 26784
rect 35348 26741 35357 26775
rect 35357 26741 35391 26775
rect 35391 26741 35400 26775
rect 35348 26732 35400 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 18604 26571 18656 26580
rect 18604 26537 18613 26571
rect 18613 26537 18647 26571
rect 18647 26537 18656 26571
rect 18604 26528 18656 26537
rect 20628 26528 20680 26580
rect 20812 26528 20864 26580
rect 21916 26528 21968 26580
rect 21180 26460 21232 26512
rect 15016 26435 15068 26444
rect 15016 26401 15025 26435
rect 15025 26401 15059 26435
rect 15059 26401 15068 26435
rect 15016 26392 15068 26401
rect 16488 26435 16540 26444
rect 16488 26401 16497 26435
rect 16497 26401 16531 26435
rect 16531 26401 16540 26435
rect 16488 26392 16540 26401
rect 17224 26392 17276 26444
rect 21640 26435 21692 26444
rect 13728 26324 13780 26376
rect 21640 26401 21649 26435
rect 21649 26401 21683 26435
rect 21683 26401 21692 26435
rect 21640 26392 21692 26401
rect 22284 26460 22336 26512
rect 23388 26460 23440 26512
rect 19248 26256 19300 26308
rect 19984 26256 20036 26308
rect 21548 26299 21600 26308
rect 21548 26265 21557 26299
rect 21557 26265 21591 26299
rect 21591 26265 21600 26299
rect 21548 26256 21600 26265
rect 22192 26324 22244 26376
rect 23480 26367 23532 26376
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 23664 26460 23716 26512
rect 23756 26460 23808 26512
rect 24400 26435 24452 26444
rect 24400 26401 24409 26435
rect 24409 26401 24443 26435
rect 24443 26401 24452 26435
rect 24400 26392 24452 26401
rect 23756 26324 23808 26376
rect 28632 26528 28684 26580
rect 33140 26571 33192 26580
rect 26608 26503 26660 26512
rect 24676 26435 24728 26444
rect 24676 26401 24685 26435
rect 24685 26401 24719 26435
rect 24719 26401 24728 26435
rect 24676 26392 24728 26401
rect 24768 26392 24820 26444
rect 26240 26324 26292 26376
rect 26608 26469 26617 26503
rect 26617 26469 26651 26503
rect 26651 26469 26660 26503
rect 33140 26537 33149 26571
rect 33149 26537 33183 26571
rect 33183 26537 33192 26571
rect 33140 26528 33192 26537
rect 33876 26571 33928 26580
rect 33876 26537 33885 26571
rect 33885 26537 33919 26571
rect 33919 26537 33928 26571
rect 33876 26528 33928 26537
rect 26608 26460 26660 26469
rect 29184 26324 29236 26376
rect 25964 26256 26016 26308
rect 27436 26256 27488 26308
rect 28632 26299 28684 26308
rect 28632 26265 28641 26299
rect 28641 26265 28675 26299
rect 28675 26265 28684 26299
rect 28632 26256 28684 26265
rect 28816 26299 28868 26308
rect 28816 26265 28825 26299
rect 28825 26265 28859 26299
rect 28859 26265 28868 26299
rect 28816 26256 28868 26265
rect 22100 26188 22152 26240
rect 23848 26188 23900 26240
rect 25136 26188 25188 26240
rect 27988 26231 28040 26240
rect 27988 26197 27997 26231
rect 27997 26197 28031 26231
rect 28031 26197 28040 26231
rect 27988 26188 28040 26197
rect 29460 26324 29512 26376
rect 34612 26392 34664 26444
rect 35348 26392 35400 26444
rect 35992 26392 36044 26444
rect 42800 26392 42852 26444
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 32680 26324 32732 26376
rect 33968 26324 34020 26376
rect 34428 26324 34480 26376
rect 36912 26324 36964 26376
rect 34612 26256 34664 26308
rect 35992 26256 36044 26308
rect 37648 26299 37700 26308
rect 37648 26265 37657 26299
rect 37657 26265 37691 26299
rect 37691 26265 37700 26299
rect 37648 26256 37700 26265
rect 34888 26188 34940 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 19984 25984 20036 26036
rect 20168 25984 20220 26036
rect 24400 25984 24452 26036
rect 29460 25984 29512 26036
rect 34428 25984 34480 26036
rect 34796 25984 34848 26036
rect 35992 25984 36044 26036
rect 23572 25916 23624 25968
rect 24860 25916 24912 25968
rect 19248 25891 19300 25900
rect 19248 25857 19257 25891
rect 19257 25857 19291 25891
rect 19291 25857 19300 25891
rect 19248 25848 19300 25857
rect 19340 25848 19392 25900
rect 21180 25848 21232 25900
rect 22100 25848 22152 25900
rect 24768 25891 24820 25900
rect 24768 25857 24777 25891
rect 24777 25857 24811 25891
rect 24811 25857 24820 25891
rect 24768 25848 24820 25857
rect 12348 25823 12400 25832
rect 12348 25789 12357 25823
rect 12357 25789 12391 25823
rect 12391 25789 12400 25823
rect 12348 25780 12400 25789
rect 14280 25780 14332 25832
rect 16856 25823 16908 25832
rect 16856 25789 16865 25823
rect 16865 25789 16899 25823
rect 16899 25789 16908 25823
rect 16856 25780 16908 25789
rect 12808 25712 12860 25764
rect 16764 25712 16816 25764
rect 23296 25780 23348 25832
rect 24124 25780 24176 25832
rect 26516 25916 26568 25968
rect 27988 25916 28040 25968
rect 29644 25916 29696 25968
rect 34336 25959 34388 25968
rect 34336 25925 34345 25959
rect 34345 25925 34379 25959
rect 34379 25925 34388 25959
rect 34336 25916 34388 25925
rect 35808 25916 35860 25968
rect 25320 25848 25372 25900
rect 27252 25848 27304 25900
rect 27344 25780 27396 25832
rect 32496 25780 32548 25832
rect 34704 25891 34756 25900
rect 34704 25857 34713 25891
rect 34713 25857 34747 25891
rect 34747 25857 34756 25891
rect 34704 25848 34756 25857
rect 35532 25848 35584 25900
rect 44916 25891 44968 25900
rect 34796 25780 34848 25832
rect 34520 25712 34572 25764
rect 44916 25857 44925 25891
rect 44925 25857 44959 25891
rect 44959 25857 44968 25891
rect 44916 25848 44968 25857
rect 20076 25687 20128 25696
rect 20076 25653 20085 25687
rect 20085 25653 20119 25687
rect 20119 25653 20128 25687
rect 20076 25644 20128 25653
rect 25044 25644 25096 25696
rect 45468 25644 45520 25696
rect 46204 25644 46256 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 12348 25440 12400 25492
rect 19432 25483 19484 25492
rect 19432 25449 19441 25483
rect 19441 25449 19475 25483
rect 19475 25449 19484 25483
rect 19432 25440 19484 25449
rect 21548 25440 21600 25492
rect 21916 25440 21968 25492
rect 23296 25483 23348 25492
rect 23296 25449 23305 25483
rect 23305 25449 23339 25483
rect 23339 25449 23348 25483
rect 23296 25440 23348 25449
rect 19248 25372 19300 25424
rect 23664 25372 23716 25424
rect 8300 25304 8352 25356
rect 21640 25304 21692 25356
rect 25136 25440 25188 25492
rect 25228 25440 25280 25492
rect 29644 25483 29696 25492
rect 29644 25449 29653 25483
rect 29653 25449 29687 25483
rect 29687 25449 29696 25483
rect 29644 25440 29696 25449
rect 34520 25440 34572 25492
rect 37648 25440 37700 25492
rect 37188 25372 37240 25424
rect 45836 25372 45888 25424
rect 12256 25236 12308 25288
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 13728 25236 13780 25288
rect 13912 25236 13964 25288
rect 15292 25236 15344 25288
rect 16028 25236 16080 25288
rect 18144 25236 18196 25288
rect 20536 25236 20588 25288
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 23480 25279 23532 25288
rect 23480 25245 23489 25279
rect 23489 25245 23523 25279
rect 23523 25245 23532 25279
rect 23480 25236 23532 25245
rect 27252 25304 27304 25356
rect 36084 25304 36136 25356
rect 41788 25347 41840 25356
rect 41788 25313 41797 25347
rect 41797 25313 41831 25347
rect 41831 25313 41840 25347
rect 41788 25304 41840 25313
rect 45468 25347 45520 25356
rect 45468 25313 45477 25347
rect 45477 25313 45511 25347
rect 45511 25313 45520 25347
rect 45468 25304 45520 25313
rect 46848 25347 46900 25356
rect 46848 25313 46857 25347
rect 46857 25313 46891 25347
rect 46891 25313 46900 25347
rect 46848 25304 46900 25313
rect 13360 25168 13412 25220
rect 17408 25168 17460 25220
rect 23848 25279 23900 25288
rect 23848 25245 23857 25279
rect 23857 25245 23891 25279
rect 23891 25245 23900 25279
rect 23848 25236 23900 25245
rect 27896 25236 27948 25288
rect 28908 25236 28960 25288
rect 29736 25236 29788 25288
rect 35900 25236 35952 25288
rect 36176 25236 36228 25288
rect 37188 25279 37240 25288
rect 37188 25245 37197 25279
rect 37197 25245 37231 25279
rect 37231 25245 37240 25279
rect 37188 25236 37240 25245
rect 37832 25279 37884 25288
rect 37832 25245 37841 25279
rect 37841 25245 37875 25279
rect 37875 25245 37884 25279
rect 37832 25236 37884 25245
rect 45008 25236 45060 25288
rect 47768 25279 47820 25288
rect 47768 25245 47777 25279
rect 47777 25245 47811 25279
rect 47811 25245 47820 25279
rect 47768 25236 47820 25245
rect 24124 25168 24176 25220
rect 25044 25211 25096 25220
rect 25044 25177 25053 25211
rect 25053 25177 25087 25211
rect 25087 25177 25096 25211
rect 25044 25168 25096 25177
rect 25596 25168 25648 25220
rect 40132 25211 40184 25220
rect 40132 25177 40141 25211
rect 40141 25177 40175 25211
rect 40175 25177 40184 25211
rect 40132 25168 40184 25177
rect 2136 25143 2188 25152
rect 2136 25109 2145 25143
rect 2145 25109 2179 25143
rect 2179 25109 2188 25143
rect 2136 25100 2188 25109
rect 12532 25100 12584 25152
rect 14188 25143 14240 25152
rect 14188 25109 14197 25143
rect 14197 25109 14231 25143
rect 14231 25109 14240 25143
rect 14188 25100 14240 25109
rect 22376 25100 22428 25152
rect 27528 25100 27580 25152
rect 37464 25100 37516 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 2136 24896 2188 24948
rect 12808 24871 12860 24880
rect 12808 24837 12817 24871
rect 12817 24837 12851 24871
rect 12851 24837 12860 24871
rect 12808 24828 12860 24837
rect 14188 24828 14240 24880
rect 25872 24896 25924 24948
rect 27804 24896 27856 24948
rect 27896 24896 27948 24948
rect 40132 24939 40184 24948
rect 40132 24905 40141 24939
rect 40141 24905 40175 24939
rect 40175 24905 40184 24939
rect 40132 24896 40184 24905
rect 12256 24760 12308 24812
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 14096 24760 14148 24812
rect 15660 24760 15712 24812
rect 15752 24803 15804 24812
rect 15752 24769 15761 24803
rect 15761 24769 15795 24803
rect 15795 24769 15804 24803
rect 15752 24760 15804 24769
rect 17132 24760 17184 24812
rect 17316 24803 17368 24812
rect 17316 24769 17325 24803
rect 17325 24769 17359 24803
rect 17359 24769 17368 24803
rect 17316 24760 17368 24769
rect 17408 24803 17460 24812
rect 17408 24769 17417 24803
rect 17417 24769 17451 24803
rect 17451 24769 17460 24803
rect 18144 24803 18196 24812
rect 17408 24760 17460 24769
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 19340 24803 19392 24812
rect 19340 24769 19349 24803
rect 19349 24769 19383 24803
rect 19383 24769 19392 24803
rect 19340 24760 19392 24769
rect 14280 24735 14332 24744
rect 14280 24701 14289 24735
rect 14289 24701 14323 24735
rect 14323 24701 14332 24735
rect 14280 24692 14332 24701
rect 14832 24735 14884 24744
rect 14832 24701 14841 24735
rect 14841 24701 14875 24735
rect 14875 24701 14884 24735
rect 14832 24692 14884 24701
rect 15292 24735 15344 24744
rect 15292 24701 15301 24735
rect 15301 24701 15335 24735
rect 15335 24701 15344 24735
rect 15292 24692 15344 24701
rect 15936 24692 15988 24744
rect 20996 24692 21048 24744
rect 23572 24803 23624 24812
rect 23572 24769 23581 24803
rect 23581 24769 23615 24803
rect 23615 24769 23624 24803
rect 23572 24760 23624 24769
rect 23664 24692 23716 24744
rect 24768 24692 24820 24744
rect 25596 24803 25648 24812
rect 25596 24769 25605 24803
rect 25605 24769 25639 24803
rect 25639 24769 25648 24803
rect 25596 24760 25648 24769
rect 26792 24760 26844 24812
rect 27528 24735 27580 24744
rect 27528 24701 27537 24735
rect 27537 24701 27571 24735
rect 27571 24701 27580 24735
rect 27528 24692 27580 24701
rect 27804 24760 27856 24812
rect 31300 24760 31352 24812
rect 31484 24760 31536 24812
rect 31576 24692 31628 24744
rect 33508 24803 33560 24812
rect 33232 24692 33284 24744
rect 33508 24769 33517 24803
rect 33517 24769 33551 24803
rect 33551 24769 33560 24803
rect 33508 24760 33560 24769
rect 34796 24760 34848 24812
rect 36912 24760 36964 24812
rect 34612 24735 34664 24744
rect 34612 24701 34621 24735
rect 34621 24701 34655 24735
rect 34655 24701 34664 24735
rect 34612 24692 34664 24701
rect 35532 24692 35584 24744
rect 37464 24735 37516 24744
rect 37464 24701 37473 24735
rect 37473 24701 37507 24735
rect 37507 24701 37516 24735
rect 37464 24692 37516 24701
rect 38476 24735 38528 24744
rect 38476 24701 38485 24735
rect 38485 24701 38519 24735
rect 38519 24701 38528 24735
rect 38476 24692 38528 24701
rect 44824 24828 44876 24880
rect 40040 24803 40092 24812
rect 40040 24769 40049 24803
rect 40049 24769 40083 24803
rect 40083 24769 40092 24803
rect 40040 24760 40092 24769
rect 46204 24828 46256 24880
rect 46572 24828 46624 24880
rect 46756 24828 46808 24880
rect 47032 24871 47084 24880
rect 47032 24837 47041 24871
rect 47041 24837 47075 24871
rect 47075 24837 47084 24871
rect 47032 24828 47084 24837
rect 47492 24760 47544 24812
rect 46572 24692 46624 24744
rect 11796 24599 11848 24608
rect 11796 24565 11805 24599
rect 11805 24565 11839 24599
rect 11839 24565 11848 24599
rect 11796 24556 11848 24565
rect 13452 24556 13504 24608
rect 14372 24556 14424 24608
rect 19340 24624 19392 24676
rect 15844 24599 15896 24608
rect 15844 24565 15853 24599
rect 15853 24565 15887 24599
rect 15887 24565 15896 24599
rect 15844 24556 15896 24565
rect 16764 24599 16816 24608
rect 16764 24565 16773 24599
rect 16773 24565 16807 24599
rect 16807 24565 16816 24599
rect 16764 24556 16816 24565
rect 18328 24599 18380 24608
rect 18328 24565 18337 24599
rect 18337 24565 18371 24599
rect 18371 24565 18380 24599
rect 23296 24624 23348 24676
rect 27896 24624 27948 24676
rect 46388 24624 46440 24676
rect 18328 24556 18380 24565
rect 28264 24556 28316 24608
rect 30748 24556 30800 24608
rect 33968 24556 34020 24608
rect 35440 24556 35492 24608
rect 37832 24556 37884 24608
rect 40040 24556 40092 24608
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 12072 24352 12124 24404
rect 15936 24352 15988 24404
rect 16028 24352 16080 24404
rect 17316 24352 17368 24404
rect 22468 24352 22520 24404
rect 19340 24284 19392 24336
rect 22192 24284 22244 24336
rect 11796 24259 11848 24268
rect 11796 24225 11805 24259
rect 11805 24225 11839 24259
rect 11839 24225 11848 24259
rect 11796 24216 11848 24225
rect 15844 24216 15896 24268
rect 17868 24216 17920 24268
rect 20536 24216 20588 24268
rect 24308 24284 24360 24336
rect 27896 24284 27948 24336
rect 46020 24352 46072 24404
rect 33232 24327 33284 24336
rect 33232 24293 33241 24327
rect 33241 24293 33275 24327
rect 33275 24293 33284 24327
rect 33232 24284 33284 24293
rect 36912 24327 36964 24336
rect 36912 24293 36921 24327
rect 36921 24293 36955 24327
rect 36955 24293 36964 24327
rect 36912 24284 36964 24293
rect 13360 24148 13412 24200
rect 14372 24191 14424 24200
rect 14372 24157 14381 24191
rect 14381 24157 14415 24191
rect 14415 24157 14424 24191
rect 14372 24148 14424 24157
rect 12072 24123 12124 24132
rect 12072 24089 12081 24123
rect 12081 24089 12115 24123
rect 12115 24089 12124 24123
rect 12072 24080 12124 24089
rect 14004 24080 14056 24132
rect 16764 24148 16816 24200
rect 17408 24148 17460 24200
rect 18328 24148 18380 24200
rect 15200 24080 15252 24132
rect 15384 24080 15436 24132
rect 20076 24148 20128 24200
rect 20996 24191 21048 24200
rect 20996 24157 21005 24191
rect 21005 24157 21039 24191
rect 21039 24157 21048 24191
rect 20996 24148 21048 24157
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 24768 24148 24820 24200
rect 30748 24259 30800 24268
rect 30748 24225 30757 24259
rect 30757 24225 30791 24259
rect 30791 24225 30800 24259
rect 30748 24216 30800 24225
rect 35440 24259 35492 24268
rect 35440 24225 35449 24259
rect 35449 24225 35483 24259
rect 35483 24225 35492 24259
rect 35440 24216 35492 24225
rect 35808 24216 35860 24268
rect 40316 24259 40368 24268
rect 40316 24225 40325 24259
rect 40325 24225 40359 24259
rect 40359 24225 40368 24259
rect 40316 24216 40368 24225
rect 47768 24284 47820 24336
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 26516 24148 26568 24200
rect 29552 24191 29604 24200
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 30472 24191 30524 24200
rect 30472 24157 30481 24191
rect 30481 24157 30515 24191
rect 30515 24157 30524 24191
rect 30472 24148 30524 24157
rect 32956 24148 33008 24200
rect 34520 24148 34572 24200
rect 34796 24148 34848 24200
rect 39856 24191 39908 24200
rect 39856 24157 39865 24191
rect 39865 24157 39899 24191
rect 39899 24157 39908 24191
rect 39856 24148 39908 24157
rect 20352 24080 20404 24132
rect 31760 24080 31812 24132
rect 32680 24123 32732 24132
rect 32680 24089 32689 24123
rect 32689 24089 32723 24123
rect 32723 24089 32732 24123
rect 32680 24080 32732 24089
rect 32772 24080 32824 24132
rect 12348 24012 12400 24064
rect 14096 24012 14148 24064
rect 15660 24012 15712 24064
rect 17132 24012 17184 24064
rect 18328 24012 18380 24064
rect 20812 24012 20864 24064
rect 21824 24012 21876 24064
rect 25412 24055 25464 24064
rect 25412 24021 25421 24055
rect 25421 24021 25455 24055
rect 25455 24021 25464 24055
rect 25412 24012 25464 24021
rect 29644 24055 29696 24064
rect 29644 24021 29653 24055
rect 29653 24021 29687 24055
rect 29687 24021 29696 24055
rect 29644 24012 29696 24021
rect 32128 24012 32180 24064
rect 34060 24055 34112 24064
rect 34060 24021 34069 24055
rect 34069 24021 34103 24055
rect 34103 24021 34112 24055
rect 34060 24012 34112 24021
rect 35992 24080 36044 24132
rect 37648 24123 37700 24132
rect 37648 24089 37657 24123
rect 37657 24089 37691 24123
rect 37691 24089 37700 24123
rect 37648 24080 37700 24089
rect 39304 24123 39356 24132
rect 39304 24089 39313 24123
rect 39313 24089 39347 24123
rect 39347 24089 39356 24123
rect 39304 24080 39356 24089
rect 40040 24123 40092 24132
rect 40040 24089 40049 24123
rect 40049 24089 40083 24123
rect 40083 24089 40092 24123
rect 40040 24080 40092 24089
rect 36084 24012 36136 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 11704 23808 11756 23860
rect 13452 23851 13504 23860
rect 12992 23740 13044 23792
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 11980 23715 12032 23724
rect 11980 23681 11989 23715
rect 11989 23681 12023 23715
rect 12023 23681 12032 23715
rect 11980 23672 12032 23681
rect 12348 23715 12400 23724
rect 11612 23604 11664 23656
rect 12348 23681 12357 23715
rect 12357 23681 12391 23715
rect 12391 23681 12400 23715
rect 13452 23817 13461 23851
rect 13461 23817 13495 23851
rect 13495 23817 13504 23851
rect 13452 23808 13504 23817
rect 14004 23851 14056 23860
rect 14004 23817 14013 23851
rect 14013 23817 14047 23851
rect 14047 23817 14056 23851
rect 14004 23808 14056 23817
rect 14096 23808 14148 23860
rect 15200 23808 15252 23860
rect 20812 23851 20864 23860
rect 20812 23817 20821 23851
rect 20821 23817 20855 23851
rect 20855 23817 20864 23851
rect 20812 23808 20864 23817
rect 21364 23808 21416 23860
rect 15016 23740 15068 23792
rect 20536 23740 20588 23792
rect 26792 23808 26844 23860
rect 30472 23851 30524 23860
rect 28264 23783 28316 23792
rect 28264 23749 28273 23783
rect 28273 23749 28307 23783
rect 28307 23749 28316 23783
rect 28264 23740 28316 23749
rect 29644 23740 29696 23792
rect 30472 23817 30481 23851
rect 30481 23817 30515 23851
rect 30515 23817 30524 23851
rect 30472 23808 30524 23817
rect 33508 23808 33560 23860
rect 12348 23672 12400 23681
rect 13360 23672 13412 23724
rect 13912 23715 13964 23724
rect 13912 23681 13921 23715
rect 13921 23681 13955 23715
rect 13955 23681 13964 23715
rect 13912 23672 13964 23681
rect 14280 23672 14332 23724
rect 13728 23604 13780 23656
rect 16948 23672 17000 23724
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 17132 23672 17184 23681
rect 19616 23672 19668 23724
rect 19892 23715 19944 23724
rect 19892 23681 19901 23715
rect 19901 23681 19935 23715
rect 19935 23681 19944 23715
rect 19892 23672 19944 23681
rect 19984 23715 20036 23724
rect 19984 23681 19993 23715
rect 19993 23681 20027 23715
rect 20027 23681 20036 23715
rect 20628 23715 20680 23724
rect 19984 23672 20036 23681
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 20720 23715 20772 23724
rect 20720 23681 20729 23715
rect 20729 23681 20763 23715
rect 20763 23681 20772 23715
rect 21824 23715 21876 23724
rect 20720 23672 20772 23681
rect 21824 23681 21833 23715
rect 21833 23681 21867 23715
rect 21867 23681 21876 23715
rect 21824 23672 21876 23681
rect 23204 23672 23256 23724
rect 25872 23672 25924 23724
rect 27896 23672 27948 23724
rect 32128 23783 32180 23792
rect 32128 23749 32137 23783
rect 32137 23749 32171 23783
rect 32171 23749 32180 23783
rect 32128 23740 32180 23749
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 16028 23604 16080 23656
rect 21456 23604 21508 23656
rect 22100 23647 22152 23656
rect 22100 23613 22109 23647
rect 22109 23613 22143 23647
rect 22143 23613 22152 23647
rect 22100 23604 22152 23613
rect 14280 23536 14332 23588
rect 16396 23536 16448 23588
rect 12348 23511 12400 23520
rect 12348 23477 12357 23511
rect 12357 23477 12391 23511
rect 12391 23477 12400 23511
rect 12348 23468 12400 23477
rect 12992 23468 13044 23520
rect 18052 23536 18104 23588
rect 27896 23536 27948 23588
rect 30840 23604 30892 23656
rect 31300 23579 31352 23588
rect 31300 23545 31309 23579
rect 31309 23545 31343 23579
rect 31343 23545 31352 23579
rect 31300 23536 31352 23545
rect 17132 23468 17184 23520
rect 19524 23511 19576 23520
rect 19524 23477 19533 23511
rect 19533 23477 19567 23511
rect 19567 23477 19576 23511
rect 19524 23468 19576 23477
rect 25228 23468 25280 23520
rect 31576 23715 31628 23724
rect 31576 23681 31585 23715
rect 31585 23681 31619 23715
rect 31619 23681 31628 23715
rect 32680 23740 32732 23792
rect 35532 23808 35584 23860
rect 35992 23851 36044 23860
rect 35992 23817 36001 23851
rect 36001 23817 36035 23851
rect 36035 23817 36044 23851
rect 35992 23808 36044 23817
rect 37648 23808 37700 23860
rect 40040 23808 40092 23860
rect 46572 23808 46624 23860
rect 33968 23783 34020 23792
rect 33968 23749 33977 23783
rect 33977 23749 34011 23783
rect 34011 23749 34020 23783
rect 33968 23740 34020 23749
rect 34060 23740 34112 23792
rect 31576 23672 31628 23681
rect 33048 23672 33100 23724
rect 37464 23715 37516 23724
rect 31484 23536 31536 23588
rect 33692 23647 33744 23656
rect 33692 23613 33701 23647
rect 33701 23613 33735 23647
rect 33735 23613 33744 23647
rect 33692 23604 33744 23613
rect 34520 23604 34572 23656
rect 37464 23681 37473 23715
rect 37473 23681 37507 23715
rect 37507 23681 37516 23715
rect 37464 23672 37516 23681
rect 39212 23715 39264 23724
rect 39212 23681 39221 23715
rect 39221 23681 39255 23715
rect 39255 23681 39264 23715
rect 44916 23740 44968 23792
rect 39212 23672 39264 23681
rect 42984 23715 43036 23724
rect 42984 23681 42993 23715
rect 42993 23681 43027 23715
rect 43027 23681 43036 23715
rect 42984 23672 43036 23681
rect 47032 23715 47084 23724
rect 43444 23604 43496 23656
rect 47032 23681 47041 23715
rect 47041 23681 47075 23715
rect 47075 23681 47084 23715
rect 47032 23672 47084 23681
rect 47584 23715 47636 23724
rect 47584 23681 47593 23715
rect 47593 23681 47627 23715
rect 47627 23681 47636 23715
rect 47584 23672 47636 23681
rect 48044 23604 48096 23656
rect 32772 23468 32824 23520
rect 33784 23468 33836 23520
rect 37832 23468 37884 23520
rect 42800 23511 42852 23520
rect 42800 23477 42809 23511
rect 42809 23477 42843 23511
rect 42843 23477 42852 23511
rect 42800 23468 42852 23477
rect 45744 23511 45796 23520
rect 45744 23477 45753 23511
rect 45753 23477 45787 23511
rect 45787 23477 45796 23511
rect 45744 23468 45796 23477
rect 46572 23468 46624 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 12072 23264 12124 23316
rect 16580 23264 16632 23316
rect 16948 23264 17000 23316
rect 17868 23307 17920 23316
rect 17868 23273 17877 23307
rect 17877 23273 17911 23307
rect 17911 23273 17920 23307
rect 17868 23264 17920 23273
rect 22100 23264 22152 23316
rect 23204 23307 23256 23316
rect 23204 23273 23213 23307
rect 23213 23273 23247 23307
rect 23247 23273 23256 23307
rect 23204 23264 23256 23273
rect 12348 23103 12400 23112
rect 12348 23069 12357 23103
rect 12357 23069 12391 23103
rect 12391 23069 12400 23103
rect 12348 23060 12400 23069
rect 13452 23060 13504 23112
rect 16028 23128 16080 23180
rect 16396 23171 16448 23180
rect 16396 23137 16405 23171
rect 16405 23137 16439 23171
rect 16439 23137 16448 23171
rect 16396 23128 16448 23137
rect 19524 23128 19576 23180
rect 29552 23264 29604 23316
rect 27804 23128 27856 23180
rect 27988 23171 28040 23180
rect 27988 23137 27997 23171
rect 27997 23137 28031 23171
rect 28031 23137 28040 23171
rect 27988 23128 28040 23137
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 19340 23060 19392 23112
rect 19892 23060 19944 23112
rect 20812 23060 20864 23112
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 21456 23103 21508 23112
rect 20996 23060 21048 23069
rect 21456 23069 21465 23103
rect 21465 23069 21499 23103
rect 21499 23069 21508 23103
rect 21456 23060 21508 23069
rect 22192 23103 22244 23112
rect 22192 23069 22201 23103
rect 22201 23069 22235 23103
rect 22235 23069 22244 23103
rect 22192 23060 22244 23069
rect 22376 23103 22428 23112
rect 22376 23069 22385 23103
rect 22385 23069 22419 23103
rect 22419 23069 22428 23103
rect 22376 23060 22428 23069
rect 23940 23060 23992 23112
rect 26792 23103 26844 23112
rect 26792 23069 26801 23103
rect 26801 23069 26835 23103
rect 26835 23069 26844 23103
rect 26792 23060 26844 23069
rect 17132 22992 17184 23044
rect 19616 22992 19668 23044
rect 20168 22992 20220 23044
rect 24768 23035 24820 23044
rect 24768 23001 24777 23035
rect 24777 23001 24811 23035
rect 24811 23001 24820 23035
rect 24768 22992 24820 23001
rect 25412 22992 25464 23044
rect 26976 23035 27028 23044
rect 18328 22924 18380 22976
rect 19432 22924 19484 22976
rect 20536 22924 20588 22976
rect 20812 22967 20864 22976
rect 20812 22933 20821 22967
rect 20821 22933 20855 22967
rect 20855 22933 20864 22967
rect 20812 22924 20864 22933
rect 21824 22924 21876 22976
rect 23296 22924 23348 22976
rect 26148 22924 26200 22976
rect 26976 23001 26985 23035
rect 26985 23001 27019 23035
rect 27019 23001 27028 23035
rect 26976 22992 27028 23001
rect 29644 23060 29696 23112
rect 31760 23264 31812 23316
rect 33692 23307 33744 23316
rect 33692 23273 33701 23307
rect 33701 23273 33735 23307
rect 33735 23273 33744 23307
rect 33692 23264 33744 23273
rect 34796 23307 34848 23316
rect 34796 23273 34805 23307
rect 34805 23273 34839 23307
rect 34839 23273 34848 23307
rect 34796 23264 34848 23273
rect 38108 23264 38160 23316
rect 38660 23264 38712 23316
rect 42984 23264 43036 23316
rect 29920 23196 29972 23248
rect 30840 23103 30892 23112
rect 30840 23069 30849 23103
rect 30849 23069 30883 23103
rect 30883 23069 30892 23103
rect 30840 23060 30892 23069
rect 38384 23128 38436 23180
rect 39856 23128 39908 23180
rect 42340 23128 42392 23180
rect 38936 23103 38988 23112
rect 32128 22992 32180 23044
rect 33876 22992 33928 23044
rect 38936 23069 38945 23103
rect 38945 23069 38979 23103
rect 38979 23069 38988 23103
rect 38936 23060 38988 23069
rect 45744 23128 45796 23180
rect 46388 23171 46440 23180
rect 46388 23137 46397 23171
rect 46397 23137 46431 23171
rect 46431 23137 46440 23171
rect 46388 23128 46440 23137
rect 40132 23035 40184 23044
rect 30932 22924 30984 22976
rect 37280 22924 37332 22976
rect 39580 22924 39632 22976
rect 40132 23001 40141 23035
rect 40141 23001 40175 23035
rect 40175 23001 40184 23035
rect 40132 22992 40184 23001
rect 41788 23035 41840 23044
rect 41788 23001 41797 23035
rect 41797 23001 41831 23035
rect 41831 23001 41840 23035
rect 41788 22992 41840 23001
rect 41880 22992 41932 23044
rect 45008 23060 45060 23112
rect 47308 23060 47360 23112
rect 47952 23035 48004 23044
rect 47952 23001 47961 23035
rect 47961 23001 47995 23035
rect 47995 23001 48004 23035
rect 47952 22992 48004 23001
rect 43260 22924 43312 22976
rect 43444 22967 43496 22976
rect 43444 22933 43453 22967
rect 43453 22933 43487 22967
rect 43487 22933 43496 22967
rect 43444 22924 43496 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 16028 22763 16080 22772
rect 16028 22729 16037 22763
rect 16037 22729 16071 22763
rect 16071 22729 16080 22763
rect 16028 22720 16080 22729
rect 16212 22720 16264 22772
rect 16856 22720 16908 22772
rect 17868 22720 17920 22772
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 14648 22584 14700 22636
rect 15476 22652 15528 22704
rect 17684 22652 17736 22704
rect 18328 22652 18380 22704
rect 19340 22720 19392 22772
rect 19432 22720 19484 22772
rect 20076 22720 20128 22772
rect 24768 22763 24820 22772
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 16672 22627 16724 22636
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 11980 22516 12032 22568
rect 12532 22516 12584 22568
rect 15200 22516 15252 22568
rect 17316 22559 17368 22568
rect 17316 22525 17325 22559
rect 17325 22525 17359 22559
rect 17359 22525 17368 22559
rect 17316 22516 17368 22525
rect 18604 22516 18656 22568
rect 20536 22652 20588 22704
rect 20812 22652 20864 22704
rect 24768 22729 24777 22763
rect 24777 22729 24811 22763
rect 24811 22729 24820 22763
rect 24768 22720 24820 22729
rect 26976 22720 27028 22772
rect 27344 22720 27396 22772
rect 27804 22720 27856 22772
rect 32864 22720 32916 22772
rect 39856 22720 39908 22772
rect 41788 22720 41840 22772
rect 46388 22720 46440 22772
rect 48044 22763 48096 22772
rect 48044 22729 48053 22763
rect 48053 22729 48087 22763
rect 48087 22729 48096 22763
rect 48044 22720 48096 22729
rect 20628 22627 20680 22636
rect 11796 22380 11848 22432
rect 12348 22380 12400 22432
rect 13728 22380 13780 22432
rect 15200 22423 15252 22432
rect 15200 22389 15209 22423
rect 15209 22389 15243 22423
rect 15243 22389 15252 22423
rect 15200 22380 15252 22389
rect 20628 22593 20637 22627
rect 20637 22593 20671 22627
rect 20671 22593 20680 22627
rect 20628 22584 20680 22593
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 21824 22627 21876 22636
rect 20720 22584 20772 22593
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 23940 22584 23992 22636
rect 20168 22516 20220 22568
rect 26516 22652 26568 22704
rect 38108 22695 38160 22704
rect 38108 22661 38117 22695
rect 38117 22661 38151 22695
rect 38151 22661 38160 22695
rect 38108 22652 38160 22661
rect 24676 22627 24728 22636
rect 24676 22593 24685 22627
rect 24685 22593 24719 22627
rect 24719 22593 24728 22627
rect 24676 22584 24728 22593
rect 19340 22380 19392 22432
rect 19984 22380 20036 22432
rect 25596 22448 25648 22500
rect 26148 22584 26200 22636
rect 31852 22584 31904 22636
rect 32128 22627 32180 22636
rect 32128 22593 32137 22627
rect 32137 22593 32171 22627
rect 32171 22593 32180 22627
rect 32128 22584 32180 22593
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 35348 22584 35400 22636
rect 37280 22627 37332 22636
rect 37280 22593 37289 22627
rect 37289 22593 37323 22627
rect 37323 22593 37332 22627
rect 37280 22584 37332 22593
rect 31484 22516 31536 22568
rect 39580 22559 39632 22568
rect 39580 22525 39589 22559
rect 39589 22525 39623 22559
rect 39623 22525 39632 22559
rect 39580 22516 39632 22525
rect 40040 22584 40092 22636
rect 41880 22627 41932 22636
rect 40224 22516 40276 22568
rect 41880 22593 41889 22627
rect 41889 22593 41923 22627
rect 41923 22593 41932 22627
rect 41880 22584 41932 22593
rect 42800 22584 42852 22636
rect 45836 22652 45888 22704
rect 42340 22516 42392 22568
rect 42892 22559 42944 22568
rect 42892 22525 42901 22559
rect 42901 22525 42935 22559
rect 42935 22525 42944 22559
rect 42892 22516 42944 22525
rect 45192 22559 45244 22568
rect 45192 22525 45201 22559
rect 45201 22525 45235 22559
rect 45235 22525 45244 22559
rect 45192 22516 45244 22525
rect 46388 22559 46440 22568
rect 33876 22448 33928 22500
rect 35900 22448 35952 22500
rect 46388 22525 46397 22559
rect 46397 22525 46431 22559
rect 46431 22525 46440 22559
rect 46388 22516 46440 22525
rect 45928 22448 45980 22500
rect 20352 22380 20404 22432
rect 22192 22380 22244 22432
rect 27896 22380 27948 22432
rect 31208 22380 31260 22432
rect 32220 22423 32272 22432
rect 32220 22389 32229 22423
rect 32229 22389 32263 22423
rect 32263 22389 32272 22423
rect 32220 22380 32272 22389
rect 32956 22380 33008 22432
rect 33692 22380 33744 22432
rect 34796 22380 34848 22432
rect 40592 22423 40644 22432
rect 40592 22389 40601 22423
rect 40601 22389 40635 22423
rect 40635 22389 40644 22423
rect 40592 22380 40644 22389
rect 40868 22380 40920 22432
rect 41788 22423 41840 22432
rect 41788 22389 41797 22423
rect 41797 22389 41831 22423
rect 41831 22389 41840 22423
rect 41788 22380 41840 22389
rect 45100 22380 45152 22432
rect 45652 22380 45704 22432
rect 47216 22380 47268 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 11796 22219 11848 22228
rect 11796 22185 11826 22219
rect 11826 22185 11848 22219
rect 11796 22176 11848 22185
rect 17316 22176 17368 22228
rect 14648 22108 14700 22160
rect 15844 22108 15896 22160
rect 26148 22176 26200 22228
rect 31208 22219 31260 22228
rect 31208 22185 31238 22219
rect 31238 22185 31260 22219
rect 31208 22176 31260 22185
rect 18604 22108 18656 22160
rect 11796 22040 11848 22092
rect 15200 22040 15252 22092
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 19340 22083 19392 22092
rect 15292 22040 15344 22049
rect 19340 22049 19349 22083
rect 19349 22049 19383 22083
rect 19383 22049 19392 22083
rect 19340 22040 19392 22049
rect 22192 22040 22244 22092
rect 25964 22108 26016 22160
rect 35348 22176 35400 22228
rect 35624 22176 35676 22228
rect 40132 22176 40184 22228
rect 45192 22176 45244 22228
rect 45468 22176 45520 22228
rect 45652 22219 45704 22228
rect 45652 22185 45661 22219
rect 45661 22185 45695 22219
rect 45695 22185 45704 22219
rect 45652 22176 45704 22185
rect 45836 22219 45888 22228
rect 45836 22185 45845 22219
rect 45845 22185 45879 22219
rect 45879 22185 45888 22219
rect 45836 22176 45888 22185
rect 28908 22040 28960 22092
rect 30932 22083 30984 22092
rect 11520 22015 11572 22024
rect 11520 21981 11529 22015
rect 11529 21981 11563 22015
rect 11563 21981 11572 22015
rect 11520 21972 11572 21981
rect 13084 21904 13136 21956
rect 16212 21972 16264 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 24860 21972 24912 22024
rect 25228 22015 25280 22024
rect 25228 21981 25237 22015
rect 25237 21981 25271 22015
rect 25271 21981 25280 22015
rect 25228 21972 25280 21981
rect 25688 21972 25740 22024
rect 27436 22015 27488 22024
rect 27436 21981 27445 22015
rect 27445 21981 27479 22015
rect 27479 21981 27488 22015
rect 27436 21972 27488 21981
rect 27896 21972 27948 22024
rect 29000 22015 29052 22024
rect 29000 21981 29009 22015
rect 29009 21981 29043 22015
rect 29043 21981 29052 22015
rect 29000 21972 29052 21981
rect 30932 22049 30941 22083
rect 30941 22049 30975 22083
rect 30975 22049 30984 22083
rect 30932 22040 30984 22049
rect 31760 22040 31812 22092
rect 33048 22040 33100 22092
rect 40224 22040 40276 22092
rect 45928 22108 45980 22160
rect 32496 21972 32548 22024
rect 32956 22015 33008 22024
rect 32956 21981 32965 22015
rect 32965 21981 32999 22015
rect 32999 21981 33008 22015
rect 32956 21972 33008 21981
rect 34704 22015 34756 22024
rect 34704 21981 34713 22015
rect 34713 21981 34747 22015
rect 34747 21981 34756 22015
rect 34704 21972 34756 21981
rect 16580 21904 16632 21956
rect 24676 21904 24728 21956
rect 32220 21904 32272 21956
rect 33784 21947 33836 21956
rect 24400 21879 24452 21888
rect 24400 21845 24409 21879
rect 24409 21845 24443 21879
rect 24443 21845 24452 21879
rect 24400 21836 24452 21845
rect 25320 21879 25372 21888
rect 25320 21845 25329 21879
rect 25329 21845 25363 21879
rect 25363 21845 25372 21879
rect 25320 21836 25372 21845
rect 27712 21836 27764 21888
rect 28448 21836 28500 21888
rect 28816 21879 28868 21888
rect 28816 21845 28825 21879
rect 28825 21845 28859 21879
rect 28859 21845 28868 21879
rect 28816 21836 28868 21845
rect 29736 21836 29788 21888
rect 30196 21836 30248 21888
rect 33784 21913 33793 21947
rect 33793 21913 33827 21947
rect 33827 21913 33836 21947
rect 33784 21904 33836 21913
rect 40040 21972 40092 22024
rect 40592 21972 40644 22024
rect 40868 22015 40920 22024
rect 40868 21981 40877 22015
rect 40877 21981 40911 22015
rect 40911 21981 40920 22015
rect 40868 21972 40920 21981
rect 41788 21972 41840 22024
rect 42800 21972 42852 22024
rect 45468 22040 45520 22092
rect 46480 22083 46532 22092
rect 46480 22049 46489 22083
rect 46489 22049 46523 22083
rect 46523 22049 46532 22083
rect 46480 22040 46532 22049
rect 46756 22083 46808 22092
rect 46756 22049 46765 22083
rect 46765 22049 46799 22083
rect 46799 22049 46808 22083
rect 46756 22040 46808 22049
rect 44456 22015 44508 22024
rect 44456 21981 44465 22015
rect 44465 21981 44499 22015
rect 44499 21981 44508 22015
rect 44456 21972 44508 21981
rect 45560 22015 45612 22024
rect 36360 21879 36412 21888
rect 36360 21845 36369 21879
rect 36369 21845 36403 21879
rect 36403 21845 36412 21879
rect 36360 21836 36412 21845
rect 36636 21904 36688 21956
rect 40224 21947 40276 21956
rect 37188 21836 37240 21888
rect 40224 21913 40233 21947
rect 40233 21913 40267 21947
rect 40267 21913 40276 21947
rect 40224 21904 40276 21913
rect 43444 21904 43496 21956
rect 45100 21904 45152 21956
rect 45560 21981 45569 22015
rect 45569 21981 45603 22015
rect 45603 21981 45612 22015
rect 45560 21972 45612 21981
rect 46020 21904 46072 21956
rect 45652 21836 45704 21888
rect 46296 21836 46348 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11520 21632 11572 21684
rect 13084 21675 13136 21684
rect 13084 21641 13093 21675
rect 13093 21641 13127 21675
rect 13127 21641 13136 21675
rect 13084 21632 13136 21641
rect 22192 21632 22244 21684
rect 3608 21564 3660 21616
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 12348 21496 12400 21548
rect 13820 21496 13872 21548
rect 20 21360 72 21412
rect 11428 21360 11480 21412
rect 15384 21564 15436 21616
rect 18512 21496 18564 21548
rect 18880 21539 18932 21548
rect 18880 21505 18889 21539
rect 18889 21505 18923 21539
rect 18923 21505 18932 21539
rect 18880 21496 18932 21505
rect 22284 21539 22336 21548
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 24676 21632 24728 21684
rect 25136 21632 25188 21684
rect 25596 21632 25648 21684
rect 36636 21675 36688 21684
rect 24400 21564 24452 21616
rect 25320 21564 25372 21616
rect 14464 21428 14516 21480
rect 24308 21428 24360 21480
rect 28816 21564 28868 21616
rect 29736 21564 29788 21616
rect 26884 21496 26936 21548
rect 27252 21496 27304 21548
rect 28448 21539 28500 21548
rect 28448 21505 28457 21539
rect 28457 21505 28491 21539
rect 28491 21505 28500 21539
rect 28448 21496 28500 21505
rect 32496 21539 32548 21548
rect 32496 21505 32505 21539
rect 32505 21505 32539 21539
rect 32539 21505 32548 21539
rect 32496 21496 32548 21505
rect 35348 21539 35400 21548
rect 35348 21505 35357 21539
rect 35357 21505 35391 21539
rect 35391 21505 35400 21539
rect 35348 21496 35400 21505
rect 27160 21428 27212 21480
rect 30196 21471 30248 21480
rect 30196 21437 30205 21471
rect 30205 21437 30239 21471
rect 30239 21437 30248 21471
rect 30196 21428 30248 21437
rect 32772 21471 32824 21480
rect 32772 21437 32781 21471
rect 32781 21437 32815 21471
rect 32815 21437 32824 21471
rect 32772 21428 32824 21437
rect 20904 21360 20956 21412
rect 15752 21292 15804 21344
rect 16672 21292 16724 21344
rect 17960 21335 18012 21344
rect 17960 21301 17969 21335
rect 17969 21301 18003 21335
rect 18003 21301 18012 21335
rect 17960 21292 18012 21301
rect 18972 21335 19024 21344
rect 18972 21301 18981 21335
rect 18981 21301 19015 21335
rect 19015 21301 19024 21335
rect 18972 21292 19024 21301
rect 30288 21360 30340 21412
rect 36636 21641 36645 21675
rect 36645 21641 36679 21675
rect 36679 21641 36688 21675
rect 36636 21632 36688 21641
rect 40040 21632 40092 21684
rect 46020 21632 46072 21684
rect 37280 21564 37332 21616
rect 38936 21564 38988 21616
rect 43536 21564 43588 21616
rect 45468 21607 45520 21616
rect 45468 21573 45477 21607
rect 45477 21573 45511 21607
rect 45511 21573 45520 21607
rect 45468 21564 45520 21573
rect 42708 21539 42760 21548
rect 42708 21505 42717 21539
rect 42717 21505 42751 21539
rect 42751 21505 42760 21539
rect 42708 21496 42760 21505
rect 43812 21539 43864 21548
rect 25688 21292 25740 21344
rect 25964 21292 26016 21344
rect 27896 21292 27948 21344
rect 32772 21292 32824 21344
rect 38200 21360 38252 21412
rect 42616 21428 42668 21480
rect 43812 21505 43821 21539
rect 43821 21505 43855 21539
rect 43855 21505 43864 21539
rect 43812 21496 43864 21505
rect 43996 21539 44048 21548
rect 43996 21505 44005 21539
rect 44005 21505 44039 21539
rect 44039 21505 44048 21539
rect 43996 21496 44048 21505
rect 45836 21496 45888 21548
rect 46572 21564 46624 21616
rect 46204 21539 46256 21548
rect 46204 21505 46213 21539
rect 46213 21505 46247 21539
rect 46247 21505 46256 21539
rect 46204 21496 46256 21505
rect 46296 21496 46348 21548
rect 46112 21428 46164 21480
rect 44364 21360 44416 21412
rect 44456 21360 44508 21412
rect 38936 21335 38988 21344
rect 38936 21301 38945 21335
rect 38945 21301 38979 21335
rect 38979 21301 38988 21335
rect 38936 21292 38988 21301
rect 43168 21292 43220 21344
rect 44272 21292 44324 21344
rect 44732 21335 44784 21344
rect 44732 21301 44741 21335
rect 44741 21301 44775 21335
rect 44775 21301 44784 21335
rect 44732 21292 44784 21301
rect 45284 21360 45336 21412
rect 47216 21292 47268 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2228 21088 2280 21140
rect 25688 21020 25740 21072
rect 33416 21020 33468 21072
rect 3700 20952 3752 21004
rect 11428 20952 11480 21004
rect 22836 20995 22888 21004
rect 22836 20961 22845 20995
rect 22845 20961 22879 20995
rect 22879 20961 22888 20995
rect 22836 20952 22888 20961
rect 24308 20952 24360 21004
rect 24860 20995 24912 21004
rect 24860 20961 24869 20995
rect 24869 20961 24903 20995
rect 24903 20961 24912 20995
rect 24860 20952 24912 20961
rect 25596 20995 25648 21004
rect 25596 20961 25605 20995
rect 25605 20961 25639 20995
rect 25639 20961 25648 20995
rect 25596 20952 25648 20961
rect 25964 20952 26016 21004
rect 27712 20995 27764 21004
rect 27712 20961 27721 20995
rect 27721 20961 27755 20995
rect 27755 20961 27764 20995
rect 27712 20952 27764 20961
rect 13820 20884 13872 20936
rect 14372 20884 14424 20936
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 14648 20884 14700 20893
rect 15752 20927 15804 20936
rect 15752 20893 15761 20927
rect 15761 20893 15795 20927
rect 15795 20893 15804 20927
rect 15752 20884 15804 20893
rect 16396 20927 16448 20936
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 17960 20884 18012 20936
rect 20352 20884 20404 20936
rect 22560 20884 22612 20936
rect 25504 20884 25556 20936
rect 11060 20859 11112 20868
rect 11060 20825 11069 20859
rect 11069 20825 11103 20859
rect 11103 20825 11112 20859
rect 11060 20816 11112 20825
rect 21272 20859 21324 20868
rect 21272 20825 21281 20859
rect 21281 20825 21315 20859
rect 21315 20825 21324 20859
rect 21272 20816 21324 20825
rect 25320 20816 25372 20868
rect 26056 20884 26108 20936
rect 26976 20927 27028 20936
rect 26976 20893 26985 20927
rect 26985 20893 27019 20927
rect 27019 20893 27028 20927
rect 26976 20884 27028 20893
rect 27436 20884 27488 20936
rect 30288 20952 30340 21004
rect 31760 20952 31812 21004
rect 11888 20748 11940 20800
rect 13268 20791 13320 20800
rect 13268 20757 13277 20791
rect 13277 20757 13311 20791
rect 13311 20757 13320 20791
rect 13268 20748 13320 20757
rect 16672 20748 16724 20800
rect 17500 20748 17552 20800
rect 20352 20748 20404 20800
rect 25780 20748 25832 20800
rect 26148 20816 26200 20868
rect 27896 20884 27948 20936
rect 28908 20884 28960 20936
rect 33692 20927 33744 20936
rect 33692 20893 33701 20927
rect 33701 20893 33735 20927
rect 33735 20893 33744 20927
rect 33692 20884 33744 20893
rect 42800 21088 42852 21140
rect 44364 21088 44416 21140
rect 47584 21088 47636 21140
rect 35440 21020 35492 21072
rect 47492 21020 47544 21072
rect 38936 20952 38988 21004
rect 37280 20927 37332 20936
rect 37280 20893 37289 20927
rect 37289 20893 37323 20927
rect 37323 20893 37332 20927
rect 37280 20884 37332 20893
rect 38016 20927 38068 20936
rect 38016 20893 38025 20927
rect 38025 20893 38059 20927
rect 38059 20893 38068 20927
rect 38016 20884 38068 20893
rect 42248 20927 42300 20936
rect 28724 20816 28776 20868
rect 31392 20859 31444 20868
rect 27896 20748 27948 20800
rect 28172 20791 28224 20800
rect 28172 20757 28181 20791
rect 28181 20757 28215 20791
rect 28215 20757 28224 20791
rect 28172 20748 28224 20757
rect 28540 20748 28592 20800
rect 29828 20748 29880 20800
rect 31392 20825 31401 20859
rect 31401 20825 31435 20859
rect 31435 20825 31444 20859
rect 31392 20816 31444 20825
rect 33048 20859 33100 20868
rect 33048 20825 33057 20859
rect 33057 20825 33091 20859
rect 33091 20825 33100 20859
rect 33048 20816 33100 20825
rect 35072 20859 35124 20868
rect 35072 20825 35081 20859
rect 35081 20825 35115 20859
rect 35115 20825 35124 20859
rect 35992 20859 36044 20868
rect 35072 20816 35124 20825
rect 35992 20825 36001 20859
rect 36001 20825 36035 20859
rect 36035 20825 36044 20859
rect 35992 20816 36044 20825
rect 42248 20893 42257 20927
rect 42257 20893 42291 20927
rect 42291 20893 42300 20927
rect 42248 20884 42300 20893
rect 42892 20927 42944 20936
rect 42892 20893 42901 20927
rect 42901 20893 42935 20927
rect 42935 20893 42944 20927
rect 42892 20884 42944 20893
rect 44732 20952 44784 21004
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 43168 20927 43220 20936
rect 43168 20893 43177 20927
rect 43177 20893 43211 20927
rect 43211 20893 43220 20927
rect 43720 20927 43772 20936
rect 43168 20884 43220 20893
rect 43720 20893 43729 20927
rect 43729 20893 43763 20927
rect 43763 20893 43772 20927
rect 43720 20884 43772 20893
rect 43904 20927 43956 20936
rect 43904 20893 43913 20927
rect 43913 20893 43947 20927
rect 43947 20893 43956 20927
rect 43904 20884 43956 20893
rect 45284 20884 45336 20936
rect 43536 20816 43588 20868
rect 42800 20748 42852 20800
rect 42892 20748 42944 20800
rect 43168 20748 43220 20800
rect 43812 20791 43864 20800
rect 43812 20757 43821 20791
rect 43821 20757 43855 20791
rect 43855 20757 43864 20791
rect 43812 20748 43864 20757
rect 45376 20748 45428 20800
rect 45560 20748 45612 20800
rect 46020 20748 46072 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 11060 20544 11112 20596
rect 3976 20476 4028 20528
rect 13268 20476 13320 20528
rect 15384 20519 15436 20528
rect 15384 20485 15393 20519
rect 15393 20485 15427 20519
rect 15427 20485 15436 20519
rect 15384 20476 15436 20485
rect 18972 20519 19024 20528
rect 18972 20485 18981 20519
rect 18981 20485 19015 20519
rect 19015 20485 19024 20519
rect 18972 20476 19024 20485
rect 19156 20544 19208 20596
rect 22652 20544 22704 20596
rect 25596 20544 25648 20596
rect 26056 20544 26108 20596
rect 26976 20587 27028 20596
rect 26976 20553 26985 20587
rect 26985 20553 27019 20587
rect 27019 20553 27028 20587
rect 26976 20544 27028 20553
rect 29000 20544 29052 20596
rect 30288 20587 30340 20596
rect 30288 20553 30297 20587
rect 30297 20553 30331 20587
rect 30331 20553 30340 20587
rect 30288 20544 30340 20553
rect 31392 20587 31444 20596
rect 31392 20553 31401 20587
rect 31401 20553 31435 20587
rect 31435 20553 31444 20587
rect 31392 20544 31444 20553
rect 42248 20544 42300 20596
rect 42984 20544 43036 20596
rect 46480 20544 46532 20596
rect 25780 20519 25832 20528
rect 11428 20408 11480 20460
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 15752 20408 15804 20460
rect 16212 20408 16264 20460
rect 17408 20408 17460 20460
rect 17500 20451 17552 20460
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 22192 20408 22244 20460
rect 23296 20408 23348 20460
rect 24676 20408 24728 20460
rect 25780 20485 25789 20519
rect 25789 20485 25823 20519
rect 25823 20485 25832 20519
rect 25780 20476 25832 20485
rect 25872 20519 25924 20528
rect 25872 20485 25881 20519
rect 25881 20485 25915 20519
rect 25915 20485 25924 20519
rect 25872 20476 25924 20485
rect 26516 20476 26568 20528
rect 27988 20476 28040 20528
rect 28172 20476 28224 20528
rect 29828 20476 29880 20528
rect 33876 20519 33928 20528
rect 33876 20485 33885 20519
rect 33885 20485 33919 20519
rect 33919 20485 33928 20519
rect 33876 20476 33928 20485
rect 34704 20476 34756 20528
rect 35624 20476 35676 20528
rect 35992 20476 36044 20528
rect 27160 20451 27212 20460
rect 27160 20417 27169 20451
rect 27169 20417 27203 20451
rect 27203 20417 27212 20451
rect 27712 20451 27764 20460
rect 27160 20408 27212 20417
rect 27712 20417 27721 20451
rect 27721 20417 27755 20451
rect 27755 20417 27764 20451
rect 27712 20408 27764 20417
rect 27896 20451 27948 20460
rect 27896 20417 27905 20451
rect 27905 20417 27939 20451
rect 27939 20417 27948 20451
rect 27896 20408 27948 20417
rect 28540 20451 28592 20460
rect 28540 20417 28549 20451
rect 28549 20417 28583 20451
rect 28583 20417 28592 20451
rect 28540 20408 28592 20417
rect 31300 20451 31352 20460
rect 31300 20417 31309 20451
rect 31309 20417 31343 20451
rect 31343 20417 31352 20451
rect 31300 20408 31352 20417
rect 11520 20383 11572 20392
rect 11520 20349 11529 20383
rect 11529 20349 11563 20383
rect 11563 20349 11572 20383
rect 11520 20340 11572 20349
rect 12348 20340 12400 20392
rect 19432 20340 19484 20392
rect 22468 20383 22520 20392
rect 11888 20204 11940 20256
rect 19340 20272 19392 20324
rect 13728 20247 13780 20256
rect 13728 20213 13737 20247
rect 13737 20213 13771 20247
rect 13771 20213 13780 20247
rect 13728 20204 13780 20213
rect 16948 20247 17000 20256
rect 16948 20213 16957 20247
rect 16957 20213 16991 20247
rect 16991 20213 17000 20247
rect 16948 20204 17000 20213
rect 17224 20204 17276 20256
rect 18420 20204 18472 20256
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 22560 20340 22612 20392
rect 33692 20408 33744 20460
rect 43720 20476 43772 20528
rect 43904 20476 43956 20528
rect 45376 20519 45428 20528
rect 35440 20383 35492 20392
rect 35440 20349 35449 20383
rect 35449 20349 35483 20383
rect 35483 20349 35492 20383
rect 35440 20340 35492 20349
rect 42616 20408 42668 20460
rect 43076 20408 43128 20460
rect 45376 20485 45385 20519
rect 45385 20485 45419 20519
rect 45419 20485 45428 20519
rect 45376 20476 45428 20485
rect 46572 20408 46624 20460
rect 42708 20340 42760 20392
rect 42892 20383 42944 20392
rect 42892 20349 42901 20383
rect 42901 20349 42935 20383
rect 42935 20349 42944 20383
rect 42892 20340 42944 20349
rect 43536 20383 43588 20392
rect 43536 20349 43545 20383
rect 43545 20349 43579 20383
rect 43579 20349 43588 20383
rect 43536 20340 43588 20349
rect 46388 20383 46440 20392
rect 46388 20349 46397 20383
rect 46397 20349 46431 20383
rect 46431 20349 46440 20383
rect 46388 20340 46440 20349
rect 25044 20272 25096 20324
rect 25596 20315 25648 20324
rect 25596 20281 25605 20315
rect 25605 20281 25639 20315
rect 25639 20281 25648 20315
rect 25596 20272 25648 20281
rect 25780 20272 25832 20324
rect 27160 20272 27212 20324
rect 32220 20272 32272 20324
rect 42524 20272 42576 20324
rect 23756 20204 23808 20256
rect 25320 20204 25372 20256
rect 26332 20204 26384 20256
rect 31300 20204 31352 20256
rect 37464 20204 37516 20256
rect 42892 20204 42944 20256
rect 44180 20204 44232 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 11520 20000 11572 20052
rect 12348 20043 12400 20052
rect 12348 20009 12357 20043
rect 12357 20009 12391 20043
rect 12391 20009 12400 20043
rect 12348 20000 12400 20009
rect 15568 20043 15620 20052
rect 15568 20009 15577 20043
rect 15577 20009 15611 20043
rect 15611 20009 15620 20043
rect 15568 20000 15620 20009
rect 15844 20000 15896 20052
rect 20536 20000 20588 20052
rect 18512 19932 18564 19984
rect 22192 20000 22244 20052
rect 32496 20000 32548 20052
rect 25596 19932 25648 19984
rect 25964 19932 26016 19984
rect 36360 19932 36412 19984
rect 43812 20000 43864 20052
rect 43996 20043 44048 20052
rect 43996 20009 44005 20043
rect 44005 20009 44039 20043
rect 44039 20009 44048 20043
rect 43996 20000 44048 20009
rect 42524 19932 42576 19984
rect 46112 19932 46164 19984
rect 1768 19796 1820 19848
rect 11796 19839 11848 19848
rect 11796 19805 11805 19839
rect 11805 19805 11839 19839
rect 11839 19805 11848 19839
rect 11796 19796 11848 19805
rect 17224 19864 17276 19916
rect 18604 19864 18656 19916
rect 19156 19864 19208 19916
rect 20352 19907 20404 19916
rect 20352 19873 20361 19907
rect 20361 19873 20395 19907
rect 20395 19873 20404 19907
rect 20352 19864 20404 19873
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14372 19796 14424 19848
rect 16856 19796 16908 19848
rect 18696 19796 18748 19848
rect 19064 19796 19116 19848
rect 19984 19796 20036 19848
rect 25688 19839 25740 19848
rect 25688 19805 25697 19839
rect 25697 19805 25731 19839
rect 25731 19805 25740 19839
rect 25688 19796 25740 19805
rect 26240 19796 26292 19848
rect 32404 19839 32456 19848
rect 32404 19805 32413 19839
rect 32413 19805 32447 19839
rect 32447 19805 32456 19839
rect 32404 19796 32456 19805
rect 11888 19728 11940 19780
rect 15476 19728 15528 19780
rect 16764 19728 16816 19780
rect 17224 19771 17276 19780
rect 17224 19737 17233 19771
rect 17233 19737 17267 19771
rect 17267 19737 17276 19771
rect 17224 19728 17276 19737
rect 18972 19728 19024 19780
rect 19340 19771 19392 19780
rect 19340 19737 19349 19771
rect 19349 19737 19383 19771
rect 19383 19737 19392 19771
rect 19340 19728 19392 19737
rect 22560 19771 22612 19780
rect 13820 19660 13872 19712
rect 14188 19703 14240 19712
rect 14188 19669 14197 19703
rect 14197 19669 14231 19703
rect 14231 19669 14240 19703
rect 14188 19660 14240 19669
rect 15752 19703 15804 19712
rect 15752 19669 15761 19703
rect 15761 19669 15795 19703
rect 15795 19669 15804 19703
rect 15752 19660 15804 19669
rect 16396 19660 16448 19712
rect 18052 19660 18104 19712
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 18788 19660 18840 19712
rect 20260 19660 20312 19712
rect 22560 19737 22569 19771
rect 22569 19737 22603 19771
rect 22603 19737 22612 19771
rect 22560 19728 22612 19737
rect 25780 19728 25832 19780
rect 25872 19771 25924 19780
rect 25872 19737 25881 19771
rect 25881 19737 25915 19771
rect 25915 19737 25924 19771
rect 25872 19728 25924 19737
rect 22192 19660 22244 19712
rect 22376 19660 22428 19712
rect 26332 19728 26384 19780
rect 35440 19796 35492 19848
rect 36360 19728 36412 19780
rect 26516 19703 26568 19712
rect 26516 19669 26525 19703
rect 26525 19669 26559 19703
rect 26559 19669 26568 19703
rect 26516 19660 26568 19669
rect 26792 19660 26844 19712
rect 33232 19660 33284 19712
rect 33508 19660 33560 19712
rect 42708 19796 42760 19848
rect 42800 19839 42852 19848
rect 42800 19805 42809 19839
rect 42809 19805 42843 19839
rect 42843 19805 42852 19839
rect 42800 19796 42852 19805
rect 42616 19771 42668 19780
rect 42616 19737 42625 19771
rect 42625 19737 42659 19771
rect 42659 19737 42668 19771
rect 42616 19728 42668 19737
rect 43444 19660 43496 19712
rect 43720 19864 43772 19916
rect 43812 19864 43864 19916
rect 46572 19864 46624 19916
rect 43720 19728 43772 19780
rect 43904 19728 43956 19780
rect 47676 19728 47728 19780
rect 48136 19771 48188 19780
rect 48136 19737 48145 19771
rect 48145 19737 48179 19771
rect 48179 19737 48188 19771
rect 48136 19728 48188 19737
rect 45928 19660 45980 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3424 19456 3476 19508
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 13728 19388 13780 19440
rect 14188 19388 14240 19440
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 14096 19252 14148 19304
rect 14464 19252 14516 19304
rect 15568 19431 15620 19440
rect 15568 19397 15593 19431
rect 15593 19397 15620 19431
rect 15568 19388 15620 19397
rect 17224 19388 17276 19440
rect 13820 19116 13872 19168
rect 14188 19116 14240 19168
rect 15844 19320 15896 19372
rect 16764 19363 16816 19372
rect 16764 19329 16773 19363
rect 16773 19329 16807 19363
rect 16807 19329 16816 19363
rect 18788 19388 18840 19440
rect 19800 19388 19852 19440
rect 20168 19388 20220 19440
rect 16764 19320 16816 19329
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 18604 19320 18656 19372
rect 19064 19320 19116 19372
rect 19892 19363 19944 19372
rect 19892 19329 19901 19363
rect 19901 19329 19935 19363
rect 19935 19329 19944 19363
rect 19892 19320 19944 19329
rect 20536 19456 20588 19508
rect 43076 19499 43128 19508
rect 20628 19388 20680 19440
rect 20812 19320 20864 19372
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 22008 19431 22060 19440
rect 22008 19397 22033 19431
rect 22033 19397 22060 19431
rect 22008 19388 22060 19397
rect 22284 19388 22336 19440
rect 25872 19388 25924 19440
rect 21088 19320 21140 19329
rect 22192 19320 22244 19372
rect 23388 19320 23440 19372
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 23756 19320 23808 19329
rect 18972 19227 19024 19236
rect 18972 19193 18981 19227
rect 18981 19193 19015 19227
rect 19015 19193 19024 19227
rect 18972 19184 19024 19193
rect 20996 19184 21048 19236
rect 15476 19116 15528 19168
rect 16856 19159 16908 19168
rect 16856 19125 16865 19159
rect 16865 19125 16899 19159
rect 16899 19125 16908 19159
rect 16856 19116 16908 19125
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 26148 19431 26200 19440
rect 26148 19397 26173 19431
rect 26173 19397 26200 19431
rect 32220 19431 32272 19440
rect 26148 19388 26200 19397
rect 32220 19397 32229 19431
rect 32229 19397 32263 19431
rect 32263 19397 32272 19431
rect 32220 19388 32272 19397
rect 33324 19388 33376 19440
rect 33508 19431 33560 19440
rect 33508 19397 33517 19431
rect 33517 19397 33551 19431
rect 33551 19397 33560 19431
rect 33508 19388 33560 19397
rect 43076 19465 43085 19499
rect 43085 19465 43119 19499
rect 43119 19465 43128 19499
rect 43076 19456 43128 19465
rect 43444 19456 43496 19508
rect 42892 19388 42944 19440
rect 45008 19431 45060 19440
rect 26056 19320 26108 19372
rect 26792 19320 26844 19372
rect 42984 19363 43036 19372
rect 42984 19329 42993 19363
rect 42993 19329 43027 19363
rect 43027 19329 43036 19363
rect 42984 19320 43036 19329
rect 43168 19363 43220 19372
rect 43168 19329 43177 19363
rect 43177 19329 43211 19363
rect 43211 19329 43220 19363
rect 43168 19320 43220 19329
rect 43996 19363 44048 19372
rect 43996 19329 44005 19363
rect 44005 19329 44039 19363
rect 44039 19329 44048 19363
rect 43996 19320 44048 19329
rect 44272 19320 44324 19372
rect 45008 19397 45017 19431
rect 45017 19397 45051 19431
rect 45051 19397 45060 19431
rect 45008 19388 45060 19397
rect 45652 19456 45704 19508
rect 47676 19499 47728 19508
rect 47676 19465 47685 19499
rect 47685 19465 47719 19499
rect 47719 19465 47728 19499
rect 47676 19456 47728 19465
rect 46756 19388 46808 19440
rect 45744 19363 45796 19372
rect 26516 19252 26568 19304
rect 32496 19295 32548 19304
rect 32496 19261 32505 19295
rect 32505 19261 32539 19295
rect 32539 19261 32548 19295
rect 32496 19252 32548 19261
rect 33232 19252 33284 19304
rect 45744 19329 45753 19363
rect 45753 19329 45787 19363
rect 45787 19329 45796 19363
rect 45744 19320 45796 19329
rect 47492 19320 47544 19372
rect 26332 19227 26384 19236
rect 26332 19193 26341 19227
rect 26341 19193 26375 19227
rect 26375 19193 26384 19227
rect 26332 19184 26384 19193
rect 25320 19116 25372 19168
rect 25504 19159 25556 19168
rect 25504 19125 25513 19159
rect 25513 19125 25547 19159
rect 25547 19125 25556 19159
rect 25504 19116 25556 19125
rect 46296 19116 46348 19168
rect 46940 19159 46992 19168
rect 46940 19125 46949 19159
rect 46949 19125 46983 19159
rect 46983 19125 46992 19159
rect 46940 19116 46992 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 14464 18912 14516 18964
rect 21088 18912 21140 18964
rect 25872 18912 25924 18964
rect 29828 18912 29880 18964
rect 30288 18912 30340 18964
rect 32404 18912 32456 18964
rect 32588 18955 32640 18964
rect 32588 18921 32597 18955
rect 32597 18921 32631 18955
rect 32631 18921 32640 18955
rect 32588 18912 32640 18921
rect 33324 18955 33376 18964
rect 33324 18921 33333 18955
rect 33333 18921 33367 18955
rect 33367 18921 33376 18955
rect 33324 18912 33376 18921
rect 45836 18955 45888 18964
rect 45836 18921 45845 18955
rect 45845 18921 45879 18955
rect 45879 18921 45888 18955
rect 45836 18912 45888 18921
rect 13544 18844 13596 18896
rect 4896 18776 4948 18828
rect 2320 18708 2372 18760
rect 13636 18708 13688 18760
rect 14188 18751 14240 18760
rect 14188 18717 14230 18751
rect 14230 18717 14240 18751
rect 14188 18708 14240 18717
rect 15200 18776 15252 18828
rect 15752 18776 15804 18828
rect 15476 18708 15528 18760
rect 16856 18844 16908 18896
rect 19892 18844 19944 18896
rect 20996 18844 21048 18896
rect 20720 18776 20772 18828
rect 22100 18844 22152 18896
rect 25228 18844 25280 18896
rect 25780 18844 25832 18896
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 16304 18751 16356 18760
rect 16304 18717 16313 18751
rect 16313 18717 16347 18751
rect 16347 18717 16356 18751
rect 16304 18708 16356 18717
rect 17960 18708 18012 18760
rect 20904 18708 20956 18760
rect 21916 18708 21968 18760
rect 22100 18708 22152 18760
rect 23388 18708 23440 18760
rect 25044 18640 25096 18692
rect 25320 18708 25372 18760
rect 25780 18708 25832 18760
rect 26884 18751 26936 18760
rect 26884 18717 26893 18751
rect 26893 18717 26927 18751
rect 26927 18717 26936 18751
rect 26884 18708 26936 18717
rect 13084 18572 13136 18624
rect 13544 18572 13596 18624
rect 15384 18572 15436 18624
rect 15568 18615 15620 18624
rect 15568 18581 15577 18615
rect 15577 18581 15611 18615
rect 15611 18581 15620 18615
rect 15568 18572 15620 18581
rect 15660 18572 15712 18624
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 25228 18615 25280 18624
rect 25504 18640 25556 18692
rect 28724 18708 28776 18760
rect 32496 18844 32548 18896
rect 33232 18844 33284 18896
rect 30288 18708 30340 18760
rect 31392 18776 31444 18828
rect 46756 18844 46808 18896
rect 29184 18640 29236 18692
rect 25228 18581 25243 18615
rect 25243 18581 25277 18615
rect 25277 18581 25280 18615
rect 25228 18572 25280 18581
rect 25872 18572 25924 18624
rect 29092 18572 29144 18624
rect 35072 18776 35124 18828
rect 46112 18776 46164 18828
rect 46296 18819 46348 18828
rect 46296 18785 46305 18819
rect 46305 18785 46339 18819
rect 46339 18785 46348 18819
rect 46296 18776 46348 18785
rect 46940 18776 46992 18828
rect 45836 18708 45888 18760
rect 35440 18640 35492 18692
rect 36544 18683 36596 18692
rect 36544 18649 36553 18683
rect 36553 18649 36587 18683
rect 36587 18649 36596 18683
rect 36544 18640 36596 18649
rect 45376 18640 45428 18692
rect 47860 18640 47912 18692
rect 45560 18615 45612 18624
rect 45560 18581 45569 18615
rect 45569 18581 45603 18615
rect 45603 18581 45612 18615
rect 45560 18572 45612 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3976 18368 4028 18420
rect 15200 18300 15252 18352
rect 17684 18343 17736 18352
rect 17684 18309 17693 18343
rect 17693 18309 17727 18343
rect 17727 18309 17736 18343
rect 17684 18300 17736 18309
rect 21548 18300 21600 18352
rect 22744 18300 22796 18352
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 11428 18232 11480 18284
rect 12256 18232 12308 18284
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 15476 18232 15528 18284
rect 25872 18300 25924 18352
rect 35716 18368 35768 18420
rect 45560 18368 45612 18420
rect 25228 18232 25280 18284
rect 26056 18232 26108 18284
rect 29000 18275 29052 18284
rect 29000 18241 29009 18275
rect 29009 18241 29043 18275
rect 29043 18241 29052 18275
rect 29000 18232 29052 18241
rect 29460 18232 29512 18284
rect 35072 18275 35124 18284
rect 35072 18241 35081 18275
rect 35081 18241 35115 18275
rect 35115 18241 35124 18275
rect 35072 18232 35124 18241
rect 35440 18232 35492 18284
rect 38108 18232 38160 18284
rect 45376 18232 45428 18284
rect 45836 18275 45888 18284
rect 45836 18241 45845 18275
rect 45845 18241 45879 18275
rect 45879 18241 45888 18275
rect 45836 18232 45888 18241
rect 46112 18275 46164 18284
rect 46112 18241 46121 18275
rect 46121 18241 46155 18275
rect 46155 18241 46164 18275
rect 46112 18232 46164 18241
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 16304 18164 16356 18216
rect 17132 18164 17184 18216
rect 19156 18207 19208 18216
rect 19156 18173 19165 18207
rect 19165 18173 19199 18207
rect 19199 18173 19208 18207
rect 19156 18164 19208 18173
rect 15384 18139 15436 18148
rect 11888 18028 11940 18080
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 14464 18071 14516 18080
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 14464 18028 14516 18037
rect 15384 18105 15393 18139
rect 15393 18105 15427 18139
rect 15427 18105 15436 18139
rect 15384 18096 15436 18105
rect 17040 18028 17092 18080
rect 22100 18164 22152 18216
rect 23848 18207 23900 18216
rect 23848 18173 23857 18207
rect 23857 18173 23891 18207
rect 23891 18173 23900 18207
rect 23848 18164 23900 18173
rect 25044 18164 25096 18216
rect 26516 18164 26568 18216
rect 26792 18164 26844 18216
rect 31208 18164 31260 18216
rect 30656 18096 30708 18148
rect 33876 18164 33928 18216
rect 32864 18096 32916 18148
rect 36544 18164 36596 18216
rect 43536 18164 43588 18216
rect 43904 18207 43956 18216
rect 43904 18173 43913 18207
rect 43913 18173 43947 18207
rect 43947 18173 43956 18207
rect 43904 18164 43956 18173
rect 46204 18164 46256 18216
rect 47400 18232 47452 18284
rect 34520 18096 34572 18148
rect 48044 18164 48096 18216
rect 22100 18028 22152 18080
rect 25044 18071 25096 18080
rect 25044 18037 25053 18071
rect 25053 18037 25087 18071
rect 25087 18037 25096 18071
rect 25044 18028 25096 18037
rect 25320 18028 25372 18080
rect 29736 18028 29788 18080
rect 35348 18071 35400 18080
rect 35348 18037 35357 18071
rect 35357 18037 35391 18071
rect 35391 18037 35400 18071
rect 45560 18071 45612 18080
rect 35348 18028 35400 18037
rect 45560 18037 45569 18071
rect 45569 18037 45603 18071
rect 45603 18037 45612 18071
rect 45560 18028 45612 18037
rect 47032 18071 47084 18080
rect 47032 18037 47041 18071
rect 47041 18037 47075 18071
rect 47075 18037 47084 18071
rect 47032 18028 47084 18037
rect 47676 18071 47728 18080
rect 47676 18037 47685 18071
rect 47685 18037 47719 18071
rect 47719 18037 47728 18071
rect 47676 18028 47728 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3976 17756 4028 17808
rect 11612 17688 11664 17740
rect 11888 17731 11940 17740
rect 11888 17697 11897 17731
rect 11897 17697 11931 17731
rect 11931 17697 11940 17731
rect 11888 17688 11940 17697
rect 12256 17688 12308 17740
rect 16672 17824 16724 17876
rect 17132 17867 17184 17876
rect 17132 17833 17141 17867
rect 17141 17833 17175 17867
rect 17175 17833 17184 17867
rect 17132 17824 17184 17833
rect 22100 17867 22152 17876
rect 22100 17833 22109 17867
rect 22109 17833 22143 17867
rect 22143 17833 22152 17867
rect 22744 17867 22796 17876
rect 22100 17824 22152 17833
rect 22744 17833 22753 17867
rect 22753 17833 22787 17867
rect 22787 17833 22796 17867
rect 22744 17824 22796 17833
rect 26792 17867 26844 17876
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 16764 17620 16816 17672
rect 18880 17688 18932 17740
rect 22376 17688 22428 17740
rect 17868 17620 17920 17672
rect 21180 17620 21232 17672
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 24400 17663 24452 17672
rect 24400 17629 24409 17663
rect 24409 17629 24443 17663
rect 24443 17629 24452 17663
rect 26792 17833 26801 17867
rect 26801 17833 26835 17867
rect 26835 17833 26844 17867
rect 26792 17824 26844 17833
rect 31208 17867 31260 17876
rect 31208 17833 31217 17867
rect 31217 17833 31251 17867
rect 31251 17833 31260 17867
rect 31208 17824 31260 17833
rect 33876 17867 33928 17876
rect 33876 17833 33885 17867
rect 33885 17833 33919 17867
rect 33919 17833 33928 17867
rect 33876 17824 33928 17833
rect 35716 17824 35768 17876
rect 43996 17824 44048 17876
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 25320 17731 25372 17740
rect 25320 17697 25329 17731
rect 25329 17697 25363 17731
rect 25363 17697 25372 17731
rect 25320 17688 25372 17697
rect 28724 17731 28776 17740
rect 28724 17697 28733 17731
rect 28733 17697 28767 17731
rect 28767 17697 28776 17731
rect 28724 17688 28776 17697
rect 29828 17731 29880 17740
rect 29828 17697 29837 17731
rect 29837 17697 29871 17731
rect 29871 17697 29880 17731
rect 30656 17731 30708 17740
rect 29828 17688 29880 17697
rect 30656 17697 30665 17731
rect 30665 17697 30699 17731
rect 30699 17697 30708 17731
rect 30656 17688 30708 17697
rect 35072 17756 35124 17808
rect 44640 17756 44692 17808
rect 28356 17663 28408 17672
rect 24400 17620 24452 17629
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 28540 17620 28592 17672
rect 29184 17620 29236 17672
rect 29736 17620 29788 17672
rect 31116 17663 31168 17672
rect 31116 17629 31125 17663
rect 31125 17629 31159 17663
rect 31159 17629 31168 17663
rect 31116 17620 31168 17629
rect 34520 17620 34572 17672
rect 35348 17663 35400 17672
rect 19432 17552 19484 17604
rect 20168 17552 20220 17604
rect 26056 17552 26108 17604
rect 35348 17629 35357 17663
rect 35357 17629 35391 17663
rect 35391 17629 35400 17663
rect 35348 17620 35400 17629
rect 35440 17663 35492 17672
rect 35440 17629 35449 17663
rect 35449 17629 35483 17663
rect 35483 17629 35492 17663
rect 47032 17688 47084 17740
rect 35440 17620 35492 17629
rect 45376 17663 45428 17672
rect 45376 17629 45385 17663
rect 45385 17629 45419 17663
rect 45419 17629 45428 17663
rect 45376 17620 45428 17629
rect 35716 17552 35768 17604
rect 44088 17595 44140 17604
rect 44088 17561 44097 17595
rect 44097 17561 44131 17595
rect 44131 17561 44140 17595
rect 44088 17552 44140 17561
rect 20996 17527 21048 17536
rect 20996 17493 21005 17527
rect 21005 17493 21039 17527
rect 21039 17493 21048 17527
rect 20996 17484 21048 17493
rect 23664 17484 23716 17536
rect 28632 17484 28684 17536
rect 28816 17484 28868 17536
rect 31116 17484 31168 17536
rect 39212 17484 39264 17536
rect 43628 17527 43680 17536
rect 43628 17493 43637 17527
rect 43637 17493 43671 17527
rect 43671 17493 43680 17527
rect 43628 17484 43680 17493
rect 45284 17552 45336 17604
rect 45652 17620 45704 17672
rect 47676 17552 47728 17604
rect 48228 17552 48280 17604
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 5448 17280 5500 17332
rect 16764 17323 16816 17332
rect 13360 17212 13412 17264
rect 14464 17212 14516 17264
rect 12256 17144 12308 17196
rect 14188 17076 14240 17128
rect 1400 16940 1452 16992
rect 11888 16940 11940 16992
rect 12992 16940 13044 16992
rect 15568 16940 15620 16992
rect 16764 17289 16773 17323
rect 16773 17289 16807 17323
rect 16807 17289 16816 17323
rect 16764 17280 16816 17289
rect 17868 17323 17920 17332
rect 17868 17289 17877 17323
rect 17877 17289 17911 17323
rect 17911 17289 17920 17323
rect 17868 17280 17920 17289
rect 20076 17280 20128 17332
rect 26056 17280 26108 17332
rect 28724 17323 28776 17332
rect 28724 17289 28733 17323
rect 28733 17289 28767 17323
rect 28767 17289 28776 17323
rect 28724 17280 28776 17289
rect 28816 17280 28868 17332
rect 16948 17212 17000 17264
rect 20352 17212 20404 17264
rect 23664 17255 23716 17264
rect 16764 17144 16816 17196
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 23664 17221 23673 17255
rect 23673 17221 23707 17255
rect 23707 17221 23716 17255
rect 23664 17212 23716 17221
rect 23848 17212 23900 17264
rect 27896 17212 27948 17264
rect 28632 17255 28684 17264
rect 28632 17221 28641 17255
rect 28641 17221 28675 17255
rect 28675 17221 28684 17255
rect 28632 17212 28684 17221
rect 22376 17144 22428 17196
rect 23388 17144 23440 17196
rect 25780 17144 25832 17196
rect 26056 17187 26108 17196
rect 26056 17153 26065 17187
rect 26065 17153 26099 17187
rect 26099 17153 26108 17187
rect 26056 17144 26108 17153
rect 27528 17187 27580 17196
rect 18512 17119 18564 17128
rect 18512 17085 18521 17119
rect 18521 17085 18555 17119
rect 18555 17085 18564 17119
rect 18512 17076 18564 17085
rect 19340 17076 19392 17128
rect 19984 17076 20036 17128
rect 20352 17076 20404 17128
rect 20720 17076 20772 17128
rect 25320 17119 25372 17128
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 27528 17153 27537 17187
rect 27537 17153 27571 17187
rect 27571 17153 27580 17187
rect 27528 17144 27580 17153
rect 27712 17187 27764 17196
rect 27712 17153 27721 17187
rect 27721 17153 27755 17187
rect 27755 17153 27764 17187
rect 27712 17144 27764 17153
rect 29092 17144 29144 17196
rect 36544 17280 36596 17332
rect 41880 17280 41932 17332
rect 45744 17280 45796 17332
rect 35072 17255 35124 17264
rect 35072 17221 35081 17255
rect 35081 17221 35115 17255
rect 35115 17221 35124 17255
rect 35072 17212 35124 17221
rect 44272 17255 44324 17264
rect 44272 17221 44281 17255
rect 44281 17221 44315 17255
rect 44315 17221 44324 17255
rect 44272 17212 44324 17221
rect 45560 17212 45612 17264
rect 29460 17119 29512 17128
rect 29460 17085 29469 17119
rect 29469 17085 29503 17119
rect 29503 17085 29512 17119
rect 29460 17076 29512 17085
rect 43628 17144 43680 17196
rect 47584 17187 47636 17196
rect 47584 17153 47593 17187
rect 47593 17153 47627 17187
rect 47627 17153 47636 17187
rect 47584 17144 47636 17153
rect 30656 17076 30708 17128
rect 36544 17119 36596 17128
rect 36544 17085 36553 17119
rect 36553 17085 36587 17119
rect 36587 17085 36596 17119
rect 36544 17076 36596 17085
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 21364 16940 21416 16992
rect 24860 16940 24912 16992
rect 25044 16940 25096 16992
rect 28724 16940 28776 16992
rect 29460 16940 29512 16992
rect 29828 16983 29880 16992
rect 29828 16949 29837 16983
rect 29837 16949 29871 16983
rect 29871 16949 29880 16983
rect 29828 16940 29880 16949
rect 30380 16983 30432 16992
rect 30380 16949 30389 16983
rect 30389 16949 30423 16983
rect 30423 16949 30432 16983
rect 30380 16940 30432 16949
rect 42524 17008 42576 17060
rect 45284 17076 45336 17128
rect 45744 17119 45796 17128
rect 45744 17085 45753 17119
rect 45753 17085 45787 17119
rect 45787 17085 45796 17119
rect 45744 17076 45796 17085
rect 47676 16983 47728 16992
rect 47676 16949 47685 16983
rect 47685 16949 47719 16983
rect 47719 16949 47728 16983
rect 47676 16940 47728 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 18512 16736 18564 16788
rect 19432 16736 19484 16788
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25044 16779 25096 16788
rect 25044 16745 25053 16779
rect 25053 16745 25087 16779
rect 25087 16745 25096 16779
rect 25044 16736 25096 16745
rect 25780 16736 25832 16788
rect 29000 16736 29052 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 12992 16668 13044 16720
rect 20260 16668 20312 16720
rect 23664 16668 23716 16720
rect 29092 16668 29144 16720
rect 11888 16643 11940 16652
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 12440 16600 12492 16609
rect 16672 16600 16724 16652
rect 17684 16600 17736 16652
rect 14188 16575 14240 16584
rect 14188 16541 14197 16575
rect 14197 16541 14231 16575
rect 14231 16541 14240 16575
rect 16212 16575 16264 16584
rect 14188 16532 14240 16541
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 20076 16600 20128 16652
rect 20352 16600 20404 16652
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 2136 16464 2188 16516
rect 20720 16532 20772 16584
rect 24400 16600 24452 16652
rect 27528 16600 27580 16652
rect 24860 16532 24912 16584
rect 20996 16464 21048 16516
rect 23388 16464 23440 16516
rect 23572 16464 23624 16516
rect 25596 16532 25648 16584
rect 25780 16532 25832 16584
rect 27712 16600 27764 16652
rect 27896 16600 27948 16652
rect 30656 16643 30708 16652
rect 30656 16609 30665 16643
rect 30665 16609 30699 16643
rect 30699 16609 30708 16643
rect 30656 16600 30708 16609
rect 44088 16668 44140 16720
rect 28356 16532 28408 16584
rect 29644 16575 29696 16584
rect 29644 16541 29653 16575
rect 29653 16541 29687 16575
rect 29687 16541 29696 16575
rect 29644 16532 29696 16541
rect 29828 16575 29880 16584
rect 29828 16541 29837 16575
rect 29837 16541 29871 16575
rect 29871 16541 29880 16575
rect 29828 16532 29880 16541
rect 46572 16668 46624 16720
rect 45652 16600 45704 16652
rect 47768 16600 47820 16652
rect 48136 16643 48188 16652
rect 48136 16609 48145 16643
rect 48145 16609 48179 16643
rect 48179 16609 48188 16643
rect 48136 16600 48188 16609
rect 25872 16464 25924 16516
rect 28540 16464 28592 16516
rect 28632 16507 28684 16516
rect 28632 16473 28641 16507
rect 28641 16473 28675 16507
rect 28675 16473 28684 16507
rect 32496 16507 32548 16516
rect 28632 16464 28684 16473
rect 32496 16473 32505 16507
rect 32505 16473 32539 16507
rect 32539 16473 32548 16507
rect 32496 16464 32548 16473
rect 42800 16464 42852 16516
rect 45376 16464 45428 16516
rect 47676 16464 47728 16516
rect 16304 16439 16356 16448
rect 16304 16405 16313 16439
rect 16313 16405 16347 16439
rect 16347 16405 16356 16439
rect 16304 16396 16356 16405
rect 20076 16396 20128 16448
rect 20904 16396 20956 16448
rect 23848 16396 23900 16448
rect 25596 16396 25648 16448
rect 25964 16396 26016 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 20168 16124 20220 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 16212 16056 16264 16108
rect 22744 16192 22796 16244
rect 23572 16235 23624 16244
rect 23572 16201 23581 16235
rect 23581 16201 23615 16235
rect 23615 16201 23624 16235
rect 23572 16192 23624 16201
rect 25872 16235 25924 16244
rect 25872 16201 25881 16235
rect 25881 16201 25915 16235
rect 25915 16201 25924 16235
rect 25872 16192 25924 16201
rect 28724 16192 28776 16244
rect 29644 16192 29696 16244
rect 32496 16192 32548 16244
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 22192 16124 22244 16176
rect 23112 16124 23164 16176
rect 25964 16124 26016 16176
rect 21180 16099 21232 16108
rect 21180 16065 21189 16099
rect 21189 16065 21223 16099
rect 21223 16065 21232 16099
rect 21180 16056 21232 16065
rect 26148 16056 26200 16108
rect 28540 16056 28592 16108
rect 28632 16099 28684 16108
rect 28632 16065 28641 16099
rect 28641 16065 28675 16099
rect 28675 16065 28684 16099
rect 29092 16099 29144 16108
rect 28632 16056 28684 16065
rect 29092 16065 29101 16099
rect 29101 16065 29135 16099
rect 29135 16065 29144 16099
rect 29092 16056 29144 16065
rect 30380 16056 30432 16108
rect 32772 16056 32824 16108
rect 44272 16124 44324 16176
rect 47768 16099 47820 16108
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 24124 16031 24176 16040
rect 22100 15988 22152 15997
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 24860 15988 24912 16040
rect 44180 16031 44232 16040
rect 44180 15997 44189 16031
rect 44189 15997 44223 16031
rect 44223 15997 44232 16031
rect 44180 15988 44232 15997
rect 45836 16031 45888 16040
rect 45836 15997 45845 16031
rect 45845 15997 45879 16031
rect 45879 15997 45888 16031
rect 45836 15988 45888 15997
rect 21272 15852 21324 15904
rect 22192 15852 22244 15904
rect 26792 15852 26844 15904
rect 27160 15852 27212 15904
rect 30564 15852 30616 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19340 15648 19392 15700
rect 22100 15648 22152 15700
rect 23112 15648 23164 15700
rect 23388 15648 23440 15700
rect 24860 15691 24912 15700
rect 3516 15580 3568 15632
rect 16304 15555 16356 15564
rect 16304 15521 16313 15555
rect 16313 15521 16347 15555
rect 16347 15521 16356 15555
rect 16304 15512 16356 15521
rect 1768 15444 1820 15496
rect 20076 15512 20128 15564
rect 23572 15580 23624 15632
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 44180 15648 44232 15700
rect 45560 15580 45612 15632
rect 20260 15444 20312 15496
rect 20720 15444 20772 15496
rect 24124 15512 24176 15564
rect 24676 15555 24728 15564
rect 24676 15521 24685 15555
rect 24685 15521 24719 15555
rect 24719 15521 24728 15555
rect 24676 15512 24728 15521
rect 30564 15555 30616 15564
rect 22744 15444 22796 15496
rect 23664 15376 23716 15428
rect 21180 15308 21232 15360
rect 23940 15444 23992 15496
rect 24768 15444 24820 15496
rect 25228 15376 25280 15428
rect 25780 15444 25832 15496
rect 26056 15376 26108 15428
rect 25688 15308 25740 15360
rect 26608 15376 26660 15428
rect 27160 15376 27212 15428
rect 30564 15521 30573 15555
rect 30573 15521 30607 15555
rect 30607 15521 30616 15555
rect 30564 15512 30616 15521
rect 30656 15512 30708 15564
rect 43812 15444 43864 15496
rect 43996 15487 44048 15496
rect 43996 15453 44005 15487
rect 44005 15453 44039 15487
rect 44039 15453 44048 15487
rect 43996 15444 44048 15453
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 25964 15147 26016 15156
rect 25964 15113 25973 15147
rect 25973 15113 26007 15147
rect 26007 15113 26016 15147
rect 25964 15104 26016 15113
rect 26608 15104 26660 15156
rect 23848 15036 23900 15088
rect 25688 15036 25740 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 26148 14968 26200 15020
rect 42524 14968 42576 15020
rect 2320 14900 2372 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 23940 14900 23992 14952
rect 43812 14943 43864 14952
rect 14740 14832 14792 14884
rect 43812 14909 43821 14943
rect 43821 14909 43855 14943
rect 43855 14909 43864 14943
rect 43812 14900 43864 14909
rect 45100 14943 45152 14952
rect 45100 14909 45109 14943
rect 45109 14909 45143 14943
rect 45143 14909 45152 14943
rect 45100 14900 45152 14909
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 24676 14560 24728 14612
rect 43812 14603 43864 14612
rect 43812 14569 43821 14603
rect 43821 14569 43855 14603
rect 43855 14569 43864 14603
rect 43812 14560 43864 14569
rect 2688 14356 2740 14408
rect 25228 14424 25280 14476
rect 25780 14356 25832 14408
rect 43996 14356 44048 14408
rect 33876 14288 33928 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 43996 13880 44048 13932
rect 3976 13744 4028 13796
rect 15292 13744 15344 13796
rect 47676 13719 47728 13728
rect 47676 13685 47685 13719
rect 47685 13685 47719 13719
rect 47719 13685 47728 13719
rect 47676 13676 47728 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 47676 13336 47728 13388
rect 46296 13311 46348 13320
rect 46296 13277 46305 13311
rect 46305 13277 46339 13311
rect 46339 13277 46348 13311
rect 46296 13268 46348 13277
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 46296 12792 46348 12844
rect 29368 12588 29420 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 47676 11135 47728 11144
rect 47676 11101 47685 11135
rect 47685 11101 47719 11135
rect 47719 11101 47728 11135
rect 47676 11092 47728 11101
rect 4068 10956 4120 11008
rect 12440 10956 12492 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 27620 10684 27672 10736
rect 27804 10684 27856 10736
rect 47492 10616 47544 10668
rect 46480 10412 46532 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 25504 10072 25556 10124
rect 26148 10115 26200 10124
rect 26148 10081 26157 10115
rect 26157 10081 26191 10115
rect 26191 10081 26200 10115
rect 26148 10072 26200 10081
rect 47676 10140 47728 10192
rect 46480 10115 46532 10124
rect 46480 10081 46489 10115
rect 46489 10081 46523 10115
rect 46523 10081 46532 10115
rect 46480 10072 46532 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 24584 9979 24636 9988
rect 24584 9945 24593 9979
rect 24593 9945 24627 9979
rect 24627 9945 24636 9979
rect 24584 9936 24636 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 24584 9707 24636 9716
rect 24584 9673 24593 9707
rect 24593 9673 24627 9707
rect 24627 9673 24636 9707
rect 24584 9664 24636 9673
rect 24400 9528 24452 9580
rect 38936 9528 38988 9580
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 46664 9392 46716 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47768 8891 47820 8900
rect 47768 8857 47777 8891
rect 47777 8857 47811 8891
rect 47811 8857 47820 8891
rect 47768 8848 47820 8857
rect 27344 8780 27396 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 44824 8619 44876 8628
rect 44824 8585 44833 8619
rect 44833 8585 44867 8619
rect 44867 8585 44876 8619
rect 44824 8576 44876 8585
rect 45560 8440 45612 8492
rect 44824 8236 44876 8288
rect 45652 8279 45704 8288
rect 45652 8245 45661 8279
rect 45661 8245 45695 8279
rect 45695 8245 45704 8279
rect 45652 8236 45704 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 42800 8032 42852 8084
rect 46848 8032 46900 8084
rect 46572 7939 46624 7948
rect 46572 7905 46581 7939
rect 46581 7905 46615 7939
rect 46615 7905 46624 7939
rect 46572 7896 46624 7905
rect 45652 7828 45704 7880
rect 45928 7803 45980 7812
rect 45928 7769 45937 7803
rect 45937 7769 45971 7803
rect 45971 7769 45980 7803
rect 45928 7760 45980 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 45928 7488 45980 7540
rect 45652 7463 45704 7472
rect 45652 7429 45661 7463
rect 45661 7429 45695 7463
rect 45695 7429 45704 7463
rect 45652 7420 45704 7429
rect 46572 7463 46624 7472
rect 46572 7429 46581 7463
rect 46581 7429 46615 7463
rect 46615 7429 46624 7463
rect 46572 7420 46624 7429
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 45560 7327 45612 7336
rect 45560 7293 45569 7327
rect 45569 7293 45603 7327
rect 45603 7293 45612 7327
rect 45560 7284 45612 7293
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4068 6808 4120 6860
rect 18512 6808 18564 6860
rect 42340 6851 42392 6860
rect 42340 6817 42349 6851
rect 42349 6817 42383 6851
rect 42383 6817 42392 6851
rect 42340 6808 42392 6817
rect 47308 6851 47360 6860
rect 47308 6817 47317 6851
rect 47317 6817 47351 6851
rect 47351 6817 47360 6851
rect 47308 6808 47360 6817
rect 46020 6740 46072 6792
rect 3976 6604 4028 6656
rect 41420 6715 41472 6724
rect 41420 6681 41429 6715
rect 41429 6681 41463 6715
rect 41463 6681 41472 6715
rect 41420 6672 41472 6681
rect 42616 6604 42668 6656
rect 45560 6604 45612 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 41420 6400 41472 6452
rect 43812 6400 43864 6452
rect 44180 6332 44232 6384
rect 41328 6264 41380 6316
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 41604 6196 41656 6248
rect 42616 6196 42668 6248
rect 42340 6128 42392 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 38476 5856 38528 5908
rect 41328 5899 41380 5908
rect 41328 5865 41337 5899
rect 41337 5865 41371 5899
rect 41371 5865 41380 5899
rect 41328 5856 41380 5865
rect 44180 5652 44232 5704
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 6644 5108 6696 5160
rect 37464 5287 37516 5296
rect 37464 5253 37473 5287
rect 37473 5253 37507 5287
rect 37507 5253 37516 5287
rect 37464 5244 37516 5253
rect 41328 5176 41380 5228
rect 47768 5219 47820 5228
rect 47768 5185 47777 5219
rect 47777 5185 47811 5219
rect 47811 5185 47820 5219
rect 47768 5176 47820 5185
rect 38384 5151 38436 5160
rect 38384 5117 38393 5151
rect 38393 5117 38427 5151
rect 38427 5117 38436 5151
rect 38384 5108 38436 5117
rect 23480 5040 23532 5092
rect 39120 4972 39172 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 20444 4700 20496 4752
rect 28632 4700 28684 4752
rect 45652 4700 45704 4752
rect 7656 4564 7708 4616
rect 31116 4632 31168 4684
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 16672 4564 16724 4616
rect 20260 4564 20312 4616
rect 21088 4607 21140 4616
rect 21088 4573 21097 4607
rect 21097 4573 21131 4607
rect 21131 4573 21140 4607
rect 21088 4564 21140 4573
rect 22468 4607 22520 4616
rect 22468 4573 22477 4607
rect 22477 4573 22511 4607
rect 22511 4573 22520 4607
rect 22468 4564 22520 4573
rect 39120 4607 39172 4616
rect 39120 4573 39129 4607
rect 39129 4573 39163 4607
rect 39163 4573 39172 4607
rect 39120 4564 39172 4573
rect 47492 4632 47544 4684
rect 46848 4564 46900 4616
rect 16856 4496 16908 4548
rect 40040 4539 40092 4548
rect 40040 4505 40049 4539
rect 40049 4505 40083 4539
rect 40083 4505 40092 4539
rect 40040 4496 40092 4505
rect 41696 4539 41748 4548
rect 41696 4505 41705 4539
rect 41705 4505 41739 4539
rect 41739 4505 41748 4539
rect 41696 4496 41748 4505
rect 42248 4496 42300 4548
rect 8300 4428 8352 4480
rect 17316 4428 17368 4480
rect 21732 4428 21784 4480
rect 22284 4428 22336 4480
rect 22652 4428 22704 4480
rect 45744 4428 45796 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 21088 4224 21140 4276
rect 22468 4224 22520 4276
rect 40040 4224 40092 4276
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 8300 4020 8352 4072
rect 4068 3952 4120 4004
rect 1584 3884 1636 3936
rect 2780 3884 2832 3936
rect 7104 3884 7156 3936
rect 13636 4088 13688 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 14924 4088 14976 4140
rect 15200 4088 15252 4140
rect 16948 4156 17000 4208
rect 17132 4156 17184 4208
rect 16764 4088 16816 4140
rect 19156 4156 19208 4208
rect 21456 4156 21508 4208
rect 27620 4199 27672 4208
rect 27620 4165 27629 4199
rect 27629 4165 27663 4199
rect 27663 4165 27672 4199
rect 27620 4156 27672 4165
rect 37372 4199 37424 4208
rect 37372 4165 37381 4199
rect 37381 4165 37415 4199
rect 37415 4165 37424 4199
rect 37372 4156 37424 4165
rect 37556 4156 37608 4208
rect 38384 4199 38436 4208
rect 38384 4165 38393 4199
rect 38393 4165 38427 4199
rect 38427 4165 38436 4199
rect 38384 4156 38436 4165
rect 40224 4156 40276 4208
rect 46388 4156 46440 4208
rect 46756 4156 46808 4208
rect 17960 4131 18012 4140
rect 17960 4097 17969 4131
rect 17969 4097 18003 4131
rect 18003 4097 18012 4131
rect 17960 4088 18012 4097
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 19340 4088 19392 4140
rect 20812 4088 20864 4140
rect 21916 4088 21968 4140
rect 22284 4088 22336 4140
rect 25136 4088 25188 4140
rect 25228 4088 25280 4140
rect 17132 3952 17184 4004
rect 25320 4020 25372 4072
rect 31392 4088 31444 4140
rect 36728 4131 36780 4140
rect 36728 4097 36737 4131
rect 36737 4097 36771 4131
rect 36771 4097 36780 4131
rect 36728 4088 36780 4097
rect 39120 4131 39172 4140
rect 39120 4097 39129 4131
rect 39129 4097 39163 4131
rect 39163 4097 39172 4131
rect 39120 4088 39172 4097
rect 39856 4088 39908 4140
rect 28540 4063 28592 4072
rect 28540 4029 28549 4063
rect 28549 4029 28583 4063
rect 28583 4029 28592 4063
rect 28540 4020 28592 4029
rect 38016 4020 38068 4072
rect 41328 4131 41380 4140
rect 41328 4097 41337 4131
rect 41337 4097 41371 4131
rect 41371 4097 41380 4131
rect 42432 4131 42484 4140
rect 41328 4088 41380 4097
rect 42432 4097 42441 4131
rect 42441 4097 42475 4131
rect 42475 4097 42484 4131
rect 42432 4088 42484 4097
rect 9220 3884 9272 3936
rect 11704 3884 11756 3936
rect 14280 3884 14332 3936
rect 14832 3884 14884 3936
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15476 3884 15528 3936
rect 16580 3884 16632 3936
rect 17224 3884 17276 3936
rect 17868 3884 17920 3936
rect 18512 3884 18564 3936
rect 18788 3884 18840 3936
rect 20536 3884 20588 3936
rect 20628 3927 20680 3936
rect 20628 3893 20637 3927
rect 20637 3893 20671 3927
rect 20671 3893 20680 3927
rect 20628 3884 20680 3893
rect 20904 3884 20956 3936
rect 22836 3884 22888 3936
rect 22928 3884 22980 3936
rect 23848 3884 23900 3936
rect 25228 3884 25280 3936
rect 26424 3884 26476 3936
rect 37464 3884 37516 3936
rect 37556 3884 37608 3936
rect 41788 3884 41840 3936
rect 42616 3884 42668 3936
rect 46296 3884 46348 3936
rect 46664 3927 46716 3936
rect 46664 3893 46673 3927
rect 46673 3893 46707 3927
rect 46707 3893 46716 3927
rect 46664 3884 46716 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8024 3680 8076 3732
rect 9312 3612 9364 3664
rect 16488 3612 16540 3664
rect 16764 3612 16816 3664
rect 17960 3680 18012 3732
rect 19248 3680 19300 3732
rect 20812 3723 20864 3732
rect 20812 3689 20821 3723
rect 20821 3689 20855 3723
rect 20855 3689 20864 3723
rect 20812 3680 20864 3689
rect 21456 3680 21508 3732
rect 20076 3612 20128 3664
rect 35532 3680 35584 3732
rect 29092 3612 29144 3664
rect 31392 3612 31444 3664
rect 37372 3680 37424 3732
rect 38568 3680 38620 3732
rect 42432 3680 42484 3732
rect 39304 3612 39356 3664
rect 42340 3612 42392 3664
rect 1860 3544 1912 3596
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 7288 3476 7340 3528
rect 8944 3544 8996 3596
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9220 3544 9272 3553
rect 9404 3544 9456 3596
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 14464 3544 14516 3596
rect 18604 3544 18656 3596
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 11520 3476 11572 3528
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 1308 3408 1360 3460
rect 2044 3340 2096 3392
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 8116 3383 8168 3392
rect 8116 3349 8125 3383
rect 8125 3349 8159 3383
rect 8159 3349 8168 3383
rect 8116 3340 8168 3349
rect 10048 3408 10100 3460
rect 14648 3408 14700 3460
rect 18604 3408 18656 3460
rect 20444 3544 20496 3596
rect 22468 3544 22520 3596
rect 23848 3544 23900 3596
rect 27896 3544 27948 3596
rect 19984 3476 20036 3528
rect 20536 3476 20588 3528
rect 22284 3519 22336 3528
rect 22284 3485 22293 3519
rect 22293 3485 22327 3519
rect 22327 3485 22336 3519
rect 22652 3519 22704 3528
rect 22284 3476 22336 3485
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 22744 3476 22796 3528
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 25504 3519 25556 3528
rect 25504 3485 25513 3519
rect 25513 3485 25547 3519
rect 25547 3485 25556 3519
rect 25504 3476 25556 3485
rect 27620 3519 27672 3528
rect 27620 3485 27629 3519
rect 27629 3485 27663 3519
rect 27663 3485 27672 3519
rect 27620 3476 27672 3485
rect 32864 3544 32916 3596
rect 33876 3544 33928 3596
rect 46296 3587 46348 3596
rect 37924 3476 37976 3528
rect 38568 3476 38620 3528
rect 40408 3519 40460 3528
rect 40408 3485 40417 3519
rect 40417 3485 40451 3519
rect 40451 3485 40460 3519
rect 40408 3476 40460 3485
rect 40868 3519 40920 3528
rect 40868 3485 40877 3519
rect 40877 3485 40911 3519
rect 40911 3485 40920 3519
rect 40868 3476 40920 3485
rect 42432 3476 42484 3528
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 24768 3451 24820 3460
rect 19432 3340 19484 3392
rect 20168 3340 20220 3392
rect 20628 3340 20680 3392
rect 20720 3340 20772 3392
rect 22100 3340 22152 3392
rect 24768 3417 24777 3451
rect 24777 3417 24811 3451
rect 24811 3417 24820 3451
rect 24768 3408 24820 3417
rect 25044 3408 25096 3460
rect 40776 3408 40828 3460
rect 27896 3340 27948 3392
rect 29184 3340 29236 3392
rect 33048 3383 33100 3392
rect 33048 3349 33057 3383
rect 33057 3349 33091 3383
rect 33091 3349 33100 3383
rect 33048 3340 33100 3349
rect 42248 3408 42300 3460
rect 48964 3408 49016 3460
rect 41144 3340 41196 3392
rect 45468 3340 45520 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3792 3136 3844 3188
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 7472 3111 7524 3120
rect 7472 3077 7481 3111
rect 7481 3077 7515 3111
rect 7515 3077 7524 3111
rect 7472 3068 7524 3077
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 664 2932 716 2984
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 14648 3136 14700 3188
rect 14924 3179 14976 3188
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 15660 3136 15712 3188
rect 16672 3136 16724 3188
rect 16948 3136 17000 3188
rect 19248 3136 19300 3188
rect 36728 3179 36780 3188
rect 10048 3111 10100 3120
rect 10048 3077 10057 3111
rect 10057 3077 10091 3111
rect 10091 3077 10100 3111
rect 11704 3111 11756 3120
rect 10048 3068 10100 3077
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 19432 3068 19484 3120
rect 19708 3068 19760 3120
rect 22928 3111 22980 3120
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 16856 3000 16908 3052
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 11888 2932 11940 2984
rect 12256 2975 12308 2984
rect 12256 2941 12265 2975
rect 12265 2941 12299 2975
rect 12299 2941 12308 2975
rect 12256 2932 12308 2941
rect 12394 2932 12446 2984
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 16488 2932 16540 2984
rect 19340 2932 19392 2984
rect 19984 2932 20036 2984
rect 20352 2975 20404 2984
rect 20352 2941 20361 2975
rect 20361 2941 20395 2975
rect 20395 2941 20404 2975
rect 20352 2932 20404 2941
rect 22928 3077 22937 3111
rect 22937 3077 22971 3111
rect 22971 3077 22980 3111
rect 22928 3068 22980 3077
rect 23020 3068 23072 3120
rect 24400 3068 24452 3120
rect 25412 3068 25464 3120
rect 21732 3000 21784 3052
rect 21916 3043 21968 3052
rect 21916 3009 21925 3043
rect 21925 3009 21959 3043
rect 21959 3009 21968 3043
rect 22744 3043 22796 3052
rect 21916 3000 21968 3009
rect 22744 3009 22753 3043
rect 22753 3009 22787 3043
rect 22787 3009 22796 3043
rect 22744 3000 22796 3009
rect 24492 3000 24544 3052
rect 23020 2932 23072 2984
rect 23112 2932 23164 2984
rect 23480 2932 23532 2984
rect 27896 3068 27948 3120
rect 28540 3111 28592 3120
rect 28540 3077 28549 3111
rect 28549 3077 28583 3111
rect 28583 3077 28592 3111
rect 28540 3068 28592 3077
rect 33048 3111 33100 3120
rect 33048 3077 33057 3111
rect 33057 3077 33091 3111
rect 33091 3077 33100 3111
rect 33048 3068 33100 3077
rect 36728 3145 36737 3179
rect 36737 3145 36771 3179
rect 36771 3145 36780 3179
rect 36728 3136 36780 3145
rect 39120 3136 39172 3188
rect 40040 3136 40092 3188
rect 40684 3136 40736 3188
rect 40868 3136 40920 3188
rect 48044 3179 48096 3188
rect 48044 3145 48053 3179
rect 48053 3145 48087 3179
rect 48087 3145 48096 3179
rect 48044 3136 48096 3145
rect 42248 3068 42300 3120
rect 42616 3111 42668 3120
rect 42616 3077 42625 3111
rect 42625 3077 42659 3111
rect 42659 3077 42668 3111
rect 42616 3068 42668 3077
rect 45744 3068 45796 3120
rect 29184 3043 29236 3052
rect 29184 3009 29193 3043
rect 29193 3009 29227 3043
rect 29227 3009 29236 3043
rect 29184 3000 29236 3009
rect 32864 3043 32916 3052
rect 32864 3009 32873 3043
rect 32873 3009 32907 3043
rect 32907 3009 32916 3043
rect 32864 3000 32916 3009
rect 37556 3000 37608 3052
rect 25596 2932 25648 2984
rect 32772 2932 32824 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 37372 2932 37424 2984
rect 39856 2932 39908 2984
rect 40132 3000 40184 3052
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 48320 3000 48372 3052
rect 40592 2975 40644 2984
rect 3884 2864 3936 2916
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 10968 2864 11020 2916
rect 11980 2864 12032 2916
rect 24124 2864 24176 2916
rect 27620 2864 27672 2916
rect 40040 2864 40092 2916
rect 40592 2941 40601 2975
rect 40601 2941 40635 2975
rect 40635 2941 40644 2975
rect 40592 2932 40644 2941
rect 40684 2932 40736 2984
rect 43168 2975 43220 2984
rect 41604 2864 41656 2916
rect 43168 2941 43177 2975
rect 43177 2941 43211 2975
rect 43211 2941 43220 2975
rect 43168 2932 43220 2941
rect 47676 2932 47728 2984
rect 43904 2864 43956 2916
rect 12164 2796 12216 2848
rect 19248 2796 19300 2848
rect 27896 2796 27948 2848
rect 29092 2796 29144 2848
rect 32220 2796 32272 2848
rect 36360 2839 36412 2848
rect 36360 2805 36369 2839
rect 36369 2805 36403 2839
rect 36403 2805 36412 2839
rect 36360 2796 36412 2805
rect 39856 2796 39908 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 12348 2592 12400 2644
rect 15200 2592 15252 2644
rect 2780 2524 2832 2576
rect 6460 2524 6512 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 6828 2456 6880 2508
rect 2596 2320 2648 2372
rect 5172 2388 5224 2440
rect 3240 2320 3292 2372
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 8116 2320 8168 2372
rect 8392 2320 8444 2372
rect 17684 2524 17736 2576
rect 20444 2592 20496 2644
rect 20628 2592 20680 2644
rect 22284 2592 22336 2644
rect 23480 2592 23532 2644
rect 24952 2592 25004 2644
rect 35532 2635 35584 2644
rect 35532 2601 35541 2635
rect 35541 2601 35575 2635
rect 35575 2601 35584 2635
rect 35532 2592 35584 2601
rect 35624 2592 35676 2644
rect 40224 2635 40276 2644
rect 40224 2601 40233 2635
rect 40233 2601 40267 2635
rect 40267 2601 40276 2635
rect 40224 2592 40276 2601
rect 40408 2592 40460 2644
rect 42524 2592 42576 2644
rect 24032 2456 24084 2508
rect 15108 2388 15160 2440
rect 15476 2388 15528 2440
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 20168 2388 20220 2440
rect 23204 2388 23256 2440
rect 16120 2320 16172 2372
rect 20628 2320 20680 2372
rect 21916 2320 21968 2372
rect 25504 2524 25556 2576
rect 27804 2524 27856 2576
rect 32128 2524 32180 2576
rect 24768 2499 24820 2508
rect 24768 2465 24777 2499
rect 24777 2465 24811 2499
rect 24811 2465 24820 2499
rect 24768 2456 24820 2465
rect 25136 2499 25188 2508
rect 25136 2465 25145 2499
rect 25145 2465 25179 2499
rect 25179 2465 25188 2499
rect 25136 2456 25188 2465
rect 27712 2456 27764 2508
rect 32496 2456 32548 2508
rect 40592 2456 40644 2508
rect 41788 2456 41840 2508
rect 26424 2388 26476 2440
rect 28356 2388 28408 2440
rect 29644 2388 29696 2440
rect 35440 2388 35492 2440
rect 38016 2388 38068 2440
rect 39856 2388 39908 2440
rect 41236 2388 41288 2440
rect 43812 2388 43864 2440
rect 44180 2388 44232 2440
rect 46572 2456 46624 2508
rect 47032 2388 47084 2440
rect 48044 2388 48096 2440
rect 26148 2320 26200 2372
rect 27068 2320 27120 2372
rect 36084 2320 36136 2372
rect 39304 2320 39356 2372
rect 40592 2320 40644 2372
rect 46848 2320 46900 2372
rect 38476 2252 38528 2304
rect 45468 2295 45520 2304
rect 45468 2261 45477 2295
rect 45477 2261 45511 2295
rect 45511 2261 45520 2295
rect 45468 2252 45520 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 15568 1980 15620 2032
rect 36360 1980 36412 2032
rect 3976 1912 4028 1964
rect 16028 1912 16080 1964
rect 29276 1912 29328 1964
rect 45468 1912 45520 1964
rect 19340 1504 19392 1556
rect 25596 1504 25648 1556
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4844 49314
rect 4498 49200 4610 49286
rect 32 21418 60 49200
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 46578 1440 47631
rect 1964 47054 1992 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2608 46918 2636 49200
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3790 47016 3846 47025
rect 3790 46951 3846 46960
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1492 46368 1544 46374
rect 1492 46310 1544 46316
rect 2778 46336 2834 46345
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1504 28218 1532 46310
rect 2778 46271 2834 46280
rect 1768 45960 1820 45966
rect 1768 45902 1820 45908
rect 1780 45490 1808 45902
rect 1768 45484 1820 45490
rect 1768 45426 1820 45432
rect 2792 45422 2820 46271
rect 3804 45554 3832 46951
rect 3896 46646 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4816 47054 4844 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7328 49314
rect 7074 49200 7186 49286
rect 5828 47054 5856 49200
rect 7300 47054 7328 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7288 47048 7340 47054
rect 7288 46990 7340 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 6644 46980 6696 46986
rect 6644 46922 6696 46928
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3988 46170 4016 46446
rect 3976 46164 4028 46170
rect 3976 46106 4028 46112
rect 3804 45526 3924 45554
rect 2228 45416 2280 45422
rect 2228 45358 2280 45364
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 2240 45082 2268 45358
rect 2228 45076 2280 45082
rect 2228 45018 2280 45024
rect 3422 44976 3478 44985
rect 3422 44911 3478 44920
rect 2044 44872 2096 44878
rect 2044 44814 2096 44820
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1584 41540 1636 41546
rect 1858 41511 1914 41520
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35465 1624 35634
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1964 34202 1992 40326
rect 1952 34196 2004 34202
rect 1952 34138 2004 34144
rect 1584 33992 1636 33998
rect 1584 33934 1636 33940
rect 1596 32745 1624 33934
rect 1952 33856 2004 33862
rect 1952 33798 2004 33804
rect 1860 33448 1912 33454
rect 1860 33390 1912 33396
rect 1872 32994 1900 33390
rect 1964 33114 1992 33798
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 1872 32966 1992 32994
rect 1964 32910 1992 32966
rect 1952 32904 2004 32910
rect 1952 32846 2004 32852
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1964 31890 1992 32846
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1952 31884 2004 31890
rect 1952 31826 2004 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 2056 31346 2084 44814
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2320 36168 2372 36174
rect 2320 36110 2372 36116
rect 2228 35488 2280 35494
rect 2228 35430 2280 35436
rect 2240 32434 2268 35430
rect 2228 32428 2280 32434
rect 2228 32370 2280 32376
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 1492 28212 1544 28218
rect 1492 28154 1544 28160
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 2148 24954 2176 25094
rect 2136 24948 2188 24954
rect 2136 24890 2188 24896
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 20 21412 72 21418
rect 20 21354 72 21360
rect 2240 21146 2268 31282
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 1964 18970 1992 19246
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2332 18766 2360 36110
rect 2412 32768 2464 32774
rect 2412 32710 2464 32716
rect 2424 32502 2452 32710
rect 2412 32496 2464 32502
rect 2412 32438 2464 32444
rect 3436 19514 3464 44911
rect 3514 43616 3570 43625
rect 3514 43551 3570 43560
rect 3528 35894 3556 43551
rect 3698 39536 3754 39545
rect 3698 39471 3754 39480
rect 3528 35866 3648 35894
rect 3514 31376 3570 31385
rect 3514 31311 3570 31320
rect 3528 30297 3556 31311
rect 3514 30288 3570 30297
rect 3514 30223 3570 30232
rect 3514 28656 3570 28665
rect 3514 28591 3570 28600
rect 3528 27674 3556 28591
rect 3516 27668 3568 27674
rect 3516 27610 3568 27616
rect 3620 21622 3648 35866
rect 3608 21616 3660 21622
rect 3608 21558 3660 21564
rect 3712 21010 3740 39471
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1872 17785 1900 18226
rect 1858 17776 1914 17785
rect 1858 17711 1914 17720
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 2056 4146 2084 16050
rect 3516 15632 3568 15638
rect 3516 15574 3568 15580
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2332 14618 2360 14894
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3402
rect 1596 2514 1624 3878
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3058 1900 3538
rect 2700 3534 2728 14350
rect 3528 7585 3556 15574
rect 3514 7576 3570 7585
rect 3514 7511 3570 7520
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 3126 2084 3334
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 2792 2582 2820 3878
rect 3804 3194 3832 31758
rect 3896 29209 3924 45526
rect 3882 29200 3938 29209
rect 3882 29135 3938 29144
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 3988 19825 4016 20470
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3974 18456 4030 18465
rect 3974 18391 3976 18400
rect 4028 18391 4030 18400
rect 3976 18362 4028 18368
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 3988 17105 4016 17750
rect 3974 17096 4030 17105
rect 3974 17031 4030 17040
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3988 13705 4016 13738
rect 3974 13696 4030 13705
rect 3974 13631 4030 13640
rect 4080 12434 4108 46922
rect 4896 46912 4948 46918
rect 4896 46854 4948 46860
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4632 31890 4660 32302
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4908 18834 4936 46854
rect 5356 46504 5408 46510
rect 5356 46446 5408 46452
rect 5368 46170 5396 46446
rect 5356 46164 5408 46170
rect 5356 46106 5408 46112
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 5460 17338 5488 31826
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3988 12406 4108 12434
rect 3988 6662 4016 12406
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10305 4108 10950
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4066 10296 4122 10305
rect 4214 10288 4522 10308
rect 4066 10231 4122 10240
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 6656 5166 6684 46922
rect 7472 46912 7524 46918
rect 7472 46854 7524 46860
rect 7484 27538 7512 46854
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 7472 27532 7524 27538
rect 7472 27474 7524 27480
rect 8312 25362 8340 45526
rect 9508 36922 9536 46922
rect 10980 46646 11008 49200
rect 10968 46640 11020 46646
rect 10968 46582 11020 46588
rect 11624 46034 11652 49200
rect 12268 47122 12296 49200
rect 12624 47456 12676 47462
rect 12624 47398 12676 47404
rect 12636 47122 12664 47398
rect 12256 47116 12308 47122
rect 12256 47058 12308 47064
rect 12624 47116 12676 47122
rect 12624 47058 12676 47064
rect 12912 46918 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 13740 47122 13860 47138
rect 13740 47116 13872 47122
rect 13740 47110 13820 47116
rect 13820 47058 13872 47064
rect 12900 46912 12952 46918
rect 12900 46854 12952 46860
rect 14200 46594 14228 49200
rect 15488 47546 15516 49200
rect 15488 47518 16344 47546
rect 15844 47456 15896 47462
rect 15844 47398 15896 47404
rect 15016 46980 15068 46986
rect 15016 46922 15068 46928
rect 14200 46566 14320 46594
rect 14292 46510 14320 46566
rect 13084 46504 13136 46510
rect 13084 46446 13136 46452
rect 13820 46504 13872 46510
rect 13820 46446 13872 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 13096 46170 13124 46446
rect 13084 46164 13136 46170
rect 13084 46106 13136 46112
rect 11612 46028 11664 46034
rect 11612 45970 11664 45976
rect 13832 45490 13860 46446
rect 14200 46170 14228 46446
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14096 46096 14148 46102
rect 13924 46044 14096 46050
rect 13924 46038 14148 46044
rect 13924 46022 14136 46038
rect 13924 45966 13952 46022
rect 13912 45960 13964 45966
rect 13912 45902 13964 45908
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 14108 45830 14136 45902
rect 14096 45824 14148 45830
rect 14096 45766 14148 45772
rect 13820 45484 13872 45490
rect 13820 45426 13872 45432
rect 14108 41138 14136 45766
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 9496 36916 9548 36922
rect 9496 36858 9548 36864
rect 14464 33924 14516 33930
rect 14464 33866 14516 33872
rect 14476 33658 14504 33866
rect 14464 33652 14516 33658
rect 14464 33594 14516 33600
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 14476 33114 14504 33458
rect 14464 33108 14516 33114
rect 14464 33050 14516 33056
rect 14464 32904 14516 32910
rect 14464 32846 14516 32852
rect 14476 32230 14504 32846
rect 14740 32496 14792 32502
rect 14740 32438 14792 32444
rect 14464 32224 14516 32230
rect 14464 32166 14516 32172
rect 14476 31346 14504 32166
rect 14464 31340 14516 31346
rect 14464 31282 14516 31288
rect 14752 31278 14780 32438
rect 14740 31272 14792 31278
rect 14740 31214 14792 31220
rect 14924 31204 14976 31210
rect 14924 31146 14976 31152
rect 14936 30258 14964 31146
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 15028 28626 15056 46922
rect 15856 38350 15884 47398
rect 16316 45554 16344 47518
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49200 27150 50000
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49200 31014 50000
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49314 38098 50000
rect 37986 49286 38424 49314
rect 37986 49200 38098 49286
rect 17420 47410 17448 49200
rect 16776 47382 17448 47410
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 16316 45526 16528 45554
rect 15844 38344 15896 38350
rect 15844 38286 15896 38292
rect 16028 36780 16080 36786
rect 16028 36722 16080 36728
rect 15752 36576 15804 36582
rect 15752 36518 15804 36524
rect 15764 36106 15792 36518
rect 15292 36100 15344 36106
rect 15292 36042 15344 36048
rect 15752 36100 15804 36106
rect 15752 36042 15804 36048
rect 15304 35290 15332 36042
rect 16040 35766 16068 36722
rect 16396 36032 16448 36038
rect 16396 35974 16448 35980
rect 16028 35760 16080 35766
rect 16028 35702 16080 35708
rect 15752 35624 15804 35630
rect 15752 35566 15804 35572
rect 15292 35284 15344 35290
rect 15292 35226 15344 35232
rect 15476 34400 15528 34406
rect 15476 34342 15528 34348
rect 15488 33930 15516 34342
rect 15476 33924 15528 33930
rect 15476 33866 15528 33872
rect 15764 33590 15792 35566
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15948 35290 15976 35430
rect 15936 35284 15988 35290
rect 15936 35226 15988 35232
rect 15936 35080 15988 35086
rect 15936 35022 15988 35028
rect 15752 33584 15804 33590
rect 15752 33526 15804 33532
rect 15764 33046 15792 33526
rect 15948 33454 15976 35022
rect 16040 34610 16068 35702
rect 16408 35630 16436 35974
rect 16120 35624 16172 35630
rect 16120 35566 16172 35572
rect 16396 35624 16448 35630
rect 16396 35566 16448 35572
rect 16028 34604 16080 34610
rect 16028 34546 16080 34552
rect 15936 33448 15988 33454
rect 15936 33390 15988 33396
rect 15936 33108 15988 33114
rect 15936 33050 15988 33056
rect 15752 33040 15804 33046
rect 15752 32982 15804 32988
rect 15108 32904 15160 32910
rect 15108 32846 15160 32852
rect 15120 32502 15148 32846
rect 15844 32768 15896 32774
rect 15844 32710 15896 32716
rect 15108 32496 15160 32502
rect 15108 32438 15160 32444
rect 15856 32434 15884 32710
rect 15948 32434 15976 33050
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 16040 31754 16068 34546
rect 16132 32842 16160 35566
rect 16304 33924 16356 33930
rect 16304 33866 16356 33872
rect 16316 33402 16344 33866
rect 16396 33856 16448 33862
rect 16396 33798 16448 33804
rect 16408 33522 16436 33798
rect 16396 33516 16448 33522
rect 16396 33458 16448 33464
rect 16316 33374 16436 33402
rect 16408 33046 16436 33374
rect 16304 33040 16356 33046
rect 16304 32982 16356 32988
rect 16396 33040 16448 33046
rect 16396 32982 16448 32988
rect 16120 32836 16172 32842
rect 16120 32778 16172 32784
rect 16132 31890 16160 32778
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 16224 32026 16252 32302
rect 16316 32026 16344 32982
rect 16396 32836 16448 32842
rect 16396 32778 16448 32784
rect 16212 32020 16264 32026
rect 16212 31962 16264 31968
rect 16304 32020 16356 32026
rect 16304 31962 16356 31968
rect 16408 31958 16436 32778
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 15948 31726 16068 31754
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15304 30394 15332 31078
rect 15844 30660 15896 30666
rect 15844 30602 15896 30608
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 15488 30394 15516 30534
rect 15292 30388 15344 30394
rect 15292 30330 15344 30336
rect 15476 30388 15528 30394
rect 15476 30330 15528 30336
rect 15856 30326 15884 30602
rect 15844 30320 15896 30326
rect 15844 30262 15896 30268
rect 15948 30258 15976 31726
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15936 30252 15988 30258
rect 15936 30194 15988 30200
rect 15212 29510 15240 30194
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15016 28620 15068 28626
rect 15016 28562 15068 28568
rect 15108 27600 15160 27606
rect 15108 27542 15160 27548
rect 15120 27470 15148 27542
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 15384 27396 15436 27402
rect 15384 27338 15436 27344
rect 15396 27130 15424 27338
rect 15384 27124 15436 27130
rect 15384 27066 15436 27072
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 15028 26450 15056 26726
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 12360 25498 12388 25774
rect 12808 25764 12860 25770
rect 12808 25706 12860 25712
rect 12348 25492 12400 25498
rect 12348 25434 12400 25440
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12268 24818 12296 25230
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12544 24818 12572 25094
rect 12820 24886 12848 25706
rect 13740 25294 13768 26318
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11808 24274 11836 24550
rect 12072 24404 12124 24410
rect 11992 24364 12072 24392
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11612 23656 11664 23662
rect 11612 23598 11664 23604
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11532 21690 11560 21966
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11440 21010 11468 21354
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11072 20602 11100 20810
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11440 18290 11468 20402
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11532 20058 11560 20334
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11624 17746 11652 23598
rect 11716 22642 11744 23802
rect 11992 23730 12020 24364
rect 12072 24346 12124 24352
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11716 22114 11744 22578
rect 11992 22574 12020 23666
rect 12084 23322 12112 24074
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 12268 22930 12296 24754
rect 13372 24206 13400 25162
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12360 23730 12388 24006
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 13004 23526 13032 23734
rect 13372 23730 13400 24142
rect 13464 23866 13492 24550
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 12360 23118 12388 23462
rect 13464 23118 13492 23802
rect 13740 23662 13768 25230
rect 13924 24800 13952 25230
rect 14188 25152 14240 25158
rect 14188 25094 14240 25100
rect 14200 24886 14228 25094
rect 14188 24880 14240 24886
rect 14188 24822 14240 24828
rect 14096 24812 14148 24818
rect 13924 24772 14096 24800
rect 13924 23730 13952 24772
rect 14096 24754 14148 24760
rect 14292 24750 14320 25774
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15304 24750 15332 25230
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14832 24744 14884 24750
rect 15292 24744 15344 24750
rect 14832 24686 14884 24692
rect 15028 24704 15292 24732
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 14016 23866 14044 24074
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14108 23866 14136 24006
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14292 23730 14320 24686
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14384 24206 14412 24550
rect 14372 24200 14424 24206
rect 14844 24177 14872 24686
rect 14372 24142 14424 24148
rect 14830 24168 14886 24177
rect 14830 24103 14886 24112
rect 15028 23798 15056 24704
rect 15292 24686 15344 24692
rect 15382 24168 15438 24177
rect 15200 24132 15252 24138
rect 15382 24103 15384 24112
rect 15200 24074 15252 24080
rect 15436 24103 15438 24112
rect 15384 24074 15436 24080
rect 15212 23866 15240 24074
rect 15200 23860 15252 23866
rect 15200 23802 15252 23808
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 14292 23594 14320 23666
rect 14280 23588 14332 23594
rect 14280 23530 14332 23536
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 12268 22902 12388 22930
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 12360 22438 12388 22902
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 11808 22234 11836 22374
rect 11796 22228 11848 22234
rect 11796 22170 11848 22176
rect 11716 22098 11836 22114
rect 11716 22092 11848 22098
rect 11716 22086 11796 22092
rect 11796 22034 11848 22040
rect 11808 22003 11836 22034
rect 12360 21554 12388 22374
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 11808 19854 11836 21490
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11900 20262 11928 20742
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11900 19786 11928 20198
rect 12360 20058 12388 20334
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12544 19854 12572 22510
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 13096 21690 13124 21898
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 13268 20800 13320 20806
rect 13268 20742 13320 20748
rect 13280 20534 13308 20742
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13740 20466 13768 22374
rect 14660 22166 14688 22578
rect 15212 22574 15240 23802
rect 15488 22710 15516 26930
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15672 24070 15700 24754
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15672 23662 15700 24006
rect 15660 23656 15712 23662
rect 15764 23644 15792 24754
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15856 24274 15884 24550
rect 15948 24410 15976 24686
rect 16040 24410 16068 25230
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 16028 23656 16080 23662
rect 15764 23616 16028 23644
rect 15660 23598 15712 23604
rect 16028 23598 16080 23604
rect 16040 23186 16068 23598
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 16040 22778 16068 23122
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 14648 22160 14700 22166
rect 14648 22102 14700 22108
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13832 20942 13860 21490
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 13556 18902 13584 19790
rect 13740 19446 13768 20198
rect 14384 19854 14412 20878
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13832 19174 13860 19654
rect 14200 19446 14228 19654
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 14108 18970 14136 19246
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13556 18630 13584 18838
rect 14200 18766 14228 19110
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17746 11928 18022
rect 12268 17746 12296 18226
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12268 17202 12296 17682
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 13004 16998 13032 18226
rect 13096 18222 13124 18566
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17270 13400 18022
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 11900 16658 11928 16934
rect 13004 16726 13032 16934
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12452 11014 12480 16594
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7668 4146 7696 4558
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 8312 4078 8340 4422
rect 13648 4146 13676 18702
rect 14384 18290 14412 19790
rect 14476 19310 14504 21422
rect 14660 20942 14688 22102
rect 15212 22098 15240 22374
rect 15856 22166 15884 22578
rect 15844 22160 15896 22166
rect 15844 22102 15896 22108
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14476 18970 14504 19246
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15212 18358 15240 18770
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17270 14504 18022
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14200 16590 14228 17070
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4080 3505 4108 3946
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2608 800 2636 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2884 785 2912 2450
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3252 1465 3280 2314
rect 3238 1456 3294 1465
rect 3238 1391 3294 1400
rect 3896 800 3924 2858
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3988 1970 4016 2246
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 5184 800 5212 2382
rect 6472 800 6500 2518
rect 6840 2514 6868 2790
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7116 800 7144 3878
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8036 3534 8064 3674
rect 9232 3602 9260 3878
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 8944 3596 8996 3602
rect 9220 3596 9272 3602
rect 8996 3556 9168 3584
rect 8944 3538 8996 3544
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 9140 3482 9168 3556
rect 9220 3538 9272 3544
rect 9324 3482 9352 3606
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 7300 3058 7328 3470
rect 9140 3454 9352 3482
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7484 3126 7512 3334
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 800 7788 2926
rect 8128 2378 8156 3334
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9416 1714 9444 3538
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10060 3126 10088 3402
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 11532 3058 11560 3470
rect 11716 3126 11744 3878
rect 14292 3602 14320 3878
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 14384 2990 14412 4082
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 11888 2984 11940 2990
rect 12256 2984 12308 2990
rect 11888 2926 11940 2932
rect 11992 2932 12256 2938
rect 11992 2926 12308 2932
rect 12394 2984 12446 2990
rect 12394 2926 12446 2932
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 9048 1686 9444 1714
rect 9048 800 9076 1686
rect 10980 800 11008 2858
rect 11900 2802 11928 2926
rect 11992 2922 12296 2926
rect 11980 2916 12296 2922
rect 12032 2910 12296 2916
rect 11980 2858 12032 2864
rect 12164 2848 12216 2854
rect 11900 2796 12164 2802
rect 11900 2790 12216 2796
rect 11900 2774 12204 2790
rect 12406 2774 12434 2926
rect 14476 2774 14504 3538
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14660 3194 14688 3402
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 12360 2746 12434 2774
rect 14292 2746 14504 2774
rect 14752 2774 14780 14826
rect 15304 13802 15332 22034
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15396 20534 15424 21558
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15764 20942 15792 21286
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15764 20466 15792 20878
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15488 19174 15516 19722
rect 15580 19446 15608 19994
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 18766 15516 19110
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15396 18154 15424 18566
rect 15488 18290 15516 18702
rect 15580 18630 15608 19382
rect 15764 18834 15792 19654
rect 15856 19378 15884 19994
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15580 16998 15608 18566
rect 15672 17746 15700 18566
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14844 3058 14872 3878
rect 14936 3194 14964 4082
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14752 2746 14872 2774
rect 12360 2650 12388 2746
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 14292 1714 14320 2746
rect 14200 1686 14320 1714
rect 14200 800 14228 1686
rect 14844 800 14872 2746
rect 15120 2446 15148 3878
rect 15212 2650 15240 4082
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15488 3058 15516 3878
rect 15672 3194 15700 4558
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 16132 2774 16160 30126
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16408 29306 16436 29514
rect 16396 29300 16448 29306
rect 16396 29242 16448 29248
rect 16500 26450 16528 45526
rect 16580 35692 16632 35698
rect 16580 35634 16632 35640
rect 16592 35018 16620 35634
rect 16672 35488 16724 35494
rect 16672 35430 16724 35436
rect 16684 35154 16712 35430
rect 16672 35148 16724 35154
rect 16672 35090 16724 35096
rect 16580 35012 16632 35018
rect 16580 34954 16632 34960
rect 16592 33998 16620 34954
rect 16580 33992 16632 33998
rect 16580 33934 16632 33940
rect 16672 30048 16724 30054
rect 16672 29990 16724 29996
rect 16684 29170 16712 29990
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16776 25770 16804 47382
rect 18708 47054 18736 49200
rect 18696 47048 18748 47054
rect 18696 46990 18748 46996
rect 19522 47016 19578 47025
rect 19522 46951 19524 46960
rect 19576 46951 19578 46960
rect 19524 46922 19576 46928
rect 19996 46918 20024 49200
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 20168 46504 20220 46510
rect 20168 46446 20220 46452
rect 20180 46170 20208 46446
rect 20168 46164 20220 46170
rect 20168 46106 20220 46112
rect 17316 45892 17368 45898
rect 17316 45834 17368 45840
rect 17328 41414 17356 45834
rect 20076 45824 20128 45830
rect 20076 45766 20128 45772
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 20088 41414 20116 45766
rect 17328 41386 17448 41414
rect 17224 38344 17276 38350
rect 17224 38286 17276 38292
rect 17236 35698 17264 38286
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 17328 36786 17356 37130
rect 17316 36780 17368 36786
rect 17316 36722 17368 36728
rect 17328 36242 17356 36722
rect 17420 36242 17448 41386
rect 19574 41372 19882 41392
rect 20088 41386 20208 41414
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19248 38208 19300 38214
rect 19248 38150 19300 38156
rect 19260 37262 19288 38150
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19524 37800 19576 37806
rect 19524 37742 19576 37748
rect 19800 37800 19852 37806
rect 19800 37742 19852 37748
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 19536 37194 19564 37742
rect 19812 37466 19840 37742
rect 19800 37460 19852 37466
rect 19800 37402 19852 37408
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19524 37188 19576 37194
rect 19524 37130 19576 37136
rect 19984 37188 20036 37194
rect 19984 37130 20036 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 18328 36848 18380 36854
rect 18328 36790 18380 36796
rect 18236 36712 18288 36718
rect 18236 36654 18288 36660
rect 18248 36310 18276 36654
rect 18236 36304 18288 36310
rect 18236 36246 18288 36252
rect 17316 36236 17368 36242
rect 17316 36178 17368 36184
rect 17408 36236 17460 36242
rect 17408 36178 17460 36184
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 17132 35624 17184 35630
rect 17130 35592 17132 35601
rect 17184 35592 17186 35601
rect 16948 35556 17000 35562
rect 17130 35527 17186 35536
rect 16948 35498 17000 35504
rect 16856 34060 16908 34066
rect 16856 34002 16908 34008
rect 16868 31754 16896 34002
rect 16960 33998 16988 35498
rect 17328 34610 17356 36178
rect 18340 35834 18368 36790
rect 19064 36576 19116 36582
rect 19064 36518 19116 36524
rect 19076 36174 19104 36518
rect 19064 36168 19116 36174
rect 19064 36110 19116 36116
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 18972 36100 19024 36106
rect 18972 36042 19024 36048
rect 18328 35828 18380 35834
rect 18328 35770 18380 35776
rect 18984 35698 19012 36042
rect 19260 35766 19288 36110
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 19352 35834 19380 35974
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19248 35760 19300 35766
rect 19248 35702 19300 35708
rect 18328 35692 18380 35698
rect 18328 35634 18380 35640
rect 18972 35692 19024 35698
rect 18972 35634 19024 35640
rect 18340 35086 18368 35634
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18420 34944 18472 34950
rect 18420 34886 18472 34892
rect 18432 34678 18460 34886
rect 18420 34672 18472 34678
rect 18420 34614 18472 34620
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 17328 34134 17356 34546
rect 17684 34536 17736 34542
rect 17684 34478 17736 34484
rect 17696 34202 17724 34478
rect 19064 34400 19116 34406
rect 19064 34342 19116 34348
rect 17684 34196 17736 34202
rect 17684 34138 17736 34144
rect 17316 34128 17368 34134
rect 17316 34070 17368 34076
rect 16948 33992 17000 33998
rect 16948 33934 17000 33940
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 17788 33658 17816 33934
rect 17776 33652 17828 33658
rect 17776 33594 17828 33600
rect 17868 33516 17920 33522
rect 17868 33458 17920 33464
rect 17132 33108 17184 33114
rect 17132 33050 17184 33056
rect 17316 33108 17368 33114
rect 17316 33050 17368 33056
rect 16868 31726 17080 31754
rect 16948 31680 17000 31686
rect 16948 31622 17000 31628
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16868 30394 16896 31282
rect 16960 30734 16988 31622
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 16856 30116 16908 30122
rect 16856 30058 16908 30064
rect 16868 29170 16896 30058
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16764 25764 16816 25770
rect 16764 25706 16816 25712
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16776 24206 16804 24550
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16396 23588 16448 23594
rect 16396 23530 16448 23536
rect 16408 23186 16436 23530
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16224 22030 16252 22714
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16592 21962 16620 23258
rect 16868 22778 16896 25774
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16960 23322 16988 23666
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16684 21350 16712 22578
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16224 16590 16252 20402
rect 16408 19718 16436 20878
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16316 18222 16344 18702
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16684 17882 16712 20742
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16856 19848 16908 19854
rect 16960 19836 16988 20198
rect 16908 19808 16988 19836
rect 16856 19790 16908 19796
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16776 19378 16804 19722
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16868 18902 16896 19110
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16684 17184 16712 17818
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17338 16804 17614
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16960 17270 16988 19808
rect 17052 18086 17080 31726
rect 17144 31686 17172 33050
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17132 31680 17184 31686
rect 17132 31622 17184 31628
rect 17236 31362 17264 32370
rect 17328 31482 17356 33050
rect 17408 32904 17460 32910
rect 17408 32846 17460 32852
rect 17420 32570 17448 32846
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17880 32502 17908 33458
rect 17868 32496 17920 32502
rect 17868 32438 17920 32444
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17604 31822 17632 32166
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17972 31686 18000 33934
rect 18236 33312 18288 33318
rect 18236 33254 18288 33260
rect 18248 32298 18276 33254
rect 18236 32292 18288 32298
rect 18236 32234 18288 32240
rect 18340 32230 18368 33934
rect 19076 33930 19104 34342
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 19076 33522 19104 33866
rect 19260 33522 19288 35702
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19996 34066 20024 37130
rect 20088 36922 20116 37198
rect 20076 36916 20128 36922
rect 20076 36858 20128 36864
rect 20076 36236 20128 36242
rect 20076 36178 20128 36184
rect 19984 34060 20036 34066
rect 19984 34002 20036 34008
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19996 33658 20024 34002
rect 20088 33862 20116 36178
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 19064 33516 19116 33522
rect 19064 33458 19116 33464
rect 19248 33516 19300 33522
rect 19248 33458 19300 33464
rect 19076 32842 19104 33458
rect 19260 32910 19288 33458
rect 19984 33448 20036 33454
rect 19984 33390 20036 33396
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19064 32836 19116 32842
rect 19064 32778 19116 32784
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 18328 32224 18380 32230
rect 18328 32166 18380 32172
rect 18340 31822 18368 32166
rect 19248 32020 19300 32026
rect 19248 31962 19300 31968
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 17960 31680 18012 31686
rect 18144 31680 18196 31686
rect 18012 31628 18092 31634
rect 17960 31622 18092 31628
rect 18144 31622 18196 31628
rect 18328 31680 18380 31686
rect 18328 31622 18380 31628
rect 17972 31606 18092 31622
rect 17972 31557 18000 31606
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17132 31340 17184 31346
rect 17236 31334 17356 31362
rect 17132 31282 17184 31288
rect 17144 30938 17172 31282
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 17132 30932 17184 30938
rect 17132 30874 17184 30880
rect 17236 30870 17264 31214
rect 17224 30864 17276 30870
rect 17224 30806 17276 30812
rect 17132 29708 17184 29714
rect 17132 29650 17184 29656
rect 17144 29594 17172 29650
rect 17236 29594 17264 30806
rect 17328 30734 17356 31334
rect 18064 31278 18092 31606
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17880 30938 17908 31078
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17420 30258 17448 30534
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17788 29850 17816 30602
rect 17880 30258 17908 30874
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17776 29844 17828 29850
rect 17776 29786 17828 29792
rect 17144 29566 17264 29594
rect 17132 29504 17184 29510
rect 17132 29446 17184 29452
rect 17144 29034 17172 29446
rect 17236 29034 17264 29566
rect 17788 29238 17816 29786
rect 17776 29232 17828 29238
rect 17776 29174 17828 29180
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17132 29028 17184 29034
rect 17132 28970 17184 28976
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17236 26926 17264 28970
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17236 26450 17264 26862
rect 17224 26444 17276 26450
rect 17224 26386 17276 26392
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 17420 24818 17448 25162
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17144 24070 17172 24754
rect 17328 24410 17356 24754
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17144 23730 17172 24006
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17144 23050 17172 23462
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17328 22234 17356 22510
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17420 20466 17448 24142
rect 17512 22094 17540 29106
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17604 28082 17632 28358
rect 17788 28082 17816 28358
rect 17972 28082 18000 28494
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17868 27600 17920 27606
rect 17868 27542 17920 27548
rect 17880 24274 17908 27542
rect 17972 26790 18000 28018
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 18156 25378 18184 31622
rect 18340 31414 18368 31622
rect 18328 31408 18380 31414
rect 18328 31350 18380 31356
rect 19260 30734 19288 31962
rect 19340 31884 19392 31890
rect 19340 31826 19392 31832
rect 19352 31482 19380 31826
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19340 31340 19392 31346
rect 19340 31282 19392 31288
rect 19352 30938 19380 31282
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 19248 30728 19300 30734
rect 19248 30670 19300 30676
rect 18236 30116 18288 30122
rect 18236 30058 18288 30064
rect 18248 28626 18276 30058
rect 19260 29646 19288 30670
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19352 30122 19380 30330
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 18248 28082 18276 28562
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 18236 27872 18288 27878
rect 18236 27814 18288 27820
rect 18248 26926 18276 27814
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18616 26586 18644 26930
rect 18604 26580 18656 26586
rect 18604 26522 18656 26528
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19260 25906 19288 26250
rect 19352 25906 19380 30058
rect 19248 25900 19300 25906
rect 19248 25842 19300 25848
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19260 25430 19288 25842
rect 19444 25498 19472 30194
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19800 29096 19852 29102
rect 19800 29038 19852 29044
rect 19812 28762 19840 29038
rect 19800 28756 19852 28762
rect 19800 28698 19852 28704
rect 19996 28422 20024 33390
rect 20088 33318 20116 33798
rect 20076 33312 20128 33318
rect 20076 33254 20128 33260
rect 20076 32496 20128 32502
rect 20076 32438 20128 32444
rect 20088 31890 20116 32438
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 20076 30660 20128 30666
rect 20076 30602 20128 30608
rect 20088 29510 20116 30602
rect 20076 29504 20128 29510
rect 20076 29446 20128 29452
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19996 28014 20024 28358
rect 20088 28082 20116 28426
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19996 27010 20024 27406
rect 20180 27146 20208 41386
rect 20364 38350 20392 46990
rect 20640 46510 20668 49200
rect 21180 47116 21232 47122
rect 21180 47058 21232 47064
rect 20904 47048 20956 47054
rect 20904 46990 20956 46996
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20720 46164 20772 46170
rect 20720 46106 20772 46112
rect 20732 45490 20760 46106
rect 20916 46034 20944 46990
rect 20904 46028 20956 46034
rect 20904 45970 20956 45976
rect 20904 45892 20956 45898
rect 20904 45834 20956 45840
rect 20916 45626 20944 45834
rect 20904 45620 20956 45626
rect 20904 45562 20956 45568
rect 20720 45484 20772 45490
rect 20720 45426 20772 45432
rect 20732 41414 20760 45426
rect 20732 41386 20944 41414
rect 20536 38752 20588 38758
rect 20536 38694 20588 38700
rect 20352 38344 20404 38350
rect 20352 38286 20404 38292
rect 20260 37324 20312 37330
rect 20260 37266 20312 37272
rect 20272 35766 20300 37266
rect 20444 36780 20496 36786
rect 20444 36722 20496 36728
rect 20260 35760 20312 35766
rect 20260 35702 20312 35708
rect 20272 35562 20300 35702
rect 20260 35556 20312 35562
rect 20260 35498 20312 35504
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20364 31414 20392 33458
rect 20352 31408 20404 31414
rect 20352 31350 20404 31356
rect 20260 29504 20312 29510
rect 20260 29446 20312 29452
rect 20272 29238 20300 29446
rect 20260 29232 20312 29238
rect 20260 29174 20312 29180
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20364 28218 20392 28494
rect 20456 28234 20484 36722
rect 20548 31346 20576 38694
rect 20628 38344 20680 38350
rect 20628 38286 20680 38292
rect 20640 37262 20668 38286
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 20640 36786 20668 37198
rect 20628 36780 20680 36786
rect 20628 36722 20680 36728
rect 20812 35284 20864 35290
rect 20812 35226 20864 35232
rect 20824 34610 20852 35226
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20732 34066 20760 34342
rect 20720 34060 20772 34066
rect 20720 34002 20772 34008
rect 20628 33652 20680 33658
rect 20628 33594 20680 33600
rect 20640 32502 20668 33594
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20732 30870 20760 31282
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20824 30938 20852 31214
rect 20812 30932 20864 30938
rect 20812 30874 20864 30880
rect 20720 30864 20772 30870
rect 20720 30806 20772 30812
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 20720 30048 20772 30054
rect 20720 29990 20772 29996
rect 20536 28552 20588 28558
rect 20732 28506 20760 29990
rect 20824 29850 20852 30194
rect 20812 29844 20864 29850
rect 20812 29786 20864 29792
rect 20588 28500 20760 28506
rect 20536 28494 20760 28500
rect 20548 28478 20760 28494
rect 20352 28212 20404 28218
rect 20456 28206 20576 28234
rect 20352 28154 20404 28160
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20180 27118 20300 27146
rect 19996 26982 20208 27010
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19996 26042 20024 26250
rect 19984 26036 20036 26042
rect 19984 25978 20036 25984
rect 20088 25702 20116 26862
rect 20180 26042 20208 26982
rect 20168 26036 20220 26042
rect 20168 25978 20220 25984
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 18064 25350 18184 25378
rect 19248 25424 19300 25430
rect 19248 25366 19300 25372
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 18064 23594 18092 25350
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18156 24818 18184 25230
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19352 24682 19380 24754
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18340 24206 18368 24550
rect 19352 24342 19380 24618
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18052 23588 18104 23594
rect 18052 23530 18104 23536
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17880 22778 17908 23258
rect 18340 23118 18368 24006
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19536 23186 19564 23462
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 18340 22710 18368 22918
rect 19352 22778 19380 23054
rect 19628 23050 19656 23666
rect 19904 23118 19932 23666
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19616 23044 19668 23050
rect 19616 22986 19668 22992
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22778 19472 22918
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 17684 22704 17736 22710
rect 18328 22704 18380 22710
rect 17736 22652 18000 22658
rect 17684 22646 18000 22652
rect 18328 22646 18380 22652
rect 19352 22658 19380 22714
rect 17696 22630 18000 22646
rect 19352 22630 19472 22658
rect 17512 22066 17632 22094
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17512 20466 17540 20742
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17236 19922 17264 20198
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 17236 19446 17264 19722
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 17144 17882 17172 18158
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 16764 17196 16816 17202
rect 16684 17156 16764 17184
rect 16684 16658 16712 17156
rect 16764 17138 16816 17144
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16224 16114 16252 16526
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16316 15570 16344 16390
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 17604 12434 17632 22066
rect 17972 21350 18000 22630
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18616 22166 18644 22510
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 19352 22098 19380 22374
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19444 22030 19472 22630
rect 19996 22438 20024 23666
rect 20088 22778 20116 24142
rect 20168 23044 20220 23050
rect 20168 22986 20220 22992
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 20180 22574 20208 22986
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 20272 22094 20300 27118
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20364 22438 20392 24074
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20272 22066 20392 22094
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17972 20942 18000 21286
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17972 18766 18000 20878
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19378 18092 19654
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 18358 17724 18566
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17880 17338 17908 17614
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17696 16658 17724 17138
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17604 12406 17724 12434
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16500 2990 16528 3606
rect 16592 3534 16620 3878
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16684 3194 16712 4558
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16776 3670 16804 4082
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16868 3058 16896 4490
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 16960 3194 16988 4150
rect 17144 4010 17172 4150
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17236 3534 17264 3878
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17328 3058 17356 4422
rect 17406 3496 17462 3505
rect 17406 3431 17462 3440
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16040 2746 16160 2774
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15488 800 15516 2382
rect 15580 2038 15608 2382
rect 15568 2032 15620 2038
rect 15568 1974 15620 1980
rect 16040 1970 16068 2746
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 16132 800 16160 2314
rect 17420 800 17448 3431
rect 17696 2582 17724 12406
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17880 3534 17908 3878
rect 17972 3738 18000 4082
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 18432 2394 18460 20198
rect 18524 19990 18552 21490
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18616 19378 18644 19858
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18708 19718 18736 19790
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18800 19446 18828 19654
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18892 17746 18920 21490
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18984 20534 19012 21286
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 19168 19922 19196 20538
rect 19444 20398 19472 21966
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 20364 20942 20392 22066
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18984 19242 19012 19722
rect 19076 19378 19104 19790
rect 19352 19786 19380 20266
rect 20364 19922 20392 20742
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19800 19440 19852 19446
rect 19798 19408 19800 19417
rect 19852 19408 19854 19417
rect 19064 19372 19116 19378
rect 19798 19343 19854 19352
rect 19892 19372 19944 19378
rect 19064 19314 19116 19320
rect 19996 19360 20024 19790
rect 20260 19712 20312 19718
rect 20166 19680 20222 19689
rect 20260 19654 20312 19660
rect 20350 19680 20406 19689
rect 20166 19615 20222 19624
rect 20180 19446 20208 19615
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 19944 19332 20024 19360
rect 19892 19314 19944 19320
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 19904 18902 19932 19314
rect 20272 19174 20300 19654
rect 20350 19615 20406 19624
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18524 16794 18552 17070
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18524 6866 18552 15982
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 19168 4214 19196 18158
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19352 15706 19380 17070
rect 19444 16794 19472 17546
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19996 16250 20024 17070
rect 20088 16658 20116 17274
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 20088 15570 20116 16390
rect 20180 16182 20208 17546
rect 20364 17270 20392 19615
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20364 17134 20392 17206
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20260 16720 20312 16726
rect 20260 16662 20312 16668
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20272 15502 20300 16662
rect 20364 16658 20392 17070
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20456 12434 20484 28018
rect 20548 25294 20576 28206
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 26586 20668 27270
rect 20824 26994 20852 27338
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 20824 26586 20852 26930
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20548 23798 20576 24210
rect 20812 24064 20864 24070
rect 20812 24006 20864 24012
rect 20824 23866 20852 24006
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20536 23792 20588 23798
rect 20536 23734 20588 23740
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 22710 20576 22918
rect 20536 22704 20588 22710
rect 20536 22646 20588 22652
rect 20640 22642 20668 23666
rect 20732 22642 20760 23666
rect 20824 23118 20852 23802
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20824 22710 20852 22918
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20640 22094 20668 22578
rect 20548 22066 20668 22094
rect 20548 20058 20576 22066
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20626 19680 20682 19689
rect 20626 19615 20682 19624
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20548 19417 20576 19450
rect 20640 19446 20668 19615
rect 20732 19553 20760 22578
rect 20916 21418 20944 41386
rect 21088 38480 21140 38486
rect 21088 38422 21140 38428
rect 20996 33924 21048 33930
rect 20996 33866 21048 33872
rect 21008 33114 21036 33866
rect 20996 33108 21048 33114
rect 20996 33050 21048 33056
rect 21100 32910 21128 38422
rect 21192 34542 21220 47058
rect 21284 46034 21312 49200
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 21824 46912 21876 46918
rect 21824 46854 21876 46860
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 21836 39030 21864 46854
rect 24872 46646 24900 46990
rect 24860 46640 24912 46646
rect 24860 46582 24912 46588
rect 25148 46510 25176 49200
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25504 45892 25556 45898
rect 25504 45834 25556 45840
rect 25516 45626 25544 45834
rect 25792 45830 25820 49200
rect 27080 46889 27108 49200
rect 28368 47054 28396 49200
rect 29092 47184 29144 47190
rect 29092 47126 29144 47132
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 28816 46980 28868 46986
rect 28816 46922 28868 46928
rect 27066 46880 27122 46889
rect 27066 46815 27122 46824
rect 26240 46028 26292 46034
rect 26240 45970 26292 45976
rect 25780 45824 25832 45830
rect 25780 45766 25832 45772
rect 24768 45620 24820 45626
rect 24768 45562 24820 45568
rect 25504 45620 25556 45626
rect 25504 45562 25556 45568
rect 23572 39500 23624 39506
rect 23572 39442 23624 39448
rect 22744 39296 22796 39302
rect 22744 39238 22796 39244
rect 22756 39030 22784 39238
rect 23584 39098 23612 39442
rect 24780 39438 24808 45562
rect 26252 45422 26280 45970
rect 26240 45416 26292 45422
rect 26240 45358 26292 45364
rect 25780 43784 25832 43790
rect 25780 43726 25832 43732
rect 24768 39432 24820 39438
rect 24768 39374 24820 39380
rect 24492 39296 24544 39302
rect 24492 39238 24544 39244
rect 23572 39092 23624 39098
rect 23572 39034 23624 39040
rect 21824 39024 21876 39030
rect 21824 38966 21876 38972
rect 22744 39024 22796 39030
rect 22744 38966 22796 38972
rect 23480 39024 23532 39030
rect 23480 38966 23532 38972
rect 21916 38888 21968 38894
rect 21916 38830 21968 38836
rect 21824 37868 21876 37874
rect 21824 37810 21876 37816
rect 21836 37466 21864 37810
rect 21824 37460 21876 37466
rect 21824 37402 21876 37408
rect 21928 37262 21956 38830
rect 23492 38554 23520 38966
rect 23480 38548 23532 38554
rect 23480 38490 23532 38496
rect 23584 38434 23612 39034
rect 24216 38752 24268 38758
rect 24216 38694 24268 38700
rect 23492 38406 23612 38434
rect 23664 38412 23716 38418
rect 22100 37732 22152 37738
rect 22100 37674 22152 37680
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 21836 35698 21864 36722
rect 22112 36718 22140 37674
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 22100 36712 22152 36718
rect 22100 36654 22152 36660
rect 22204 36310 22232 37130
rect 23204 36644 23256 36650
rect 23204 36586 23256 36592
rect 22192 36304 22244 36310
rect 22192 36246 22244 36252
rect 22928 36236 22980 36242
rect 22928 36178 22980 36184
rect 23020 36236 23072 36242
rect 23020 36178 23072 36184
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 21916 35760 21968 35766
rect 21916 35702 21968 35708
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 21180 34536 21232 34542
rect 21180 34478 21232 34484
rect 21284 34134 21312 34614
rect 21468 34610 21496 35090
rect 21732 35080 21784 35086
rect 21732 35022 21784 35028
rect 21456 34604 21508 34610
rect 21456 34546 21508 34552
rect 21744 34474 21772 35022
rect 21928 34678 21956 35702
rect 22572 35442 22600 36110
rect 22650 35728 22706 35737
rect 22650 35663 22652 35672
rect 22704 35663 22706 35672
rect 22652 35634 22704 35640
rect 22572 35414 22692 35442
rect 22664 35290 22692 35414
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 22652 35284 22704 35290
rect 22652 35226 22704 35232
rect 22100 35012 22152 35018
rect 22100 34954 22152 34960
rect 22112 34746 22140 34954
rect 22284 34944 22336 34950
rect 22284 34886 22336 34892
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 21916 34672 21968 34678
rect 21916 34614 21968 34620
rect 21732 34468 21784 34474
rect 21732 34410 21784 34416
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 21744 34202 21772 34410
rect 21824 34400 21876 34406
rect 21824 34342 21876 34348
rect 21732 34196 21784 34202
rect 21732 34138 21784 34144
rect 21272 34128 21324 34134
rect 21272 34070 21324 34076
rect 21836 34066 21864 34342
rect 21824 34060 21876 34066
rect 21824 34002 21876 34008
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 22020 33522 22048 33934
rect 22112 33930 22140 34410
rect 22192 34400 22244 34406
rect 22192 34342 22244 34348
rect 22100 33924 22152 33930
rect 22100 33866 22152 33872
rect 21640 33516 21692 33522
rect 21640 33458 21692 33464
rect 22008 33516 22060 33522
rect 22008 33458 22060 33464
rect 21548 33312 21600 33318
rect 21548 33254 21600 33260
rect 21088 32904 21140 32910
rect 21140 32852 21220 32858
rect 21088 32846 21220 32852
rect 21100 32830 21220 32846
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 21100 31482 21128 31826
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 21192 31210 21220 32830
rect 21560 31278 21588 33254
rect 21652 33114 21680 33458
rect 21640 33108 21692 33114
rect 21640 33050 21692 33056
rect 21652 31414 21680 33050
rect 22020 31754 22048 33458
rect 22112 32774 22140 33866
rect 22204 33590 22232 34342
rect 22296 34202 22324 34886
rect 22284 34196 22336 34202
rect 22284 34138 22336 34144
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22192 33584 22244 33590
rect 22192 33526 22244 33532
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 21744 31726 22048 31754
rect 21640 31408 21692 31414
rect 21640 31350 21692 31356
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21180 31204 21232 31210
rect 21180 31146 21232 31152
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 21008 30258 21036 30738
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 21008 29850 21036 30194
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 21192 29714 21220 31146
rect 21640 30116 21692 30122
rect 21640 30058 21692 30064
rect 21652 29782 21680 30058
rect 21640 29776 21692 29782
rect 21640 29718 21692 29724
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 21272 29640 21324 29646
rect 21744 29594 21772 31726
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 31362 22048 31622
rect 21836 31346 22048 31362
rect 21824 31340 22048 31346
rect 21876 31334 22048 31340
rect 21824 31282 21876 31288
rect 22020 30734 22048 31334
rect 22100 31204 22152 31210
rect 22100 31146 22152 31152
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 21272 29582 21324 29588
rect 21284 29306 21312 29582
rect 21560 29572 21772 29594
rect 21824 29640 21876 29646
rect 21824 29582 21876 29588
rect 21560 29566 21640 29572
rect 21272 29300 21324 29306
rect 21272 29242 21324 29248
rect 21560 29170 21588 29566
rect 21692 29566 21772 29572
rect 21640 29514 21692 29520
rect 21652 29483 21680 29514
rect 21732 29504 21784 29510
rect 21732 29446 21784 29452
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 21548 29164 21600 29170
rect 21548 29106 21600 29112
rect 21272 28688 21324 28694
rect 21272 28630 21324 28636
rect 21284 27470 21312 28630
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21100 26926 21128 27406
rect 21180 27328 21232 27334
rect 21180 27270 21232 27276
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 21192 26518 21220 27270
rect 21284 26790 21312 27406
rect 21560 26994 21588 29106
rect 21652 28422 21680 29174
rect 21744 28762 21772 29446
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21836 28626 21864 29582
rect 21928 29306 21956 29786
rect 22020 29646 22048 30670
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 21916 29300 21968 29306
rect 21916 29242 21968 29248
rect 21824 28620 21876 28626
rect 21824 28562 21876 28568
rect 21836 28506 21864 28562
rect 21836 28478 21956 28506
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21652 28082 21680 28358
rect 21928 28082 21956 28478
rect 21640 28076 21692 28082
rect 21640 28018 21692 28024
rect 21916 28076 21968 28082
rect 21916 28018 21968 28024
rect 22020 27962 22048 29582
rect 21836 27934 22048 27962
rect 21836 27878 21864 27934
rect 21824 27872 21876 27878
rect 21824 27814 21876 27820
rect 21916 27872 21968 27878
rect 21916 27814 21968 27820
rect 21928 27062 21956 27814
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 21916 27056 21968 27062
rect 21916 26998 21968 27004
rect 21548 26988 21600 26994
rect 21548 26930 21600 26936
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 21640 26920 21692 26926
rect 21640 26862 21692 26868
rect 21548 26852 21600 26858
rect 21548 26794 21600 26800
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21180 26512 21232 26518
rect 21180 26454 21232 26460
rect 21192 25906 21220 26454
rect 21560 26314 21588 26794
rect 21652 26450 21680 26862
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21548 26308 21600 26314
rect 21548 26250 21600 26256
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21560 25498 21588 26250
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21652 25362 21680 26386
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21744 25294 21772 26930
rect 21928 26586 21956 26998
rect 22020 26790 22048 27066
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 21928 25498 21956 26522
rect 22112 26246 22140 31146
rect 22204 26382 22232 33526
rect 22480 33386 22508 33934
rect 22468 33380 22520 33386
rect 22468 33322 22520 33328
rect 22376 32768 22428 32774
rect 22376 32710 22428 32716
rect 22388 32502 22416 32710
rect 22376 32496 22428 32502
rect 22376 32438 22428 32444
rect 22468 31816 22520 31822
rect 22468 31758 22520 31764
rect 22480 31482 22508 31758
rect 22572 31754 22600 35226
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22756 33046 22784 35090
rect 22836 35080 22888 35086
rect 22836 35022 22888 35028
rect 22848 34542 22876 35022
rect 22836 34536 22888 34542
rect 22836 34478 22888 34484
rect 22744 33040 22796 33046
rect 22744 32982 22796 32988
rect 22652 32496 22704 32502
rect 22652 32438 22704 32444
rect 22664 32026 22692 32438
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22572 31726 22692 31754
rect 22468 31476 22520 31482
rect 22468 31418 22520 31424
rect 22560 31340 22612 31346
rect 22560 31282 22612 31288
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22296 30258 22324 30670
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 22296 26518 22324 30194
rect 22572 29646 22600 31282
rect 22664 29850 22692 31726
rect 22652 29844 22704 29850
rect 22652 29786 22704 29792
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22652 29708 22704 29714
rect 22652 29650 22704 29656
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22664 29170 22692 29650
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 22664 28558 22692 28698
rect 22848 28558 22876 29786
rect 22940 29306 22968 36178
rect 23032 36038 23060 36178
rect 23020 36032 23072 36038
rect 23020 35974 23072 35980
rect 23032 35494 23060 35974
rect 23216 35834 23244 36586
rect 23204 35828 23256 35834
rect 23204 35770 23256 35776
rect 23112 35556 23164 35562
rect 23112 35498 23164 35504
rect 23020 35488 23072 35494
rect 23020 35430 23072 35436
rect 23124 35018 23152 35498
rect 23216 35494 23244 35770
rect 23204 35488 23256 35494
rect 23204 35430 23256 35436
rect 23112 35012 23164 35018
rect 23112 34954 23164 34960
rect 23296 35012 23348 35018
rect 23296 34954 23348 34960
rect 23112 33380 23164 33386
rect 23112 33322 23164 33328
rect 23124 30938 23152 33322
rect 23204 33040 23256 33046
rect 23204 32982 23256 32988
rect 23216 32774 23244 32982
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 23112 30932 23164 30938
rect 23112 30874 23164 30880
rect 23124 29510 23152 30874
rect 23020 29504 23072 29510
rect 23020 29446 23072 29452
rect 23112 29504 23164 29510
rect 23112 29446 23164 29452
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 23032 29238 23060 29446
rect 23020 29232 23072 29238
rect 23020 29174 23072 29180
rect 22928 29096 22980 29102
rect 22928 29038 22980 29044
rect 22940 28762 22968 29038
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 23216 28558 23244 32710
rect 23308 30666 23336 34954
rect 23400 34678 23428 37606
rect 23492 36938 23520 38406
rect 23664 38354 23716 38360
rect 23572 38344 23624 38350
rect 23572 38286 23624 38292
rect 23584 37874 23612 38286
rect 23572 37868 23624 37874
rect 23572 37810 23624 37816
rect 23572 37120 23624 37126
rect 23676 37074 23704 38354
rect 24228 38350 24256 38694
rect 24504 38486 24532 39238
rect 24492 38480 24544 38486
rect 24492 38422 24544 38428
rect 24216 38344 24268 38350
rect 24216 38286 24268 38292
rect 23848 37936 23900 37942
rect 23848 37878 23900 37884
rect 23756 37800 23808 37806
rect 23756 37742 23808 37748
rect 23624 37068 23704 37074
rect 23572 37062 23704 37068
rect 23584 37046 23704 37062
rect 23492 36910 23612 36938
rect 23676 36922 23704 37046
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23492 36310 23520 36722
rect 23480 36304 23532 36310
rect 23480 36246 23532 36252
rect 23480 36100 23532 36106
rect 23480 36042 23532 36048
rect 23492 35290 23520 36042
rect 23584 35714 23612 36910
rect 23664 36916 23716 36922
rect 23664 36858 23716 36864
rect 23768 35834 23796 37742
rect 23860 37126 23888 37878
rect 24952 37800 25004 37806
rect 24952 37742 25004 37748
rect 24964 37466 24992 37742
rect 24952 37460 25004 37466
rect 24952 37402 25004 37408
rect 25136 37256 25188 37262
rect 25136 37198 25188 37204
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 23860 36174 23888 37062
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 24032 36032 24084 36038
rect 24032 35974 24084 35980
rect 23756 35828 23808 35834
rect 23756 35770 23808 35776
rect 23584 35686 23704 35714
rect 23768 35698 23796 35770
rect 23572 35624 23624 35630
rect 23572 35566 23624 35572
rect 23480 35284 23532 35290
rect 23480 35226 23532 35232
rect 23584 34678 23612 35566
rect 23388 34672 23440 34678
rect 23388 34614 23440 34620
rect 23572 34672 23624 34678
rect 23572 34614 23624 34620
rect 23584 34202 23612 34614
rect 23572 34196 23624 34202
rect 23572 34138 23624 34144
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23400 31822 23428 32506
rect 23676 32366 23704 35686
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 24044 35630 24072 35974
rect 24584 35760 24636 35766
rect 24584 35702 24636 35708
rect 24032 35624 24084 35630
rect 24032 35566 24084 35572
rect 24124 35624 24176 35630
rect 24124 35566 24176 35572
rect 24044 35154 24072 35566
rect 24136 35222 24164 35566
rect 24124 35216 24176 35222
rect 24124 35158 24176 35164
rect 24032 35148 24084 35154
rect 24032 35090 24084 35096
rect 23940 35080 23992 35086
rect 23940 35022 23992 35028
rect 24492 35080 24544 35086
rect 24492 35022 24544 35028
rect 23664 32360 23716 32366
rect 23664 32302 23716 32308
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23492 31754 23520 31826
rect 23952 31754 23980 35022
rect 24504 34785 24532 35022
rect 24490 34776 24546 34785
rect 24490 34711 24546 34720
rect 24492 34196 24544 34202
rect 24492 34138 24544 34144
rect 24400 32904 24452 32910
rect 24400 32846 24452 32852
rect 24308 32428 24360 32434
rect 24308 32370 24360 32376
rect 23492 31726 23796 31754
rect 23952 31726 24072 31754
rect 23768 31482 23796 31726
rect 23756 31476 23808 31482
rect 23756 31418 23808 31424
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23584 30802 23612 31078
rect 23572 30796 23624 30802
rect 23572 30738 23624 30744
rect 23296 30660 23348 30666
rect 23296 30602 23348 30608
rect 23756 30320 23808 30326
rect 23756 30262 23808 30268
rect 23768 30122 23796 30262
rect 23756 30116 23808 30122
rect 23756 30058 23808 30064
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 23308 28626 23336 29038
rect 23296 28620 23348 28626
rect 23296 28562 23348 28568
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 22848 27606 22876 28494
rect 22836 27600 22888 27606
rect 22836 27542 22888 27548
rect 22284 26512 22336 26518
rect 22284 26454 22336 26460
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22112 25906 22140 26182
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 21916 25492 21968 25498
rect 21916 25434 21968 25440
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 21008 24206 21036 24686
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 21008 23118 21036 24142
rect 21376 23866 21404 25230
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21468 23662 21496 24142
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21836 23730 21864 24006
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 21468 23118 21496 23598
rect 22112 23322 22140 23598
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 22204 23118 22232 24278
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21836 22642 21864 22918
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22204 22098 22232 22374
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 22204 21690 22232 22034
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 20718 19544 20774 19553
rect 20718 19479 20774 19488
rect 20628 19440 20680 19446
rect 20534 19408 20590 19417
rect 20628 19382 20680 19388
rect 20534 19343 20590 19352
rect 20812 19372 20864 19378
rect 21088 19372 21140 19378
rect 20864 19332 20944 19360
rect 20812 19314 20864 19320
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20732 17134 20760 18770
rect 20916 18766 20944 19332
rect 21088 19314 21140 19320
rect 20996 19236 21048 19242
rect 20996 19178 21048 19184
rect 21008 18902 21036 19178
rect 21100 18970 21128 19314
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 16590 20760 17070
rect 20916 16998 20944 18702
rect 21008 17542 21036 18838
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20732 15502 20760 16526
rect 20916 16454 20944 16934
rect 21008 16522 21036 17478
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 21192 16114 21220 17614
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 21192 15366 21220 16050
rect 21284 15910 21312 20810
rect 22204 20618 22232 21626
rect 22296 21554 22324 26454
rect 22376 25152 22428 25158
rect 22376 25094 22428 25100
rect 22388 23118 22416 25094
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22112 20590 22232 20618
rect 22006 19544 22062 19553
rect 22006 19479 22062 19488
rect 22020 19446 22048 19479
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21560 18358 21588 18770
rect 21916 18760 21968 18766
rect 22020 18748 22048 19382
rect 22112 18902 22140 20590
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 20058 22232 20402
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22204 19378 22232 19654
rect 22296 19446 22324 21490
rect 22480 20398 22508 24346
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22572 20398 22600 20878
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22572 19786 22600 20334
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 22100 18760 22152 18766
rect 22020 18720 22100 18748
rect 21916 18702 21968 18708
rect 22100 18702 22152 18708
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21928 18204 21956 18702
rect 22100 18216 22152 18222
rect 21928 18176 22100 18204
rect 22100 18158 22152 18164
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22112 17882 22140 18022
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22388 17746 22416 19654
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22388 17202 22416 17682
rect 22664 17678 22692 20538
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22756 17882 22784 18294
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22652 17672 22704 17678
rect 22704 17620 22784 17626
rect 22652 17614 22784 17620
rect 22664 17598 22784 17614
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 16658 21404 16934
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 22756 16250 22784 17598
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22192 16176 22244 16182
rect 22192 16118 22244 16124
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 22112 15706 22140 15982
rect 22204 15910 22232 16118
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22756 15502 22784 16186
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20364 12406 20484 12434
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19156 4208 19208 4214
rect 19156 4150 19208 4156
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18524 3534 18552 3878
rect 18616 3602 18644 4082
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18694 3768 18750 3777
rect 18694 3703 18750 3712
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18512 3528 18564 3534
rect 18708 3482 18736 3703
rect 18512 3470 18564 3476
rect 18616 3466 18736 3482
rect 18604 3460 18736 3466
rect 18656 3454 18736 3460
rect 18604 3402 18656 3408
rect 18800 3058 18828 3878
rect 19260 3738 19288 4082
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19352 3210 19380 4082
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19260 3194 19380 3210
rect 19248 3188 19380 3194
rect 19300 3182 19380 3188
rect 19248 3130 19300 3136
rect 19444 3126 19472 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19708 3120 19760 3126
rect 19708 3062 19760 3068
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19340 2984 19392 2990
rect 19246 2952 19302 2961
rect 19720 2972 19748 3062
rect 19996 2990 20024 3470
rect 20088 3369 20116 3606
rect 20168 3392 20220 3398
rect 20074 3360 20130 3369
rect 20168 3334 20220 3340
rect 20074 3295 20130 3304
rect 19392 2944 19748 2972
rect 19984 2984 20036 2990
rect 19340 2926 19392 2932
rect 19984 2926 20036 2932
rect 19246 2887 19302 2896
rect 19260 2854 19288 2887
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 20180 2446 20208 3334
rect 20272 3210 20300 4558
rect 20364 3380 20392 12406
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 20456 3602 20484 4694
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 21100 4282 21128 4558
rect 21732 4480 21784 4486
rect 21732 4422 21784 4428
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 20548 3534 20576 3878
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20640 3398 20668 3878
rect 20824 3738 20852 4082
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20916 3777 20944 3878
rect 20902 3768 20958 3777
rect 20812 3732 20864 3738
rect 21468 3738 21496 4150
rect 20902 3703 20958 3712
rect 21456 3732 21508 3738
rect 20812 3674 20864 3680
rect 21456 3674 21508 3680
rect 20628 3392 20680 3398
rect 20364 3352 20576 3380
rect 20272 3182 20484 3210
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20168 2440 20220 2446
rect 18432 2366 18736 2394
rect 20168 2382 20220 2388
rect 18708 800 18736 2366
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19340 1556 19392 1562
rect 19340 1498 19392 1504
rect 19352 800 19380 1498
rect 19996 870 20208 898
rect 19996 800 20024 870
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20180 762 20208 870
rect 20364 762 20392 2926
rect 20456 2650 20484 3182
rect 20548 2774 20576 3352
rect 20628 3334 20680 3340
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20732 2961 20760 3334
rect 21744 3058 21772 4422
rect 22296 4146 22324 4422
rect 22480 4282 22508 4558
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 21928 3058 21956 4082
rect 22112 3602 22508 3618
rect 22112 3596 22520 3602
rect 22112 3590 22468 3596
rect 22112 3398 22140 3590
rect 22468 3538 22520 3544
rect 22664 3534 22692 4422
rect 22848 3942 22876 20946
rect 23032 4049 23060 28494
rect 23216 27946 23244 28494
rect 23860 28422 23888 29446
rect 23848 28416 23900 28422
rect 23848 28358 23900 28364
rect 23664 28076 23716 28082
rect 23664 28018 23716 28024
rect 23204 27940 23256 27946
rect 23204 27882 23256 27888
rect 23216 27538 23244 27882
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23400 26518 23428 26862
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23492 26382 23520 26726
rect 23676 26518 23704 28018
rect 23848 27396 23900 27402
rect 23848 27338 23900 27344
rect 23860 26994 23888 27338
rect 23756 26988 23808 26994
rect 23756 26930 23808 26936
rect 23848 26988 23900 26994
rect 23848 26930 23900 26936
rect 23768 26518 23796 26930
rect 23664 26512 23716 26518
rect 23664 26454 23716 26460
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 23768 26382 23796 26454
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23756 26376 23808 26382
rect 23756 26318 23808 26324
rect 23848 26240 23900 26246
rect 23848 26182 23900 26188
rect 23572 25968 23624 25974
rect 23572 25910 23624 25916
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 23308 25498 23336 25774
rect 23296 25492 23348 25498
rect 23296 25434 23348 25440
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23296 24676 23348 24682
rect 23296 24618 23348 24624
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23216 23322 23244 23666
rect 23204 23316 23256 23322
rect 23204 23258 23256 23264
rect 23308 22982 23336 24618
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 20466 23336 22918
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23400 18766 23428 19314
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23400 17202 23428 18702
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23112 16176 23164 16182
rect 23112 16118 23164 16124
rect 23124 15706 23152 16118
rect 23400 15706 23428 16458
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23492 5098 23520 25230
rect 23584 24818 23612 25910
rect 23664 25424 23716 25430
rect 23664 25366 23716 25372
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23676 24750 23704 25366
rect 23860 25294 23888 26182
rect 23848 25288 23900 25294
rect 23848 25230 23900 25236
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23940 23112 23992 23118
rect 23940 23054 23992 23060
rect 23952 22642 23980 23054
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23768 19378 23796 20198
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23676 17270 23704 17478
rect 23860 17270 23888 18158
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23584 16250 23612 16458
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23584 15638 23612 16186
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 23676 15434 23704 16662
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23860 15094 23888 16390
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23952 14958 23980 15438
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 23480 5092 23532 5098
rect 23480 5034 23532 5040
rect 23018 4040 23074 4049
rect 23018 3975 23074 3984
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 23848 3936 23900 3942
rect 23848 3878 23900 3884
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 20718 2952 20774 2961
rect 20718 2887 20774 2896
rect 20548 2746 20668 2774
rect 20640 2650 20668 2746
rect 22296 2650 22324 3470
rect 22756 3058 22784 3470
rect 22940 3126 22968 3878
rect 23860 3602 23888 3878
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23032 2990 23060 3062
rect 23020 2984 23072 2990
rect 23020 2926 23072 2932
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 20640 800 20668 2314
rect 21928 800 21956 2314
rect 23124 898 23152 2926
rect 23492 2650 23520 2926
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 24044 2514 24072 31726
rect 24214 31512 24270 31521
rect 24214 31447 24270 31456
rect 24228 31414 24256 31447
rect 24216 31408 24268 31414
rect 24216 31350 24268 31356
rect 24124 25832 24176 25838
rect 24124 25774 24176 25780
rect 24136 25226 24164 25774
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 24320 24342 24348 32370
rect 24412 32026 24440 32846
rect 24400 32020 24452 32026
rect 24400 31962 24452 31968
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24412 30036 24440 30194
rect 24504 30190 24532 34138
rect 24596 33998 24624 35702
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 24676 35556 24728 35562
rect 24676 35498 24728 35504
rect 24688 34202 24716 35498
rect 24780 35018 24808 35566
rect 24768 35012 24820 35018
rect 24768 34954 24820 34960
rect 24676 34196 24728 34202
rect 24676 34138 24728 34144
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24596 33522 24624 33934
rect 24584 33516 24636 33522
rect 24584 33458 24636 33464
rect 24596 31482 24624 33458
rect 24872 33046 24900 36518
rect 25148 36310 25176 37198
rect 25792 36922 25820 43726
rect 28828 41414 28856 46922
rect 28736 41386 28856 41414
rect 25964 37936 26016 37942
rect 25964 37878 26016 37884
rect 25976 37262 26004 37878
rect 27804 37868 27856 37874
rect 27804 37810 27856 37816
rect 26332 37664 26384 37670
rect 26332 37606 26384 37612
rect 26344 37262 26372 37606
rect 25964 37256 26016 37262
rect 25964 37198 26016 37204
rect 26332 37256 26384 37262
rect 26332 37198 26384 37204
rect 25780 36916 25832 36922
rect 25780 36858 25832 36864
rect 25228 36780 25280 36786
rect 25228 36722 25280 36728
rect 24952 36304 25004 36310
rect 24952 36246 25004 36252
rect 25136 36304 25188 36310
rect 25136 36246 25188 36252
rect 24964 35290 24992 36246
rect 25240 36242 25268 36722
rect 25228 36236 25280 36242
rect 25228 36178 25280 36184
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 25148 35834 25176 36042
rect 25136 35828 25188 35834
rect 25136 35770 25188 35776
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 24952 35148 25004 35154
rect 24952 35090 25004 35096
rect 24860 33040 24912 33046
rect 24860 32982 24912 32988
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24780 32502 24808 32846
rect 24768 32496 24820 32502
rect 24768 32438 24820 32444
rect 24676 32360 24728 32366
rect 24676 32302 24728 32308
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 24492 30184 24544 30190
rect 24544 30132 24624 30138
rect 24492 30126 24624 30132
rect 24504 30110 24624 30126
rect 24492 30048 24544 30054
rect 24412 30008 24492 30036
rect 24492 29990 24544 29996
rect 24504 29646 24532 29990
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24596 27946 24624 30110
rect 24688 28218 24716 32302
rect 24766 31512 24822 31521
rect 24766 31447 24822 31456
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24780 28098 24808 31447
rect 24872 30326 24900 32982
rect 24860 30320 24912 30326
rect 24860 30262 24912 30268
rect 24688 28070 24808 28098
rect 24584 27940 24636 27946
rect 24584 27882 24636 27888
rect 24688 26450 24716 28070
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24780 26450 24808 27270
rect 24872 26926 24900 30262
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24400 26444 24452 26450
rect 24400 26386 24452 26392
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24412 26042 24440 26386
rect 24400 26036 24452 26042
rect 24400 25978 24452 25984
rect 24780 25906 24808 26386
rect 24872 25974 24900 26726
rect 24860 25968 24912 25974
rect 24860 25910 24912 25916
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24308 24336 24360 24342
rect 24308 24278 24360 24284
rect 24780 24206 24808 24686
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24780 22778 24808 22986
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24688 21962 24716 22578
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21622 24440 21830
rect 24688 21690 24716 21898
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 24308 21480 24360 21486
rect 24308 21422 24360 21428
rect 24320 21010 24348 21422
rect 24308 21004 24360 21010
rect 24308 20946 24360 20952
rect 24688 20466 24716 21626
rect 24872 21010 24900 21966
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 24858 19408 24914 19417
rect 24858 19343 24914 19352
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24412 16658 24440 17614
rect 24872 16998 24900 19343
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24872 16590 24900 16730
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24872 16130 24900 16526
rect 24780 16102 24900 16130
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24136 15570 24164 15982
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24688 14618 24716 15506
rect 24780 15502 24808 16102
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24872 15706 24900 15982
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24584 9988 24636 9994
rect 24584 9930 24636 9936
rect 24596 9722 24624 9930
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24412 3126 24440 9522
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24688 3369 24716 3470
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 24674 3360 24730 3369
rect 24674 3295 24730 3304
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24122 2952 24178 2961
rect 24122 2887 24124 2896
rect 24176 2887 24178 2896
rect 24124 2858 24176 2864
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 22572 870 22784 898
rect 22572 800 22600 870
rect 20180 734 20392 762
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 22756 762 22784 870
rect 23032 870 23152 898
rect 23032 762 23060 870
rect 23216 800 23244 2382
rect 24504 800 24532 2994
rect 24780 2514 24808 3402
rect 24964 2650 24992 35090
rect 25044 34672 25096 34678
rect 25044 34614 25096 34620
rect 25056 31890 25084 34614
rect 25044 31884 25096 31890
rect 25044 31826 25096 31832
rect 25056 31482 25084 31826
rect 25240 31686 25268 36178
rect 25412 35284 25464 35290
rect 25412 35226 25464 35232
rect 25424 35086 25452 35226
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 25596 35080 25648 35086
rect 25596 35022 25648 35028
rect 25608 34678 25636 35022
rect 25596 34672 25648 34678
rect 25596 34614 25648 34620
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25424 33930 25452 34478
rect 25412 33924 25464 33930
rect 25412 33866 25464 33872
rect 25596 33448 25648 33454
rect 25596 33390 25648 33396
rect 25608 33318 25636 33390
rect 25596 33312 25648 33318
rect 25596 33254 25648 33260
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 25700 32842 25728 33254
rect 25596 32836 25648 32842
rect 25596 32778 25648 32784
rect 25688 32836 25740 32842
rect 25688 32778 25740 32784
rect 25608 32570 25636 32778
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 25228 31680 25280 31686
rect 25228 31622 25280 31628
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 25056 28150 25084 31418
rect 25240 31346 25268 31622
rect 25608 31414 25636 32506
rect 25688 31748 25740 31754
rect 25688 31690 25740 31696
rect 25596 31408 25648 31414
rect 25596 31350 25648 31356
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 25228 31204 25280 31210
rect 25228 31146 25280 31152
rect 25240 30938 25268 31146
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 25136 30864 25188 30870
rect 25136 30806 25188 30812
rect 25148 30598 25176 30806
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25136 30592 25188 30598
rect 25136 30534 25188 30540
rect 25148 30394 25176 30534
rect 25136 30388 25188 30394
rect 25136 30330 25188 30336
rect 25136 30184 25188 30190
rect 25136 30126 25188 30132
rect 25148 29850 25176 30126
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 25136 29164 25188 29170
rect 25136 29106 25188 29112
rect 25148 28966 25176 29106
rect 25608 29102 25636 30670
rect 25700 30666 25728 31690
rect 25688 30660 25740 30666
rect 25688 30602 25740 30608
rect 25700 30394 25728 30602
rect 25688 30388 25740 30394
rect 25688 30330 25740 30336
rect 25688 29504 25740 29510
rect 25688 29446 25740 29452
rect 25700 29170 25728 29446
rect 25688 29164 25740 29170
rect 25688 29106 25740 29112
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 25044 28144 25096 28150
rect 25044 28086 25096 28092
rect 25056 27470 25084 28086
rect 25148 27878 25176 28902
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25044 27464 25096 27470
rect 25044 27406 25096 27412
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25136 26240 25188 26246
rect 25136 26182 25188 26188
rect 25044 25696 25096 25702
rect 25044 25638 25096 25644
rect 25056 25226 25084 25638
rect 25148 25498 25176 26182
rect 25240 25498 25268 27338
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25240 22030 25268 23462
rect 25332 22094 25360 25842
rect 25596 25220 25648 25226
rect 25596 25162 25648 25168
rect 25608 24818 25636 25162
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25412 24064 25464 24070
rect 25412 24006 25464 24012
rect 25424 23050 25452 24006
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25596 22500 25648 22506
rect 25596 22442 25648 22448
rect 25332 22066 25452 22094
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25042 20360 25098 20369
rect 25042 20295 25044 20304
rect 25096 20295 25098 20304
rect 25044 20266 25096 20272
rect 25044 18692 25096 18698
rect 25044 18634 25096 18640
rect 25056 18222 25084 18634
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17746 25084 18022
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16794 25084 16934
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25148 4146 25176 21626
rect 25240 18902 25268 21966
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25332 21622 25360 21830
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25332 20262 25360 20810
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25332 19174 25360 20198
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25228 18896 25280 18902
rect 25228 18838 25280 18844
rect 25332 18766 25360 19110
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25240 18290 25268 18566
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25332 17746 25360 18022
rect 25320 17740 25372 17746
rect 25320 17682 25372 17688
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25240 14482 25268 15370
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25136 4140 25188 4146
rect 25136 4082 25188 4088
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 25240 3942 25268 4082
rect 25332 4078 25360 17070
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 25044 3460 25096 3466
rect 25044 3402 25096 3408
rect 25056 3369 25084 3402
rect 25042 3360 25098 3369
rect 25042 3295 25098 3304
rect 25424 3126 25452 22066
rect 25608 21690 25636 22442
rect 25792 22094 25820 36858
rect 26344 35766 26372 37198
rect 26976 37188 27028 37194
rect 26976 37130 27028 37136
rect 26988 36922 27016 37130
rect 27816 37126 27844 37810
rect 27988 37664 28040 37670
rect 27988 37606 28040 37612
rect 28000 37194 28028 37606
rect 27988 37188 28040 37194
rect 27988 37130 28040 37136
rect 27804 37120 27856 37126
rect 27804 37062 27856 37068
rect 28448 37120 28500 37126
rect 28448 37062 28500 37068
rect 27816 36922 27844 37062
rect 26976 36916 27028 36922
rect 26976 36858 27028 36864
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 27540 36786 27936 36802
rect 27252 36780 27304 36786
rect 27252 36722 27304 36728
rect 27528 36780 27936 36786
rect 27580 36774 27936 36780
rect 27528 36722 27580 36728
rect 27264 35834 27292 36722
rect 27528 36644 27580 36650
rect 27528 36586 27580 36592
rect 27540 36106 27568 36586
rect 27528 36100 27580 36106
rect 27528 36042 27580 36048
rect 27540 35850 27568 36042
rect 27804 36032 27856 36038
rect 27804 35974 27856 35980
rect 27252 35828 27304 35834
rect 27252 35770 27304 35776
rect 27448 35822 27568 35850
rect 27816 35834 27844 35974
rect 27804 35828 27856 35834
rect 26332 35760 26384 35766
rect 26332 35702 26384 35708
rect 26976 35692 27028 35698
rect 26976 35634 27028 35640
rect 26332 35624 26384 35630
rect 26332 35566 26384 35572
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26252 35154 26280 35430
rect 26344 35222 26372 35566
rect 26424 35488 26476 35494
rect 26424 35430 26476 35436
rect 26436 35290 26464 35430
rect 26424 35284 26476 35290
rect 26424 35226 26476 35232
rect 26332 35216 26384 35222
rect 26332 35158 26384 35164
rect 26240 35148 26292 35154
rect 26240 35090 26292 35096
rect 26148 34944 26200 34950
rect 26148 34886 26200 34892
rect 26160 33998 26188 34886
rect 26344 34746 26372 35158
rect 26436 35086 26464 35226
rect 26424 35080 26476 35086
rect 26424 35022 26476 35028
rect 26514 34776 26570 34785
rect 26332 34740 26384 34746
rect 26514 34711 26570 34720
rect 26332 34682 26384 34688
rect 26528 34678 26556 34711
rect 26516 34672 26568 34678
rect 26516 34614 26568 34620
rect 26988 34610 27016 35634
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 27068 35012 27120 35018
rect 27068 34954 27120 34960
rect 27080 34746 27108 34954
rect 27068 34740 27120 34746
rect 27068 34682 27120 34688
rect 26976 34604 27028 34610
rect 26976 34546 27028 34552
rect 26240 34536 26292 34542
rect 26240 34478 26292 34484
rect 26252 33998 26280 34478
rect 26988 34474 27016 34546
rect 26516 34468 26568 34474
rect 26344 34428 26516 34456
rect 26148 33992 26200 33998
rect 26148 33934 26200 33940
rect 26240 33992 26292 33998
rect 26240 33934 26292 33940
rect 25964 33856 26016 33862
rect 25964 33798 26016 33804
rect 26148 33856 26200 33862
rect 26344 33810 26372 34428
rect 26516 34410 26568 34416
rect 26976 34468 27028 34474
rect 26976 34410 27028 34416
rect 27080 34406 27108 34682
rect 27172 34610 27200 35022
rect 27448 34746 27476 35822
rect 27804 35770 27856 35776
rect 27528 35760 27580 35766
rect 27528 35702 27580 35708
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 26884 34400 26936 34406
rect 26884 34342 26936 34348
rect 27068 34400 27120 34406
rect 27068 34342 27120 34348
rect 26896 33998 26924 34342
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26148 33798 26200 33804
rect 25976 33522 26004 33798
rect 26160 33522 26188 33798
rect 26252 33782 26372 33810
rect 25964 33516 26016 33522
rect 25964 33458 26016 33464
rect 26148 33516 26200 33522
rect 26148 33458 26200 33464
rect 26056 33448 26108 33454
rect 26056 33390 26108 33396
rect 25964 31816 26016 31822
rect 25964 31758 26016 31764
rect 25976 31346 26004 31758
rect 25964 31340 26016 31346
rect 25964 31282 26016 31288
rect 25872 30252 25924 30258
rect 25872 30194 25924 30200
rect 25884 24954 25912 30194
rect 25976 30122 26004 31282
rect 26068 30598 26096 33390
rect 26148 32564 26200 32570
rect 26148 32506 26200 32512
rect 26160 31686 26188 32506
rect 26148 31680 26200 31686
rect 26148 31622 26200 31628
rect 26160 31521 26188 31622
rect 26146 31512 26202 31521
rect 26146 31447 26202 31456
rect 26252 30938 26280 33782
rect 27080 33096 27108 34342
rect 26896 33068 27108 33096
rect 26332 32020 26384 32026
rect 26332 31962 26384 31968
rect 26344 31278 26372 31962
rect 26332 31272 26384 31278
rect 26332 31214 26384 31220
rect 26240 30932 26292 30938
rect 26240 30874 26292 30880
rect 26608 30796 26660 30802
rect 26608 30738 26660 30744
rect 26620 30598 26648 30738
rect 26056 30592 26108 30598
rect 26056 30534 26108 30540
rect 26608 30592 26660 30598
rect 26608 30534 26660 30540
rect 26792 30592 26844 30598
rect 26792 30534 26844 30540
rect 25964 30116 26016 30122
rect 25964 30058 26016 30064
rect 25976 26314 26004 30058
rect 26332 29572 26384 29578
rect 26332 29514 26384 29520
rect 26344 29306 26372 29514
rect 26804 29510 26832 30534
rect 26896 29510 26924 33068
rect 27172 33046 27200 34546
rect 27344 34060 27396 34066
rect 27344 34002 27396 34008
rect 27160 33040 27212 33046
rect 27160 32982 27212 32988
rect 26976 32972 27028 32978
rect 26976 32914 27028 32920
rect 26988 31890 27016 32914
rect 27356 32910 27384 34002
rect 27448 33998 27476 34682
rect 27540 34134 27568 35702
rect 27816 35086 27844 35770
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27528 34128 27580 34134
rect 27528 34070 27580 34076
rect 27436 33992 27488 33998
rect 27436 33934 27488 33940
rect 27540 33674 27568 34070
rect 27448 33658 27568 33674
rect 27448 33652 27580 33658
rect 27448 33646 27528 33652
rect 27448 32978 27476 33646
rect 27528 33594 27580 33600
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27436 32972 27488 32978
rect 27436 32914 27488 32920
rect 27344 32904 27396 32910
rect 27344 32846 27396 32852
rect 27436 32836 27488 32842
rect 27436 32778 27488 32784
rect 27344 32292 27396 32298
rect 27344 32234 27396 32240
rect 27252 32224 27304 32230
rect 27252 32166 27304 32172
rect 27264 31890 27292 32166
rect 27356 31890 27384 32234
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 27344 31884 27396 31890
rect 27344 31826 27396 31832
rect 27448 30938 27476 32778
rect 27540 31414 27568 33458
rect 27908 32774 27936 36774
rect 28460 36718 28488 37062
rect 27988 36712 28040 36718
rect 27988 36654 28040 36660
rect 28448 36712 28500 36718
rect 28448 36654 28500 36660
rect 28000 36174 28028 36654
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 28000 35698 28028 36110
rect 27988 35692 28040 35698
rect 27988 35634 28040 35640
rect 28000 35290 28028 35634
rect 28356 35488 28408 35494
rect 28356 35430 28408 35436
rect 27988 35284 28040 35290
rect 27988 35226 28040 35232
rect 28368 33522 28396 35430
rect 28448 35080 28500 35086
rect 28448 35022 28500 35028
rect 28356 33516 28408 33522
rect 28356 33458 28408 33464
rect 28172 32904 28224 32910
rect 28172 32846 28224 32852
rect 27896 32768 27948 32774
rect 27896 32710 27948 32716
rect 27908 32450 27936 32710
rect 27816 32434 27936 32450
rect 27804 32428 27936 32434
rect 27856 32422 27936 32428
rect 27804 32370 27856 32376
rect 27896 32360 27948 32366
rect 27896 32302 27948 32308
rect 27712 32224 27764 32230
rect 27712 32166 27764 32172
rect 27528 31408 27580 31414
rect 27528 31350 27580 31356
rect 27436 30932 27488 30938
rect 27436 30874 27488 30880
rect 26976 30660 27028 30666
rect 26976 30602 27028 30608
rect 26792 29504 26844 29510
rect 26792 29446 26844 29452
rect 26884 29504 26936 29510
rect 26884 29446 26936 29452
rect 26332 29300 26384 29306
rect 26332 29242 26384 29248
rect 26516 29232 26568 29238
rect 26516 29174 26568 29180
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26068 28694 26096 29106
rect 26056 28688 26108 28694
rect 26056 28630 26108 28636
rect 26068 27606 26096 28630
rect 26056 27600 26108 27606
rect 26056 27542 26108 27548
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25884 23730 25912 24890
rect 25872 23724 25924 23730
rect 25872 23666 25924 23672
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 26160 22642 26188 22918
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 26160 22234 26188 22578
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 25964 22160 26016 22166
rect 25964 22102 26016 22108
rect 25700 22066 25820 22094
rect 25700 22030 25728 22066
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25976 21978 26004 22102
rect 26252 21978 26280 26318
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25700 21434 25728 21966
rect 25976 21950 26280 21978
rect 25608 21406 25728 21434
rect 25608 21010 25636 21406
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25700 21078 25728 21286
rect 25688 21072 25740 21078
rect 25688 21014 25740 21020
rect 25976 21010 26004 21286
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25964 21004 26016 21010
rect 25964 20946 26016 20952
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25516 20777 25544 20878
rect 25502 20768 25558 20777
rect 25502 20703 25558 20712
rect 25608 20602 25636 20946
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 25870 20768 25926 20777
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25792 20534 25820 20742
rect 25870 20703 25926 20712
rect 25884 20534 25912 20703
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 25872 20528 25924 20534
rect 25872 20470 25924 20476
rect 25596 20324 25648 20330
rect 25596 20266 25648 20272
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25608 19990 25636 20266
rect 25596 19984 25648 19990
rect 25596 19926 25648 19932
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 25516 18698 25544 19110
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25608 18578 25636 19926
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25700 19417 25728 19790
rect 25792 19786 25820 20266
rect 25976 19990 26004 20946
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26068 20602 26096 20878
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 25964 19984 26016 19990
rect 25964 19926 26016 19932
rect 25780 19780 25832 19786
rect 25780 19722 25832 19728
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25884 19553 25912 19722
rect 25870 19544 25926 19553
rect 25870 19479 25926 19488
rect 26160 19446 26188 20810
rect 26252 19854 26280 21950
rect 26330 20360 26386 20369
rect 26330 20295 26386 20304
rect 26344 20262 26372 20295
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 25872 19440 25924 19446
rect 25686 19408 25742 19417
rect 25872 19382 25924 19388
rect 26148 19440 26200 19446
rect 26148 19382 26200 19388
rect 25686 19343 25742 19352
rect 25884 18970 25912 19382
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25780 18896 25832 18902
rect 25780 18838 25832 18844
rect 25792 18766 25820 18838
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25516 18550 25636 18578
rect 25516 10130 25544 18550
rect 25792 17202 25820 18702
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25884 18358 25912 18566
rect 25872 18352 25924 18358
rect 25872 18294 25924 18300
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 25884 16946 25912 18294
rect 26068 18290 26096 19314
rect 26344 19242 26372 19722
rect 26332 19236 26384 19242
rect 26332 19178 26384 19184
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26068 17762 26096 18226
rect 25700 16918 25912 16946
rect 25976 17734 26096 17762
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25608 16454 25636 16526
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25700 15366 25728 16918
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25792 16590 25820 16730
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25792 15502 25820 16526
rect 25872 16516 25924 16522
rect 25872 16458 25924 16464
rect 25884 16250 25912 16458
rect 25976 16454 26004 17734
rect 26056 17604 26108 17610
rect 26056 17546 26108 17552
rect 26068 17338 26096 17546
rect 26056 17332 26108 17338
rect 26056 17274 26108 17280
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26068 16674 26096 17138
rect 26068 16646 26188 16674
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 25976 16266 26004 16390
rect 25872 16244 25924 16250
rect 25976 16238 26096 16266
rect 25872 16186 25924 16192
rect 25964 16176 26016 16182
rect 25964 16118 26016 16124
rect 25780 15496 25832 15502
rect 25780 15438 25832 15444
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25700 15094 25728 15302
rect 25688 15088 25740 15094
rect 25688 15030 25740 15036
rect 25792 14414 25820 15438
rect 25976 15162 26004 16118
rect 26068 15434 26096 16238
rect 26160 16114 26188 16646
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 25964 15156 26016 15162
rect 25964 15098 26016 15104
rect 26160 15026 26188 16050
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 25516 2582 25544 3470
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 25504 2576 25556 2582
rect 25504 2518 25556 2524
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 800 25176 2450
rect 25608 1562 25636 2926
rect 26160 2378 26188 10066
rect 26436 3942 26464 29106
rect 26528 28218 26556 29174
rect 26896 29102 26924 29446
rect 26988 29170 27016 30602
rect 27540 30326 27568 31350
rect 27528 30320 27580 30326
rect 27528 30262 27580 30268
rect 27252 30116 27304 30122
rect 27252 30058 27304 30064
rect 27264 29714 27292 30058
rect 27252 29708 27304 29714
rect 27252 29650 27304 29656
rect 27068 29572 27120 29578
rect 27068 29514 27120 29520
rect 27080 29306 27108 29514
rect 27068 29300 27120 29306
rect 27068 29242 27120 29248
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 26884 29096 26936 29102
rect 26884 29038 26936 29044
rect 26516 28212 26568 28218
rect 26516 28154 26568 28160
rect 26528 25974 26556 28154
rect 26608 28008 26660 28014
rect 26608 27950 26660 27956
rect 26620 27402 26648 27950
rect 26884 27872 26936 27878
rect 26884 27814 26936 27820
rect 26608 27396 26660 27402
rect 26608 27338 26660 27344
rect 26620 26518 26648 27338
rect 26896 26926 26924 27814
rect 27264 27062 27292 29650
rect 27528 27328 27580 27334
rect 27528 27270 27580 27276
rect 27540 27062 27568 27270
rect 27252 27056 27304 27062
rect 27252 26998 27304 27004
rect 27528 27056 27580 27062
rect 27528 26998 27580 27004
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26608 26512 26660 26518
rect 26608 26454 26660 26460
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 27264 25906 27292 26998
rect 27436 26308 27488 26314
rect 27436 26250 27488 26256
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27264 25362 27292 25842
rect 27344 25832 27396 25838
rect 27344 25774 27396 25780
rect 27252 25356 27304 25362
rect 27252 25298 27304 25304
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26528 22710 26556 24142
rect 26804 23866 26832 24754
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 26804 23118 26832 23802
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 26988 22778 27016 22986
rect 27356 22778 27384 25774
rect 26976 22772 27028 22778
rect 26976 22714 27028 22720
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 26516 22704 26568 22710
rect 27356 22658 27384 22714
rect 26516 22646 26568 22652
rect 27264 22630 27384 22658
rect 27264 21554 27292 22630
rect 27448 22094 27476 26250
rect 27528 25152 27580 25158
rect 27528 25094 27580 25100
rect 27540 24750 27568 25094
rect 27528 24744 27580 24750
rect 27528 24686 27580 24692
rect 27724 22094 27752 32166
rect 27908 31482 27936 32302
rect 27896 31476 27948 31482
rect 27896 31418 27948 31424
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 28000 29782 28028 31282
rect 28184 30054 28212 32846
rect 28264 32768 28316 32774
rect 28264 32710 28316 32716
rect 28276 31822 28304 32710
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28368 31278 28396 33458
rect 28460 31482 28488 35022
rect 28632 34944 28684 34950
rect 28632 34886 28684 34892
rect 28644 34610 28672 34886
rect 28632 34604 28684 34610
rect 28632 34546 28684 34552
rect 28540 34536 28592 34542
rect 28540 34478 28592 34484
rect 28448 31476 28500 31482
rect 28448 31418 28500 31424
rect 28356 31272 28408 31278
rect 28356 31214 28408 31220
rect 28552 30190 28580 34478
rect 28632 33380 28684 33386
rect 28632 33322 28684 33328
rect 28644 31822 28672 33322
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28632 30252 28684 30258
rect 28632 30194 28684 30200
rect 28540 30184 28592 30190
rect 28540 30126 28592 30132
rect 28172 30048 28224 30054
rect 28172 29990 28224 29996
rect 27988 29776 28040 29782
rect 27988 29718 28040 29724
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 27908 26790 27936 27406
rect 28000 27334 28028 29718
rect 28184 29510 28212 29990
rect 28644 29850 28672 30194
rect 28632 29844 28684 29850
rect 28632 29786 28684 29792
rect 28172 29504 28224 29510
rect 28172 29446 28224 29452
rect 28080 28008 28132 28014
rect 28080 27950 28132 27956
rect 28092 27470 28120 27950
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 27988 27328 28040 27334
rect 27988 27270 28040 27276
rect 28092 27130 28120 27406
rect 28080 27124 28132 27130
rect 28080 27066 28132 27072
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27908 25294 27936 26726
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 28644 26314 28672 26522
rect 28632 26308 28684 26314
rect 28632 26250 28684 26256
rect 27988 26240 28040 26246
rect 27988 26182 28040 26188
rect 28000 25974 28028 26182
rect 27988 25968 28040 25974
rect 27988 25910 28040 25916
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 27908 24954 27936 25230
rect 27804 24948 27856 24954
rect 27804 24890 27856 24896
rect 27896 24948 27948 24954
rect 27896 24890 27948 24896
rect 27816 24818 27844 24890
rect 27804 24812 27856 24818
rect 27804 24754 27856 24760
rect 27896 24676 27948 24682
rect 27896 24618 27948 24624
rect 27908 24342 27936 24618
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 27896 24336 27948 24342
rect 27896 24278 27948 24284
rect 28276 23798 28304 24550
rect 28264 23792 28316 23798
rect 28264 23734 28316 23740
rect 27896 23724 27948 23730
rect 27896 23666 27948 23672
rect 27908 23594 27936 23666
rect 27896 23588 27948 23594
rect 27896 23530 27948 23536
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 27816 22778 27844 23122
rect 27804 22772 27856 22778
rect 27804 22714 27856 22720
rect 27908 22438 27936 23530
rect 27988 23180 28040 23186
rect 27988 23122 28040 23128
rect 27896 22432 27948 22438
rect 27896 22374 27948 22380
rect 27356 22066 27476 22094
rect 27632 22066 27752 22094
rect 26884 21548 26936 21554
rect 26884 21490 26936 21496
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 26516 20528 26568 20534
rect 26516 20470 26568 20476
rect 26528 19718 26556 20470
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26804 19378 26832 19654
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26516 19304 26568 19310
rect 26516 19246 26568 19252
rect 26528 18222 26556 19246
rect 26896 18766 26924 21490
rect 27160 21480 27212 21486
rect 27160 21422 27212 21428
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26988 20602 27016 20878
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 27172 20466 27200 21422
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 27172 20330 27200 20402
rect 27160 20324 27212 20330
rect 27160 20266 27212 20272
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 26804 17882 26832 18158
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26804 15910 26832 17818
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27172 15434 27200 15846
rect 26608 15428 26660 15434
rect 26608 15370 26660 15376
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 26620 15162 26648 15370
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 27356 8838 27384 22066
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27448 20942 27476 21966
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27540 16658 27568 17138
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27632 10742 27660 22066
rect 27896 22024 27948 22030
rect 27896 21966 27948 21972
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27724 21010 27752 21830
rect 27908 21350 27936 21966
rect 27896 21344 27948 21350
rect 27896 21286 27948 21292
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27724 20466 27752 20946
rect 27908 20942 27936 21286
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27908 20466 27936 20742
rect 28000 20534 28028 23122
rect 28448 21888 28500 21894
rect 28448 21830 28500 21836
rect 28460 21554 28488 21830
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28736 20874 28764 41386
rect 28998 35728 29054 35737
rect 28998 35663 29054 35672
rect 28908 35488 28960 35494
rect 28908 35430 28960 35436
rect 28920 35018 28948 35430
rect 29012 35018 29040 35663
rect 28908 35012 28960 35018
rect 28908 34954 28960 34960
rect 29000 35012 29052 35018
rect 29000 34954 29052 34960
rect 28920 34610 28948 34954
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 29012 32774 29040 34954
rect 29000 32768 29052 32774
rect 29000 32710 29052 32716
rect 28816 32360 28868 32366
rect 28816 32302 28868 32308
rect 28828 31958 28856 32302
rect 28908 32292 28960 32298
rect 28908 32234 28960 32240
rect 28816 31952 28868 31958
rect 28816 31894 28868 31900
rect 28828 31346 28856 31894
rect 28920 31482 28948 32234
rect 29000 32224 29052 32230
rect 29000 32166 29052 32172
rect 29012 31890 29040 32166
rect 29000 31884 29052 31890
rect 29000 31826 29052 31832
rect 29000 31680 29052 31686
rect 29000 31622 29052 31628
rect 28908 31476 28960 31482
rect 28908 31418 28960 31424
rect 29012 31346 29040 31622
rect 28816 31340 28868 31346
rect 28816 31282 28868 31288
rect 29000 31340 29052 31346
rect 29000 31282 29052 31288
rect 29012 30598 29040 31282
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 29000 30388 29052 30394
rect 29000 30330 29052 30336
rect 29012 30190 29040 30330
rect 29000 30184 29052 30190
rect 29000 30126 29052 30132
rect 29000 29776 29052 29782
rect 29000 29718 29052 29724
rect 29012 28422 29040 29718
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29012 28218 29040 28358
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 28816 27328 28868 27334
rect 28816 27270 28868 27276
rect 28828 26314 28856 27270
rect 28816 26308 28868 26314
rect 28816 26250 28868 26256
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 28920 22098 28948 25230
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28828 21622 28856 21830
rect 28816 21616 28868 21622
rect 28816 21558 28868 21564
rect 28920 20942 28948 22034
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 28172 20800 28224 20806
rect 28172 20742 28224 20748
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28184 20534 28212 20742
rect 27988 20528 28040 20534
rect 27988 20470 28040 20476
rect 28172 20528 28224 20534
rect 28172 20470 28224 20476
rect 28552 20466 28580 20742
rect 29012 20602 29040 21966
rect 29000 20596 29052 20602
rect 29000 20538 29052 20544
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 28736 17746 28764 18702
rect 29104 18630 29132 47126
rect 29656 47054 29684 49200
rect 30380 47184 30432 47190
rect 30380 47126 30432 47132
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 29380 35766 29408 36518
rect 29368 35760 29420 35766
rect 29368 35702 29420 35708
rect 29368 35624 29420 35630
rect 29368 35566 29420 35572
rect 29380 34746 29408 35566
rect 30392 35086 30420 47126
rect 30944 47054 30972 49200
rect 30932 47048 30984 47054
rect 30932 46990 30984 46996
rect 32232 46442 32260 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 35440 47116 35492 47122
rect 35440 47058 35492 47064
rect 32312 46504 32364 46510
rect 32312 46446 32364 46452
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32324 46170 32352 46446
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 32312 46164 32364 46170
rect 32312 46106 32364 46112
rect 31760 45960 31812 45966
rect 31760 45902 31812 45908
rect 31024 45824 31076 45830
rect 31024 45766 31076 45772
rect 31036 45626 31064 45766
rect 31772 45626 31800 45902
rect 31024 45620 31076 45626
rect 31024 45562 31076 45568
rect 31760 45620 31812 45626
rect 31760 45562 31812 45568
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 31760 44328 31812 44334
rect 31760 44270 31812 44276
rect 31772 43994 31800 44270
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 31760 43988 31812 43994
rect 31760 43930 31812 43936
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35452 35894 35480 47058
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38200 45960 38252 45966
rect 38200 45902 38252 45908
rect 38212 45354 38240 45902
rect 38396 45554 38424 49286
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49200 41318 50000
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 39396 46096 39448 46102
rect 39396 46038 39448 46044
rect 39408 45626 39436 46038
rect 39396 45620 39448 45626
rect 39396 45562 39448 45568
rect 39960 45554 39988 49200
rect 40592 47252 40644 47258
rect 40592 47194 40644 47200
rect 40224 47048 40276 47054
rect 40224 46990 40276 46996
rect 38396 45526 38608 45554
rect 39960 45526 40080 45554
rect 38200 45348 38252 45354
rect 38200 45290 38252 45296
rect 35716 43240 35768 43246
rect 35716 43182 35768 43188
rect 35452 35866 35664 35894
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 29828 35080 29880 35086
rect 29828 35022 29880 35028
rect 30380 35080 30432 35086
rect 30380 35022 30432 35028
rect 29460 34944 29512 34950
rect 29460 34886 29512 34892
rect 29368 34740 29420 34746
rect 29368 34682 29420 34688
rect 29472 34678 29500 34886
rect 29460 34672 29512 34678
rect 29460 34614 29512 34620
rect 29184 34604 29236 34610
rect 29184 34546 29236 34552
rect 29196 32230 29224 34546
rect 29276 34536 29328 34542
rect 29276 34478 29328 34484
rect 29184 32224 29236 32230
rect 29184 32166 29236 32172
rect 29184 30660 29236 30666
rect 29184 30602 29236 30608
rect 29196 29170 29224 30602
rect 29184 29164 29236 29170
rect 29184 29106 29236 29112
rect 29196 26382 29224 29106
rect 29184 26376 29236 26382
rect 29184 26318 29236 26324
rect 29184 18692 29236 18698
rect 29184 18634 29236 18640
rect 29092 18624 29144 18630
rect 29092 18566 29144 18572
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 28724 17740 28776 17746
rect 28724 17682 28776 17688
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 27896 17264 27948 17270
rect 27896 17206 27948 17212
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 27724 16658 27752 17138
rect 27908 16658 27936 17206
rect 27712 16652 27764 16658
rect 27712 16594 27764 16600
rect 27896 16652 27948 16658
rect 27896 16594 27948 16600
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27344 8832 27396 8838
rect 27344 8774 27396 8780
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 27632 3641 27660 4150
rect 27618 3632 27674 3641
rect 27618 3567 27674 3576
rect 27632 3534 27660 3567
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27618 2952 27674 2961
rect 27618 2887 27620 2896
rect 27672 2887 27674 2896
rect 27620 2858 27672 2864
rect 27724 2514 27752 16594
rect 28368 16590 28396 17614
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28552 16522 28580 17614
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28644 17270 28672 17478
rect 28828 17338 28856 17478
rect 28724 17332 28776 17338
rect 28724 17274 28776 17280
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28736 16998 28764 17274
rect 28724 16992 28776 16998
rect 28724 16934 28776 16940
rect 28540 16516 28592 16522
rect 28540 16458 28592 16464
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 28552 16114 28580 16458
rect 28644 16114 28672 16458
rect 28736 16250 28764 16934
rect 29012 16794 29040 18226
rect 29196 17678 29224 18634
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29000 16788 29052 16794
rect 29000 16730 29052 16736
rect 29104 16726 29132 17138
rect 29092 16720 29144 16726
rect 29092 16662 29144 16668
rect 28724 16244 28776 16250
rect 28724 16186 28776 16192
rect 29104 16114 29132 16662
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 27804 10736 27856 10742
rect 27804 10678 27856 10684
rect 27816 2582 27844 10678
rect 28552 4078 28580 16050
rect 28644 4758 28672 16050
rect 28632 4752 28684 4758
rect 28632 4694 28684 4700
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 27908 3398 27936 3538
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28552 3126 28580 4014
rect 29092 3664 29144 3670
rect 29092 3606 29144 3612
rect 27896 3120 27948 3126
rect 27896 3062 27948 3068
rect 28540 3120 28592 3126
rect 28540 3062 28592 3068
rect 27908 2854 27936 3062
rect 29104 2854 29132 3606
rect 29184 3392 29236 3398
rect 29184 3334 29236 3340
rect 29196 3058 29224 3334
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 27896 2848 27948 2854
rect 27896 2790 27948 2796
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 27804 2576 27856 2582
rect 27804 2518 27856 2524
rect 27712 2508 27764 2514
rect 27712 2450 27764 2456
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 25596 1556 25648 1562
rect 25596 1498 25648 1504
rect 26436 800 26464 2382
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 27080 800 27108 2314
rect 28368 800 28396 2382
rect 29288 1970 29316 34478
rect 29368 33584 29420 33590
rect 29368 33526 29420 33532
rect 29380 33114 29408 33526
rect 29368 33108 29420 33114
rect 29368 33050 29420 33056
rect 29472 32858 29500 34614
rect 29840 33998 29868 35022
rect 30748 34944 30800 34950
rect 30748 34886 30800 34892
rect 30760 34610 30788 34886
rect 31392 34672 31444 34678
rect 31392 34614 31444 34620
rect 30748 34604 30800 34610
rect 30748 34546 30800 34552
rect 31024 34604 31076 34610
rect 31024 34546 31076 34552
rect 30564 34400 30616 34406
rect 30564 34342 30616 34348
rect 30576 34202 30604 34342
rect 30380 34196 30432 34202
rect 30380 34138 30432 34144
rect 30564 34196 30616 34202
rect 30564 34138 30616 34144
rect 29920 34060 29972 34066
rect 29972 34020 30052 34048
rect 29920 34002 29972 34008
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29552 33312 29604 33318
rect 29552 33254 29604 33260
rect 29564 32978 29592 33254
rect 29552 32972 29604 32978
rect 29552 32914 29604 32920
rect 29472 32830 29592 32858
rect 29460 32768 29512 32774
rect 29460 32710 29512 32716
rect 29368 32428 29420 32434
rect 29368 32370 29420 32376
rect 29380 31754 29408 32370
rect 29368 31748 29420 31754
rect 29368 31690 29420 31696
rect 29472 29782 29500 32710
rect 29564 30938 29592 32830
rect 29840 32026 29868 33934
rect 30024 33522 30052 34020
rect 30012 33516 30064 33522
rect 30012 33458 30064 33464
rect 29920 33312 29972 33318
rect 29920 33254 29972 33260
rect 29932 33046 29960 33254
rect 29920 33040 29972 33046
rect 29920 32982 29972 32988
rect 29932 32570 29960 32982
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 30024 32434 30052 33458
rect 30288 33040 30340 33046
rect 30288 32982 30340 32988
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 29828 32020 29880 32026
rect 29828 31962 29880 31968
rect 29840 31346 29868 31962
rect 30024 31822 30052 32370
rect 30208 32366 30236 32846
rect 30196 32360 30248 32366
rect 30196 32302 30248 32308
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 29828 31340 29880 31346
rect 29828 31282 29880 31288
rect 30024 31142 30052 31758
rect 30116 31278 30144 31758
rect 30104 31272 30156 31278
rect 30104 31214 30156 31220
rect 30012 31136 30064 31142
rect 30012 31078 30064 31084
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 29552 30932 29604 30938
rect 29552 30874 29604 30880
rect 29920 30864 29972 30870
rect 29920 30806 29972 30812
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 29460 29776 29512 29782
rect 29460 29718 29512 29724
rect 29552 29708 29604 29714
rect 29552 29650 29604 29656
rect 29564 28994 29592 29650
rect 29564 28966 29684 28994
rect 29552 28960 29604 28966
rect 29552 28902 29604 28908
rect 29552 28688 29604 28694
rect 29552 28630 29604 28636
rect 29460 28620 29512 28626
rect 29460 28562 29512 28568
rect 29368 28416 29420 28422
rect 29368 28358 29420 28364
rect 29380 28218 29408 28358
rect 29368 28212 29420 28218
rect 29368 28154 29420 28160
rect 29368 27940 29420 27946
rect 29368 27882 29420 27888
rect 29380 12646 29408 27882
rect 29472 27606 29500 28562
rect 29564 28014 29592 28630
rect 29656 28218 29684 28966
rect 29736 28484 29788 28490
rect 29736 28426 29788 28432
rect 29644 28212 29696 28218
rect 29644 28154 29696 28160
rect 29552 28008 29604 28014
rect 29552 27950 29604 27956
rect 29460 27600 29512 27606
rect 29460 27542 29512 27548
rect 29472 26994 29500 27542
rect 29748 27062 29776 28426
rect 29840 27538 29868 29990
rect 29932 29714 29960 30806
rect 30024 30734 30052 31078
rect 30116 30802 30144 31078
rect 30104 30796 30156 30802
rect 30104 30738 30156 30744
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 30012 29776 30064 29782
rect 30012 29718 30064 29724
rect 29920 29708 29972 29714
rect 29920 29650 29972 29656
rect 30024 29646 30052 29718
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 30208 28762 30236 32302
rect 30300 32026 30328 32982
rect 30392 32978 30420 34138
rect 31036 33862 31064 34546
rect 31024 33856 31076 33862
rect 31024 33798 31076 33804
rect 31404 33386 31432 34614
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 32128 34060 32180 34066
rect 32128 34002 32180 34008
rect 31392 33380 31444 33386
rect 31392 33322 31444 33328
rect 30380 32972 30432 32978
rect 30380 32914 30432 32920
rect 30392 32774 30420 32914
rect 31404 32910 31432 33322
rect 31668 33108 31720 33114
rect 31668 33050 31720 33056
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31484 32904 31536 32910
rect 31484 32846 31536 32852
rect 30380 32768 30432 32774
rect 30380 32710 30432 32716
rect 30932 32292 30984 32298
rect 30932 32234 30984 32240
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 30300 31414 30328 31962
rect 30944 31822 30972 32234
rect 30932 31816 30984 31822
rect 30932 31758 30984 31764
rect 30288 31408 30340 31414
rect 30288 31350 30340 31356
rect 31116 31340 31168 31346
rect 31116 31282 31168 31288
rect 30288 31272 30340 31278
rect 30288 31214 30340 31220
rect 30300 30394 30328 31214
rect 30840 31204 30892 31210
rect 30840 31146 30892 31152
rect 30748 30932 30800 30938
rect 30748 30874 30800 30880
rect 30288 30388 30340 30394
rect 30288 30330 30340 30336
rect 30656 30320 30708 30326
rect 30656 30262 30708 30268
rect 30668 29850 30696 30262
rect 30656 29844 30708 29850
rect 30656 29786 30708 29792
rect 30564 29640 30616 29646
rect 30564 29582 30616 29588
rect 30576 29510 30604 29582
rect 30564 29504 30616 29510
rect 30564 29446 30616 29452
rect 30760 28762 30788 30874
rect 30852 30802 30880 31146
rect 31128 30938 31156 31282
rect 31116 30932 31168 30938
rect 31116 30874 31168 30880
rect 30840 30796 30892 30802
rect 30840 30738 30892 30744
rect 30932 30728 30984 30734
rect 30932 30670 30984 30676
rect 30944 30054 30972 30670
rect 30932 30048 30984 30054
rect 30932 29990 30984 29996
rect 30196 28756 30248 28762
rect 30196 28698 30248 28704
rect 30748 28756 30800 28762
rect 30748 28698 30800 28704
rect 30288 28620 30340 28626
rect 30288 28562 30340 28568
rect 30300 28014 30328 28562
rect 30288 28008 30340 28014
rect 30288 27950 30340 27956
rect 29828 27532 29880 27538
rect 29828 27474 29880 27480
rect 30196 27396 30248 27402
rect 30196 27338 30248 27344
rect 30208 27130 30236 27338
rect 30300 27334 30328 27950
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 30748 27872 30800 27878
rect 30748 27814 30800 27820
rect 30288 27328 30340 27334
rect 30288 27270 30340 27276
rect 30196 27124 30248 27130
rect 30196 27066 30248 27072
rect 29736 27056 29788 27062
rect 29736 26998 29788 27004
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29472 26382 29500 26930
rect 30300 26926 30328 27270
rect 30392 26994 30420 27814
rect 30760 26994 30788 27814
rect 31208 27396 31260 27402
rect 31208 27338 31260 27344
rect 31220 27130 31248 27338
rect 31208 27124 31260 27130
rect 31208 27066 31260 27072
rect 31404 27062 31432 32846
rect 31496 32774 31524 32846
rect 31680 32842 31708 33050
rect 31668 32836 31720 32842
rect 31668 32778 31720 32784
rect 31484 32768 31536 32774
rect 31484 32710 31536 32716
rect 31760 32768 31812 32774
rect 31760 32710 31812 32716
rect 31772 31822 31800 32710
rect 32140 32434 32168 34002
rect 32864 33924 32916 33930
rect 32864 33866 32916 33872
rect 32588 33856 32640 33862
rect 32588 33798 32640 33804
rect 32312 33516 32364 33522
rect 32312 33458 32364 33464
rect 32220 33312 32272 33318
rect 32220 33254 32272 33260
rect 32232 32978 32260 33254
rect 32220 32972 32272 32978
rect 32220 32914 32272 32920
rect 32324 32842 32352 33458
rect 32600 32910 32628 33798
rect 32876 33658 32904 33866
rect 32864 33652 32916 33658
rect 32864 33594 32916 33600
rect 32864 33516 32916 33522
rect 32864 33458 32916 33464
rect 32588 32904 32640 32910
rect 32588 32846 32640 32852
rect 32312 32836 32364 32842
rect 32312 32778 32364 32784
rect 32772 32836 32824 32842
rect 32772 32778 32824 32784
rect 32128 32428 32180 32434
rect 32128 32370 32180 32376
rect 32784 32366 32812 32778
rect 32496 32360 32548 32366
rect 32496 32302 32548 32308
rect 32772 32360 32824 32366
rect 32772 32302 32824 32308
rect 32220 32224 32272 32230
rect 32220 32166 32272 32172
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31944 31816 31996 31822
rect 31944 31758 31996 31764
rect 32128 31816 32180 31822
rect 32232 31804 32260 32166
rect 32508 32026 32536 32302
rect 32496 32020 32548 32026
rect 32496 31962 32548 31968
rect 32784 31890 32812 32302
rect 32772 31884 32824 31890
rect 32772 31826 32824 31832
rect 32876 31822 32904 33458
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 33048 32496 33100 32502
rect 33048 32438 33100 32444
rect 33060 32026 33088 32438
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 33048 32020 33100 32026
rect 33048 31962 33100 31968
rect 32312 31816 32364 31822
rect 32232 31776 32312 31804
rect 32128 31758 32180 31764
rect 32312 31758 32364 31764
rect 32864 31816 32916 31822
rect 32864 31758 32916 31764
rect 31956 31414 31984 31758
rect 31944 31408 31996 31414
rect 31944 31350 31996 31356
rect 31668 28552 31720 28558
rect 31668 28494 31720 28500
rect 31680 28082 31708 28494
rect 31668 28076 31720 28082
rect 31668 28018 31720 28024
rect 31680 27674 31708 28018
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31392 27056 31444 27062
rect 31392 26998 31444 27004
rect 30380 26988 30432 26994
rect 30380 26930 30432 26936
rect 30748 26988 30800 26994
rect 30748 26930 30800 26936
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 29460 26376 29512 26382
rect 29460 26318 29512 26324
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 29472 26042 29500 26318
rect 29460 26036 29512 26042
rect 29460 25978 29512 25984
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29656 25498 29684 25910
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29564 23322 29592 24142
rect 29644 24064 29696 24070
rect 29644 24006 29696 24012
rect 29656 23798 29684 24006
rect 29644 23792 29696 23798
rect 29644 23734 29696 23740
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29748 23202 29776 25230
rect 29932 23254 29960 26318
rect 32140 25514 32168 31758
rect 32324 31482 32352 31758
rect 32312 31476 32364 31482
rect 32312 31418 32364 31424
rect 32404 31272 32456 31278
rect 32404 31214 32456 31220
rect 32220 31136 32272 31142
rect 32220 31078 32272 31084
rect 32232 30802 32260 31078
rect 32220 30796 32272 30802
rect 32220 30738 32272 30744
rect 32416 30598 32444 31214
rect 32404 30592 32456 30598
rect 32404 30534 32456 30540
rect 32416 28490 32444 30534
rect 32876 30258 32904 31758
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 33232 30660 33284 30666
rect 33232 30602 33284 30608
rect 33244 30326 33272 30602
rect 33232 30320 33284 30326
rect 33232 30262 33284 30268
rect 34886 30288 34942 30297
rect 32864 30252 32916 30258
rect 34886 30223 34942 30232
rect 32864 30194 32916 30200
rect 32876 29646 32904 30194
rect 34900 30190 34928 30223
rect 34336 30184 34388 30190
rect 34336 30126 34388 30132
rect 34796 30184 34848 30190
rect 34796 30126 34848 30132
rect 34888 30184 34940 30190
rect 34888 30126 34940 30132
rect 32864 29640 32916 29646
rect 32864 29582 32916 29588
rect 33138 29200 33194 29209
rect 33138 29135 33194 29144
rect 33152 29102 33180 29135
rect 32680 29096 32732 29102
rect 32680 29038 32732 29044
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 33140 29096 33192 29102
rect 33140 29038 33192 29044
rect 32404 28484 32456 28490
rect 32404 28426 32456 28432
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 32508 27470 32536 28018
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32312 27328 32364 27334
rect 32312 27270 32364 27276
rect 32324 26994 32352 27270
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 32508 25838 32536 27406
rect 32692 27130 32720 29038
rect 32876 28762 32904 29038
rect 34348 28762 34376 30126
rect 34808 29850 34836 30126
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 35348 29640 35400 29646
rect 35348 29582 35400 29588
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 32864 28756 32916 28762
rect 32864 28698 32916 28704
rect 34336 28756 34388 28762
rect 34336 28698 34388 28704
rect 33692 28552 33744 28558
rect 33692 28494 33744 28500
rect 33704 28218 33732 28494
rect 33692 28212 33744 28218
rect 33692 28154 33744 28160
rect 34348 28082 34376 28698
rect 34980 28484 35032 28490
rect 34980 28426 35032 28432
rect 34336 28076 34388 28082
rect 34336 28018 34388 28024
rect 34992 28014 35020 28426
rect 34704 28008 34756 28014
rect 34704 27950 34756 27956
rect 34980 28008 35032 28014
rect 34980 27950 35032 27956
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 32680 27124 32732 27130
rect 32680 27066 32732 27072
rect 32692 26382 32720 27066
rect 33336 27062 33364 27270
rect 34336 27124 34388 27130
rect 34336 27066 34388 27072
rect 33324 27056 33376 27062
rect 33324 26998 33376 27004
rect 33968 27056 34020 27062
rect 33968 26998 34020 27004
rect 33876 26988 33928 26994
rect 33876 26930 33928 26936
rect 33140 26920 33192 26926
rect 33140 26862 33192 26868
rect 33152 26586 33180 26862
rect 33888 26586 33916 26930
rect 33140 26580 33192 26586
rect 33140 26522 33192 26528
rect 33876 26580 33928 26586
rect 33876 26522 33928 26528
rect 33980 26382 34008 26998
rect 32680 26376 32732 26382
rect 32680 26318 32732 26324
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 34348 25974 34376 27066
rect 34612 27056 34664 27062
rect 34532 27016 34612 27044
rect 34428 26376 34480 26382
rect 34428 26318 34480 26324
rect 34532 26330 34560 27016
rect 34612 26998 34664 27004
rect 34612 26852 34664 26858
rect 34612 26794 34664 26800
rect 34624 26450 34652 26794
rect 34612 26444 34664 26450
rect 34612 26386 34664 26392
rect 34716 26330 34744 27950
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35360 26874 35388 29582
rect 35440 28484 35492 28490
rect 35440 28426 35492 28432
rect 35452 28218 35480 28426
rect 35440 28212 35492 28218
rect 35440 28154 35492 28160
rect 35532 28076 35584 28082
rect 35532 28018 35584 28024
rect 35544 27470 35572 28018
rect 35532 27464 35584 27470
rect 35532 27406 35584 27412
rect 35360 26846 35480 26874
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 34808 26466 34836 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34808 26438 34928 26466
rect 35360 26450 35388 26726
rect 34440 26042 34468 26318
rect 34532 26314 34652 26330
rect 34532 26308 34664 26314
rect 34532 26302 34612 26308
rect 34716 26302 34836 26330
rect 34612 26250 34664 26256
rect 34428 26036 34480 26042
rect 34428 25978 34480 25984
rect 34336 25968 34388 25974
rect 34336 25910 34388 25916
rect 34624 25922 34652 26250
rect 34808 26042 34836 26302
rect 34900 26246 34928 26438
rect 35348 26444 35400 26450
rect 35348 26386 35400 26392
rect 34888 26240 34940 26246
rect 34888 26182 34940 26188
rect 34796 26036 34848 26042
rect 34796 25978 34848 25984
rect 34900 25922 34928 26182
rect 34624 25906 34744 25922
rect 34624 25900 34756 25906
rect 34624 25894 34704 25900
rect 34704 25842 34756 25848
rect 34808 25894 34928 25922
rect 32496 25832 32548 25838
rect 32496 25774 32548 25780
rect 34520 25764 34572 25770
rect 34520 25706 34572 25712
rect 32048 25486 32168 25514
rect 34532 25498 34560 25706
rect 34520 25492 34572 25498
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31484 24812 31536 24818
rect 31484 24754 31536 24760
rect 30748 24608 30800 24614
rect 30748 24550 30800 24556
rect 30760 24274 30788 24550
rect 30748 24268 30800 24274
rect 30748 24210 30800 24216
rect 30472 24200 30524 24206
rect 30472 24142 30524 24148
rect 30484 23866 30512 24142
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30840 23656 30892 23662
rect 30840 23598 30892 23604
rect 29656 23174 29776 23202
rect 29920 23248 29972 23254
rect 29920 23190 29972 23196
rect 29656 23118 29684 23174
rect 30852 23118 30880 23598
rect 31312 23594 31340 24754
rect 31496 23594 31524 24754
rect 31576 24744 31628 24750
rect 31576 24686 31628 24692
rect 31588 23730 31616 24686
rect 31760 24132 31812 24138
rect 31760 24074 31812 24080
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31300 23588 31352 23594
rect 31300 23530 31352 23536
rect 31484 23588 31536 23594
rect 31484 23530 31536 23536
rect 29644 23112 29696 23118
rect 29644 23054 29696 23060
rect 30840 23112 30892 23118
rect 30840 23054 30892 23060
rect 30932 22976 30984 22982
rect 30932 22918 30984 22924
rect 30944 22098 30972 22918
rect 31496 22574 31524 23530
rect 31772 23322 31800 24074
rect 31760 23316 31812 23322
rect 31760 23258 31812 23264
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31484 22568 31536 22574
rect 31484 22510 31536 22516
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31220 22234 31248 22374
rect 31208 22228 31260 22234
rect 31208 22170 31260 22176
rect 30932 22092 30984 22098
rect 30932 22034 30984 22040
rect 31760 22094 31812 22098
rect 31864 22094 31892 22578
rect 31760 22092 31892 22094
rect 31812 22066 31892 22092
rect 32048 22094 32076 25486
rect 34520 25434 34572 25440
rect 33508 24812 33560 24818
rect 33508 24754 33560 24760
rect 33232 24744 33284 24750
rect 33232 24686 33284 24692
rect 33244 24342 33272 24686
rect 33232 24336 33284 24342
rect 33232 24278 33284 24284
rect 32956 24200 33008 24206
rect 33008 24148 33088 24154
rect 32956 24142 33088 24148
rect 32680 24132 32732 24138
rect 32680 24074 32732 24080
rect 32772 24132 32824 24138
rect 32968 24126 33088 24142
rect 32772 24074 32824 24080
rect 32128 24064 32180 24070
rect 32128 24006 32180 24012
rect 32140 23798 32168 24006
rect 32692 23798 32720 24074
rect 32128 23792 32180 23798
rect 32128 23734 32180 23740
rect 32680 23792 32732 23798
rect 32680 23734 32732 23740
rect 32784 23526 32812 24074
rect 33060 23730 33088 24126
rect 33520 23866 33548 24754
rect 33968 24608 34020 24614
rect 33968 24550 34020 24556
rect 33508 23860 33560 23866
rect 33508 23802 33560 23808
rect 33980 23798 34008 24550
rect 34532 24206 34560 25434
rect 34612 24744 34664 24750
rect 34716 24732 34744 25842
rect 34808 25838 34836 25894
rect 34796 25832 34848 25838
rect 34796 25774 34848 25780
rect 34808 24818 34836 25774
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34796 24812 34848 24818
rect 34796 24754 34848 24760
rect 34664 24704 34744 24732
rect 35452 24698 35480 26846
rect 35544 25906 35572 27406
rect 35532 25900 35584 25906
rect 35532 25842 35584 25848
rect 34612 24686 34664 24692
rect 35360 24670 35480 24698
rect 35532 24744 35584 24750
rect 35532 24686 35584 24692
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 35360 24154 35388 24670
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 35452 24274 35480 24550
rect 35440 24268 35492 24274
rect 35440 24210 35492 24216
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 34072 23798 34100 24006
rect 33968 23792 34020 23798
rect 33968 23734 34020 23740
rect 34060 23792 34112 23798
rect 34060 23734 34112 23740
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 32140 22642 32168 22986
rect 32864 22772 32916 22778
rect 32864 22714 32916 22720
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32220 22432 32272 22438
rect 32220 22374 32272 22380
rect 32048 22066 32168 22094
rect 31760 22034 31812 22040
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 30196 21888 30248 21894
rect 30196 21830 30248 21836
rect 29748 21622 29776 21830
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 30208 21486 30236 21830
rect 30196 21480 30248 21486
rect 30196 21422 30248 21428
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 30300 21010 30328 21354
rect 31772 21010 31800 22034
rect 30288 21004 30340 21010
rect 30288 20946 30340 20952
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29840 20534 29868 20742
rect 30300 20602 30328 20946
rect 31392 20868 31444 20874
rect 31392 20810 31444 20816
rect 31404 20602 31432 20810
rect 30288 20596 30340 20602
rect 30288 20538 30340 20544
rect 31392 20596 31444 20602
rect 31392 20538 31444 20544
rect 29828 20528 29880 20534
rect 29828 20470 29880 20476
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31312 20262 31340 20402
rect 31300 20256 31352 20262
rect 31300 20198 31352 20204
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29472 17134 29500 18226
rect 29736 18080 29788 18086
rect 29736 18022 29788 18028
rect 29748 17678 29776 18022
rect 29840 17746 29868 18906
rect 30300 18766 30328 18906
rect 31392 18828 31444 18834
rect 31392 18770 31444 18776
rect 30288 18760 30340 18766
rect 30288 18702 30340 18708
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 30656 18148 30708 18154
rect 30656 18090 30708 18096
rect 30668 17746 30696 18090
rect 31220 17882 31248 18158
rect 31208 17876 31260 17882
rect 31208 17818 31260 17824
rect 29828 17740 29880 17746
rect 29828 17682 29880 17688
rect 30656 17740 30708 17746
rect 30656 17682 30708 17688
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31128 17542 31156 17614
rect 31116 17536 31168 17542
rect 31116 17478 31168 17484
rect 29460 17128 29512 17134
rect 29460 17070 29512 17076
rect 30656 17128 30708 17134
rect 30656 17070 30708 17076
rect 29472 16998 29500 17070
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29828 16992 29880 16998
rect 29828 16934 29880 16940
rect 30380 16992 30432 16998
rect 30380 16934 30432 16940
rect 29840 16590 29868 16934
rect 29644 16584 29696 16590
rect 29644 16526 29696 16532
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 29656 16250 29684 16526
rect 29644 16244 29696 16250
rect 29644 16186 29696 16192
rect 30392 16114 30420 16934
rect 30668 16658 30696 17070
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30564 15904 30616 15910
rect 30564 15846 30616 15852
rect 30576 15570 30604 15846
rect 30564 15564 30616 15570
rect 30564 15506 30616 15512
rect 30656 15564 30708 15570
rect 30656 15506 30708 15512
rect 29368 12640 29420 12646
rect 29368 12582 29420 12588
rect 30668 2774 30696 15506
rect 31128 4690 31156 17478
rect 31116 4684 31168 4690
rect 31116 4626 31168 4632
rect 31404 4146 31432 18770
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 31404 3670 31432 4082
rect 31392 3664 31444 3670
rect 31392 3606 31444 3612
rect 30576 2746 30696 2774
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29276 1964 29328 1970
rect 29276 1906 29328 1912
rect 29656 800 29684 2382
rect 22756 734 23060 762
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30576 762 30604 2746
rect 32140 2582 32168 22066
rect 32232 21962 32260 22374
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 32220 21956 32272 21962
rect 32220 21898 32272 21904
rect 32508 21554 32536 21966
rect 32496 21548 32548 21554
rect 32496 21490 32548 21496
rect 32220 20324 32272 20330
rect 32220 20266 32272 20272
rect 32232 19446 32260 20266
rect 32508 20058 32536 21490
rect 32772 21480 32824 21486
rect 32772 21422 32824 21428
rect 32784 21350 32812 21422
rect 32772 21344 32824 21350
rect 32772 21286 32824 21292
rect 32496 20052 32548 20058
rect 32496 19994 32548 20000
rect 32404 19848 32456 19854
rect 32404 19790 32456 19796
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 32416 18970 32444 19790
rect 32496 19304 32548 19310
rect 32496 19246 32548 19252
rect 32404 18964 32456 18970
rect 32404 18906 32456 18912
rect 32508 18902 32536 19246
rect 32588 18964 32640 18970
rect 32588 18906 32640 18912
rect 32496 18896 32548 18902
rect 32496 18838 32548 18844
rect 32496 16516 32548 16522
rect 32496 16458 32548 16464
rect 32508 16250 32536 16458
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32600 6914 32628 18906
rect 32784 16114 32812 21286
rect 32876 18154 32904 22714
rect 32956 22432 33008 22438
rect 32956 22374 33008 22380
rect 32968 22030 32996 22374
rect 33060 22098 33088 23666
rect 34532 23662 34560 24142
rect 33692 23656 33744 23662
rect 33692 23598 33744 23604
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 33704 23322 33732 23598
rect 33784 23520 33836 23526
rect 33784 23462 33836 23468
rect 33692 23316 33744 23322
rect 33692 23258 33744 23264
rect 33692 22432 33744 22438
rect 33692 22374 33744 22380
rect 33048 22092 33100 22098
rect 33048 22034 33100 22040
rect 32956 22024 33008 22030
rect 32956 21966 33008 21972
rect 33416 21072 33468 21078
rect 33414 21040 33416 21049
rect 33468 21040 33470 21049
rect 33414 20975 33470 20984
rect 33704 20942 33732 22374
rect 33796 21962 33824 23462
rect 34808 23322 34836 24142
rect 35360 24126 35480 24154
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34796 23316 34848 23322
rect 34796 23258 34848 23264
rect 33876 23044 33928 23050
rect 33876 22986 33928 22992
rect 33888 22642 33916 22986
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 33876 22500 33928 22506
rect 33876 22442 33928 22448
rect 33784 21956 33836 21962
rect 33784 21898 33836 21904
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 33048 20868 33100 20874
rect 33048 20810 33100 20816
rect 32864 18148 32916 18154
rect 32864 18090 32916 18096
rect 32772 16108 32824 16114
rect 32772 16050 32824 16056
rect 33060 6914 33088 20810
rect 33704 20466 33732 20878
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 33508 19712 33560 19718
rect 33508 19654 33560 19660
rect 33244 19310 33272 19654
rect 33520 19446 33548 19654
rect 33324 19440 33376 19446
rect 33324 19382 33376 19388
rect 33508 19440 33560 19446
rect 33508 19382 33560 19388
rect 33232 19304 33284 19310
rect 33232 19246 33284 19252
rect 33244 18902 33272 19246
rect 33336 18970 33364 19382
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 33232 18896 33284 18902
rect 33232 18838 33284 18844
rect 33796 17762 33824 21898
rect 33888 20534 33916 22442
rect 34796 22432 34848 22438
rect 34796 22374 34848 22380
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 34716 20534 34744 21966
rect 34808 20856 34836 22374
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35360 22234 35388 22578
rect 35348 22228 35400 22234
rect 35348 22170 35400 22176
rect 35346 21584 35402 21593
rect 35346 21519 35348 21528
rect 35400 21519 35402 21528
rect 35348 21490 35400 21496
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35452 21078 35480 24126
rect 35544 23866 35572 24686
rect 35532 23860 35584 23866
rect 35532 23802 35584 23808
rect 35636 22234 35664 35866
rect 35624 22228 35676 22234
rect 35624 22170 35676 22176
rect 35440 21072 35492 21078
rect 35440 21014 35492 21020
rect 35072 20868 35124 20874
rect 34808 20828 35072 20856
rect 35072 20810 35124 20816
rect 33876 20528 33928 20534
rect 33876 20470 33928 20476
rect 34704 20528 34756 20534
rect 34704 20470 34756 20476
rect 35624 20528 35676 20534
rect 35624 20470 35676 20476
rect 35440 20392 35492 20398
rect 35440 20334 35492 20340
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35452 19854 35480 20334
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35072 18828 35124 18834
rect 35072 18770 35124 18776
rect 35084 18290 35112 18770
rect 35452 18698 35480 19790
rect 35440 18692 35492 18698
rect 35440 18634 35492 18640
rect 35072 18284 35124 18290
rect 35072 18226 35124 18232
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33888 17882 33916 18158
rect 34520 18148 34572 18154
rect 34520 18090 34572 18096
rect 33876 17876 33928 17882
rect 33876 17818 33928 17824
rect 33796 17734 33916 17762
rect 33888 14346 33916 17734
rect 34532 17678 34560 18090
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 35072 17808 35124 17814
rect 35072 17750 35124 17756
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 35084 17270 35112 17750
rect 35360 17678 35388 18022
rect 35452 17678 35480 18226
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 35440 17672 35492 17678
rect 35440 17614 35492 17620
rect 35072 17264 35124 17270
rect 35072 17206 35124 17212
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 33876 14340 33928 14346
rect 33876 14282 33928 14288
rect 32508 6886 32628 6914
rect 32784 6886 33088 6914
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 30760 870 30972 898
rect 30760 762 30788 870
rect 30944 800 30972 870
rect 32232 800 32260 2790
rect 32508 2514 32536 6886
rect 32784 2990 32812 6886
rect 33888 3602 33916 14282
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 32864 3596 32916 3602
rect 32864 3538 32916 3544
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 32876 3058 32904 3538
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 33060 3126 33088 3334
rect 33048 3120 33100 3126
rect 33048 3062 33100 3068
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 32772 2984 32824 2990
rect 32772 2926 32824 2932
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 32496 2508 32548 2514
rect 32496 2450 32548 2456
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35544 2650 35572 3674
rect 35636 2650 35664 20470
rect 35728 18426 35756 43182
rect 36176 28620 36228 28626
rect 36176 28562 36228 28568
rect 35808 27124 35860 27130
rect 35808 27066 35860 27072
rect 35820 26466 35848 27066
rect 35820 26450 36032 26466
rect 35820 26444 36044 26450
rect 35820 26438 35992 26444
rect 35820 25974 35848 26438
rect 35992 26386 36044 26392
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 36004 26042 36032 26250
rect 35992 26036 36044 26042
rect 35992 25978 36044 25984
rect 35808 25968 35860 25974
rect 35808 25910 35860 25916
rect 35820 24274 35848 25910
rect 36084 25356 36136 25362
rect 36084 25298 36136 25304
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35808 24268 35860 24274
rect 35808 24210 35860 24216
rect 35912 22506 35940 25230
rect 35992 24132 36044 24138
rect 35992 24074 36044 24080
rect 36004 23866 36032 24074
rect 36096 24070 36124 25298
rect 36188 25294 36216 28562
rect 36912 26376 36964 26382
rect 36912 26318 36964 26324
rect 36176 25288 36228 25294
rect 36176 25230 36228 25236
rect 36924 24818 36952 26318
rect 37648 26308 37700 26314
rect 37648 26250 37700 26256
rect 37660 25498 37688 26250
rect 37648 25492 37700 25498
rect 37648 25434 37700 25440
rect 37188 25424 37240 25430
rect 37188 25366 37240 25372
rect 37200 25294 37228 25366
rect 37188 25288 37240 25294
rect 37188 25230 37240 25236
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 37464 25152 37516 25158
rect 37464 25094 37516 25100
rect 36912 24812 36964 24818
rect 36912 24754 36964 24760
rect 36924 24342 36952 24754
rect 37476 24750 37504 25094
rect 37464 24744 37516 24750
rect 37464 24686 37516 24692
rect 37844 24614 37872 25230
rect 37832 24608 37884 24614
rect 37832 24550 37884 24556
rect 36912 24336 36964 24342
rect 36912 24278 36964 24284
rect 37648 24132 37700 24138
rect 37648 24074 37700 24080
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 37660 23866 37688 24074
rect 35992 23860 36044 23866
rect 35992 23802 36044 23808
rect 37648 23860 37700 23866
rect 37648 23802 37700 23808
rect 37464 23724 37516 23730
rect 37464 23666 37516 23672
rect 37280 22976 37332 22982
rect 37280 22918 37332 22924
rect 37292 22642 37320 22918
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 35900 22500 35952 22506
rect 35900 22442 35952 22448
rect 36636 21956 36688 21962
rect 36636 21898 36688 21904
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 35992 20868 36044 20874
rect 35992 20810 36044 20816
rect 36004 20534 36032 20810
rect 35992 20528 36044 20534
rect 35992 20470 36044 20476
rect 36372 19990 36400 21830
rect 36648 21690 36676 21898
rect 37188 21888 37240 21894
rect 37292 21842 37320 22578
rect 37240 21836 37320 21842
rect 37188 21830 37320 21836
rect 37200 21814 37320 21830
rect 36636 21684 36688 21690
rect 36636 21626 36688 21632
rect 37292 21622 37320 21814
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 37292 20942 37320 21558
rect 37280 20936 37332 20942
rect 37280 20878 37332 20884
rect 37476 20262 37504 23666
rect 37844 23526 37872 24550
rect 37832 23520 37884 23526
rect 37832 23462 37884 23468
rect 38108 23316 38160 23322
rect 38108 23258 38160 23264
rect 38120 22710 38148 23258
rect 38108 22704 38160 22710
rect 38108 22646 38160 22652
rect 38014 21040 38070 21049
rect 38014 20975 38070 20984
rect 38028 20942 38056 20975
rect 38016 20936 38068 20942
rect 38016 20878 38068 20884
rect 37464 20256 37516 20262
rect 37464 20198 37516 20204
rect 36360 19984 36412 19990
rect 36360 19926 36412 19932
rect 36372 19786 36400 19926
rect 36360 19780 36412 19786
rect 36360 19722 36412 19728
rect 38028 19334 38056 20878
rect 37936 19306 38056 19334
rect 36544 18692 36596 18698
rect 36544 18634 36596 18640
rect 35716 18420 35768 18426
rect 35716 18362 35768 18368
rect 35728 17882 35756 18362
rect 36556 18222 36584 18634
rect 36544 18216 36596 18222
rect 36544 18158 36596 18164
rect 35716 17876 35768 17882
rect 35716 17818 35768 17824
rect 35728 17610 35756 17818
rect 35716 17604 35768 17610
rect 35716 17546 35768 17552
rect 36556 17338 36584 18158
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 36556 17134 36584 17274
rect 36544 17128 36596 17134
rect 36544 17070 36596 17076
rect 37464 5296 37516 5302
rect 37464 5238 37516 5244
rect 37372 4208 37424 4214
rect 37372 4150 37424 4156
rect 36728 4140 36780 4146
rect 36728 4082 36780 4088
rect 36740 3194 36768 4082
rect 37384 3738 37412 4150
rect 37476 3942 37504 5238
rect 37556 4208 37608 4214
rect 37556 4150 37608 4156
rect 37568 3942 37596 4150
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37556 3936 37608 3942
rect 37556 3878 37608 3884
rect 37372 3732 37424 3738
rect 37372 3674 37424 3680
rect 36728 3188 36780 3194
rect 36728 3130 36780 3136
rect 37384 2990 37412 3674
rect 37568 3058 37596 3878
rect 37936 3534 37964 19306
rect 38120 18290 38148 22646
rect 38212 21418 38240 45290
rect 38580 31754 38608 45526
rect 38660 45484 38712 45490
rect 38660 45426 38712 45432
rect 38672 43790 38700 45426
rect 40052 44334 40080 45526
rect 38752 44328 38804 44334
rect 38752 44270 38804 44276
rect 40040 44328 40092 44334
rect 40040 44270 40092 44276
rect 38764 43994 38792 44270
rect 38752 43988 38804 43994
rect 38752 43930 38804 43936
rect 38660 43784 38712 43790
rect 38660 43726 38712 43732
rect 38672 38554 38700 43726
rect 38936 40928 38988 40934
rect 38936 40870 38988 40876
rect 38660 38548 38712 38554
rect 38660 38490 38712 38496
rect 38488 31726 38608 31754
rect 38488 24750 38516 31726
rect 38476 24744 38528 24750
rect 38476 24686 38528 24692
rect 38672 23322 38700 38490
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38384 23180 38436 23186
rect 38384 23122 38436 23128
rect 38200 21412 38252 21418
rect 38200 21354 38252 21360
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 38120 6914 38148 18226
rect 38028 6886 38148 6914
rect 38028 4078 38056 6886
rect 38396 5166 38424 23122
rect 38948 23118 38976 40870
rect 40236 31278 40264 46990
rect 40224 31272 40276 31278
rect 40224 31214 40276 31220
rect 40132 25220 40184 25226
rect 40132 25162 40184 25168
rect 40144 24954 40172 25162
rect 40132 24948 40184 24954
rect 40132 24890 40184 24896
rect 40040 24812 40092 24818
rect 40040 24754 40092 24760
rect 40052 24614 40080 24754
rect 40040 24608 40092 24614
rect 40040 24550 40092 24556
rect 40316 24268 40368 24274
rect 40316 24210 40368 24216
rect 39856 24200 39908 24206
rect 40328 24177 40356 24210
rect 39856 24142 39908 24148
rect 40314 24168 40370 24177
rect 39304 24132 39356 24138
rect 39304 24074 39356 24080
rect 39212 23724 39264 23730
rect 39212 23666 39264 23672
rect 38936 23112 38988 23118
rect 38936 23054 38988 23060
rect 38936 21616 38988 21622
rect 38936 21558 38988 21564
rect 38948 21350 38976 21558
rect 38936 21344 38988 21350
rect 38936 21286 38988 21292
rect 38948 21010 38976 21286
rect 38936 21004 38988 21010
rect 38936 20946 38988 20952
rect 38948 9586 38976 20946
rect 39224 17542 39252 23666
rect 39212 17536 39264 17542
rect 39212 17478 39264 17484
rect 38936 9580 38988 9586
rect 38936 9522 38988 9528
rect 38476 5908 38528 5914
rect 38476 5850 38528 5856
rect 38384 5160 38436 5166
rect 38384 5102 38436 5108
rect 38396 4214 38424 5102
rect 38384 4208 38436 4214
rect 38384 4150 38436 4156
rect 38016 4072 38068 4078
rect 38016 4014 38068 4020
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 37556 3052 37608 3058
rect 37556 2994 37608 3000
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 35624 2644 35676 2650
rect 35624 2586 35676 2592
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 36096 800 36124 2314
rect 36372 2038 36400 2790
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 36360 2032 36412 2038
rect 36360 1974 36412 1980
rect 38028 800 38056 2382
rect 38488 2310 38516 5850
rect 39120 5024 39172 5030
rect 39120 4966 39172 4972
rect 39132 4622 39160 4966
rect 39120 4616 39172 4622
rect 39120 4558 39172 4564
rect 39120 4140 39172 4146
rect 39120 4082 39172 4088
rect 38568 3732 38620 3738
rect 38568 3674 38620 3680
rect 38580 3534 38608 3674
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 39132 3194 39160 4082
rect 39316 3670 39344 24074
rect 39868 23186 39896 24142
rect 40040 24132 40092 24138
rect 40314 24103 40370 24112
rect 40040 24074 40092 24080
rect 40052 23866 40080 24074
rect 40040 23860 40092 23866
rect 40040 23802 40092 23808
rect 39856 23180 39908 23186
rect 39856 23122 39908 23128
rect 39580 22976 39632 22982
rect 39580 22918 39632 22924
rect 39592 22574 39620 22918
rect 39868 22778 39896 23122
rect 40132 23044 40184 23050
rect 40132 22986 40184 22992
rect 39856 22772 39908 22778
rect 39856 22714 39908 22720
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 39580 22568 39632 22574
rect 39580 22510 39632 22516
rect 40052 22030 40080 22578
rect 40144 22234 40172 22986
rect 40224 22568 40276 22574
rect 40224 22510 40276 22516
rect 40132 22228 40184 22234
rect 40132 22170 40184 22176
rect 40236 22098 40264 22510
rect 40604 22438 40632 47194
rect 41248 46918 41276 49200
rect 41236 46912 41288 46918
rect 41236 46854 41288 46860
rect 41788 46912 41840 46918
rect 41788 46854 41840 46860
rect 41328 46368 41380 46374
rect 41328 46310 41380 46316
rect 41340 46034 41368 46310
rect 41328 46028 41380 46034
rect 41328 45970 41380 45976
rect 41512 45892 41564 45898
rect 41512 45834 41564 45840
rect 41524 45626 41552 45834
rect 41512 45620 41564 45626
rect 41512 45562 41564 45568
rect 41328 45484 41380 45490
rect 41328 45426 41380 45432
rect 41340 44470 41368 45426
rect 41328 44464 41380 44470
rect 41328 44406 41380 44412
rect 41800 25362 41828 46854
rect 41892 46034 41920 49200
rect 42536 46442 42564 49200
rect 43180 47122 43208 49200
rect 43168 47116 43220 47122
rect 43168 47058 43220 47064
rect 43168 46980 43220 46986
rect 43168 46922 43220 46928
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 41880 46028 41932 46034
rect 41880 45970 41932 45976
rect 42628 45626 42656 46446
rect 42984 46096 43036 46102
rect 42984 46038 43036 46044
rect 42616 45620 42668 45626
rect 42616 45562 42668 45568
rect 42996 38418 43024 46038
rect 43180 45558 43208 46922
rect 43824 45966 43852 49200
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 44088 45824 44140 45830
rect 44088 45766 44140 45772
rect 43168 45552 43220 45558
rect 43168 45494 43220 45500
rect 43076 45484 43128 45490
rect 43076 45426 43128 45432
rect 43088 45014 43116 45426
rect 43904 45280 43956 45286
rect 43904 45222 43956 45228
rect 43076 45008 43128 45014
rect 43076 44950 43128 44956
rect 42984 38412 43036 38418
rect 42984 38354 43036 38360
rect 42996 37398 43024 38354
rect 42984 37392 43036 37398
rect 42984 37334 43036 37340
rect 43628 37256 43680 37262
rect 43628 37198 43680 37204
rect 42708 31952 42760 31958
rect 42708 31894 42760 31900
rect 41788 25356 41840 25362
rect 41788 25298 41840 25304
rect 42340 23180 42392 23186
rect 42340 23122 42392 23128
rect 41788 23044 41840 23050
rect 41788 22986 41840 22992
rect 41880 23044 41932 23050
rect 41880 22986 41932 22992
rect 41800 22778 41828 22986
rect 41788 22772 41840 22778
rect 41788 22714 41840 22720
rect 41800 22522 41828 22714
rect 41892 22642 41920 22986
rect 41880 22636 41932 22642
rect 41880 22578 41932 22584
rect 42352 22574 42380 23122
rect 42340 22568 42392 22574
rect 41800 22494 41920 22522
rect 42340 22510 42392 22516
rect 40592 22432 40644 22438
rect 40592 22374 40644 22380
rect 40868 22432 40920 22438
rect 40868 22374 40920 22380
rect 41788 22432 41840 22438
rect 41788 22374 41840 22380
rect 40224 22092 40276 22098
rect 40224 22034 40276 22040
rect 40604 22030 40632 22374
rect 40880 22030 40908 22374
rect 41800 22030 41828 22374
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 40592 22024 40644 22030
rect 40592 21966 40644 21972
rect 40868 22024 40920 22030
rect 40868 21966 40920 21972
rect 41788 22024 41840 22030
rect 41788 21966 41840 21972
rect 40052 21690 40080 21966
rect 40224 21956 40276 21962
rect 40224 21898 40276 21904
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 40040 4548 40092 4554
rect 40040 4490 40092 4496
rect 40052 4282 40080 4490
rect 40040 4276 40092 4282
rect 40040 4218 40092 4224
rect 40236 4214 40264 21898
rect 41892 17338 41920 22494
rect 42248 20936 42300 20942
rect 42248 20878 42300 20884
rect 42260 20602 42288 20878
rect 42248 20596 42300 20602
rect 42248 20538 42300 20544
rect 41880 17332 41932 17338
rect 41880 17274 41932 17280
rect 41892 6914 41920 17274
rect 41708 6886 41920 6914
rect 41420 6724 41472 6730
rect 41420 6666 41472 6672
rect 41432 6458 41460 6666
rect 41420 6452 41472 6458
rect 41420 6394 41472 6400
rect 41328 6316 41380 6322
rect 41328 6258 41380 6264
rect 41340 5914 41368 6258
rect 41604 6248 41656 6254
rect 41604 6190 41656 6196
rect 41328 5908 41380 5914
rect 41328 5850 41380 5856
rect 41328 5228 41380 5234
rect 41328 5170 41380 5176
rect 40224 4208 40276 4214
rect 40224 4150 40276 4156
rect 39856 4140 39908 4146
rect 39856 4082 39908 4088
rect 39304 3664 39356 3670
rect 39304 3606 39356 3612
rect 39120 3188 39172 3194
rect 39120 3130 39172 3136
rect 39868 2990 39896 4082
rect 40040 3188 40092 3194
rect 40040 3130 40092 3136
rect 39856 2984 39908 2990
rect 39856 2926 39908 2932
rect 39868 2854 39896 2926
rect 40052 2922 40080 3130
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 40040 2916 40092 2922
rect 40040 2858 40092 2864
rect 39856 2848 39908 2854
rect 40144 2802 40172 2994
rect 39856 2790 39908 2796
rect 39868 2446 39896 2790
rect 39960 2774 40172 2802
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 38476 2304 38528 2310
rect 38476 2246 38528 2252
rect 39316 800 39344 2314
rect 39960 800 39988 2774
rect 40236 2650 40264 4150
rect 41340 4146 41368 5170
rect 41328 4140 41380 4146
rect 41328 4082 41380 4088
rect 40788 3590 41184 3618
rect 40408 3528 40460 3534
rect 40408 3470 40460 3476
rect 40420 2650 40448 3470
rect 40788 3466 40816 3590
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 40776 3460 40828 3466
rect 40776 3402 40828 3408
rect 40880 3194 40908 3470
rect 41156 3398 41184 3590
rect 41144 3392 41196 3398
rect 41144 3334 41196 3340
rect 40684 3188 40736 3194
rect 40684 3130 40736 3136
rect 40868 3188 40920 3194
rect 40868 3130 40920 3136
rect 40696 2990 40724 3130
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40224 2644 40276 2650
rect 40224 2586 40276 2592
rect 40408 2644 40460 2650
rect 40408 2586 40460 2592
rect 40604 2514 40632 2926
rect 41616 2922 41644 6190
rect 41708 4554 41736 6886
rect 42352 6866 42380 22510
rect 42720 21554 42748 31894
rect 42800 28212 42852 28218
rect 42800 28154 42852 28160
rect 42812 26450 42840 28154
rect 42800 26444 42852 26450
rect 42800 26386 42852 26392
rect 43640 26234 43668 37198
rect 43916 29578 43944 45222
rect 44100 35601 44128 45766
rect 44180 45554 44232 45558
rect 44468 45554 44496 49200
rect 45112 45626 45140 49200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 45620 45152 45626
rect 45100 45562 45152 45568
rect 44180 45552 44496 45554
rect 44232 45526 44496 45552
rect 44180 45494 44232 45500
rect 44456 45416 44508 45422
rect 44456 45358 44508 45364
rect 45100 45416 45152 45422
rect 45100 45358 45152 45364
rect 44468 45082 44496 45358
rect 45112 45082 45140 45358
rect 44456 45076 44508 45082
rect 44456 45018 44508 45024
rect 45100 45076 45152 45082
rect 45100 45018 45152 45024
rect 45204 44946 45232 46990
rect 45376 46980 45428 46986
rect 45376 46922 45428 46928
rect 45192 44940 45244 44946
rect 45192 44882 45244 44888
rect 45008 44872 45060 44878
rect 45008 44814 45060 44820
rect 44272 38956 44324 38962
rect 44272 38898 44324 38904
rect 44180 38752 44232 38758
rect 44180 38694 44232 38700
rect 44192 37262 44220 38694
rect 44284 38350 44312 38898
rect 44732 38888 44784 38894
rect 44732 38830 44784 38836
rect 44272 38344 44324 38350
rect 44272 38286 44324 38292
rect 44284 37874 44312 38286
rect 44272 37868 44324 37874
rect 44272 37810 44324 37816
rect 44284 37466 44312 37810
rect 44272 37460 44324 37466
rect 44272 37402 44324 37408
rect 44180 37256 44232 37262
rect 44180 37198 44232 37204
rect 44086 35592 44142 35601
rect 44086 35527 44142 35536
rect 44180 33312 44232 33318
rect 44180 33254 44232 33260
rect 44192 32570 44220 33254
rect 44180 32564 44232 32570
rect 44180 32506 44232 32512
rect 43904 29572 43956 29578
rect 43904 29514 43956 29520
rect 43272 26206 43668 26234
rect 42984 23724 43036 23730
rect 42984 23666 43036 23672
rect 42800 23520 42852 23526
rect 42800 23462 42852 23468
rect 42812 22642 42840 23462
rect 42996 23322 43024 23666
rect 42984 23316 43036 23322
rect 42984 23258 43036 23264
rect 43272 22982 43300 26206
rect 43444 23656 43496 23662
rect 43444 23598 43496 23604
rect 43456 22982 43484 23598
rect 43260 22976 43312 22982
rect 43260 22918 43312 22924
rect 43444 22976 43496 22982
rect 43444 22918 43496 22924
rect 42800 22636 42852 22642
rect 42800 22578 42852 22584
rect 42892 22568 42944 22574
rect 42892 22510 42944 22516
rect 42904 22094 42932 22510
rect 42812 22066 42932 22094
rect 42812 22030 42840 22066
rect 42800 22024 42852 22030
rect 42800 21966 42852 21972
rect 42708 21548 42760 21554
rect 42708 21490 42760 21496
rect 42616 21480 42668 21486
rect 42616 21422 42668 21428
rect 42628 20466 42656 21422
rect 42616 20460 42668 20466
rect 42616 20402 42668 20408
rect 42524 20324 42576 20330
rect 42524 20266 42576 20272
rect 42536 19990 42564 20266
rect 42524 19984 42576 19990
rect 42524 19926 42576 19932
rect 42628 19786 42656 20402
rect 42720 20398 42748 21490
rect 42812 21146 42840 21966
rect 43456 21962 43484 22918
rect 44744 22094 44772 38830
rect 45020 38418 45048 44814
rect 45388 44538 45416 46922
rect 45468 46436 45520 46442
rect 45468 46378 45520 46384
rect 45376 44532 45428 44538
rect 45376 44474 45428 44480
rect 45480 43314 45508 46378
rect 45756 45966 45784 49200
rect 46400 47410 46428 49200
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46400 47382 46796 47410
rect 46386 47016 46442 47025
rect 46386 46951 46442 46960
rect 45836 46028 45888 46034
rect 45836 45970 45888 45976
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45652 45552 45704 45558
rect 45848 45554 45876 45970
rect 45652 45494 45704 45500
rect 45756 45526 45876 45554
rect 45664 44878 45692 45494
rect 45652 44872 45704 44878
rect 45652 44814 45704 44820
rect 45560 44464 45612 44470
rect 45560 44406 45612 44412
rect 45468 43308 45520 43314
rect 45468 43250 45520 43256
rect 45008 38412 45060 38418
rect 45008 38354 45060 38360
rect 45020 26234 45048 38354
rect 45572 38282 45600 44406
rect 45756 44402 45784 45526
rect 46296 44872 46348 44878
rect 46296 44814 46348 44820
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 46204 44396 46256 44402
rect 46204 44338 46256 44344
rect 45928 44192 45980 44198
rect 45928 44134 45980 44140
rect 45940 43858 45968 44134
rect 45928 43852 45980 43858
rect 45928 43794 45980 43800
rect 45836 38956 45888 38962
rect 45836 38898 45888 38904
rect 45468 38276 45520 38282
rect 45468 38218 45520 38224
rect 45560 38276 45612 38282
rect 45560 38218 45612 38224
rect 45480 26234 45508 38218
rect 45560 37800 45612 37806
rect 45560 37742 45612 37748
rect 45572 36378 45600 37742
rect 45560 36372 45612 36378
rect 45560 36314 45612 36320
rect 45572 32434 45600 36314
rect 45560 32428 45612 32434
rect 45560 32370 45612 32376
rect 45650 26616 45706 26625
rect 45650 26551 45706 26560
rect 44928 26206 45048 26234
rect 45388 26206 45508 26234
rect 44928 25906 44956 26206
rect 44916 25900 44968 25906
rect 44916 25842 44968 25848
rect 44824 24880 44876 24886
rect 44824 24822 44876 24828
rect 44652 22066 44772 22094
rect 44456 22024 44508 22030
rect 44456 21966 44508 21972
rect 43444 21956 43496 21962
rect 43444 21898 43496 21904
rect 43536 21616 43588 21622
rect 43536 21558 43588 21564
rect 43168 21344 43220 21350
rect 43168 21286 43220 21292
rect 42800 21140 42852 21146
rect 42800 21082 42852 21088
rect 43180 20942 43208 21286
rect 42892 20936 42944 20942
rect 43168 20936 43220 20942
rect 42944 20884 43024 20890
rect 42892 20878 43024 20884
rect 43168 20878 43220 20884
rect 42904 20862 43024 20878
rect 43548 20874 43576 21558
rect 43812 21548 43864 21554
rect 43812 21490 43864 21496
rect 43996 21548 44048 21554
rect 43996 21490 44048 21496
rect 43720 20936 43772 20942
rect 43720 20878 43772 20884
rect 42800 20800 42852 20806
rect 42800 20742 42852 20748
rect 42892 20800 42944 20806
rect 42892 20742 42944 20748
rect 42708 20392 42760 20398
rect 42708 20334 42760 20340
rect 42720 19854 42748 20334
rect 42812 19854 42840 20742
rect 42904 20398 42932 20742
rect 42996 20602 43024 20862
rect 43536 20868 43588 20874
rect 43536 20810 43588 20816
rect 43168 20800 43220 20806
rect 43168 20742 43220 20748
rect 42984 20596 43036 20602
rect 42984 20538 43036 20544
rect 42892 20392 42944 20398
rect 42892 20334 42944 20340
rect 42892 20256 42944 20262
rect 42892 20198 42944 20204
rect 42708 19848 42760 19854
rect 42708 19790 42760 19796
rect 42800 19848 42852 19854
rect 42800 19790 42852 19796
rect 42616 19780 42668 19786
rect 42616 19722 42668 19728
rect 42524 17060 42576 17066
rect 42524 17002 42576 17008
rect 42536 15026 42564 17002
rect 42524 15020 42576 15026
rect 42524 14962 42576 14968
rect 42628 6914 42656 19722
rect 42904 19446 42932 20198
rect 42892 19440 42944 19446
rect 42892 19382 42944 19388
rect 42996 19378 43024 20538
rect 43076 20460 43128 20466
rect 43076 20402 43128 20408
rect 43088 19514 43116 20402
rect 43076 19508 43128 19514
rect 43076 19450 43128 19456
rect 43180 19378 43208 20742
rect 43732 20534 43760 20878
rect 43824 20806 43852 21490
rect 43904 20936 43956 20942
rect 43904 20878 43956 20884
rect 43812 20800 43864 20806
rect 43812 20742 43864 20748
rect 43916 20534 43944 20878
rect 43720 20528 43772 20534
rect 43720 20470 43772 20476
rect 43904 20528 43956 20534
rect 43904 20470 43956 20476
rect 43536 20392 43588 20398
rect 43536 20334 43588 20340
rect 43444 19712 43496 19718
rect 43444 19654 43496 19660
rect 43456 19514 43484 19654
rect 43444 19508 43496 19514
rect 43444 19450 43496 19456
rect 42984 19372 43036 19378
rect 42984 19314 43036 19320
rect 43168 19372 43220 19378
rect 43168 19314 43220 19320
rect 43548 18222 43576 20334
rect 43732 19922 43760 20470
rect 43812 20052 43864 20058
rect 43812 19994 43864 20000
rect 43824 19922 43852 19994
rect 43720 19916 43772 19922
rect 43720 19858 43772 19864
rect 43812 19916 43864 19922
rect 43812 19858 43864 19864
rect 43720 19780 43772 19786
rect 43720 19722 43772 19728
rect 43536 18216 43588 18222
rect 43536 18158 43588 18164
rect 43628 17536 43680 17542
rect 43628 17478 43680 17484
rect 43640 17202 43668 17478
rect 43628 17196 43680 17202
rect 43628 17138 43680 17144
rect 42800 16516 42852 16522
rect 42800 16458 42852 16464
rect 42812 8090 42840 16458
rect 42800 8084 42852 8090
rect 42800 8026 42852 8032
rect 42536 6886 42656 6914
rect 43732 6914 43760 19722
rect 43824 15502 43852 19858
rect 43916 19786 43944 20470
rect 44008 20058 44036 21490
rect 44468 21418 44496 21966
rect 44364 21412 44416 21418
rect 44364 21354 44416 21360
rect 44456 21412 44508 21418
rect 44456 21354 44508 21360
rect 44272 21344 44324 21350
rect 44272 21286 44324 21292
rect 44180 20256 44232 20262
rect 44100 20216 44180 20244
rect 43996 20052 44048 20058
rect 43996 19994 44048 20000
rect 43904 19780 43956 19786
rect 43904 19722 43956 19728
rect 43996 19372 44048 19378
rect 44100 19360 44128 20216
rect 44180 20198 44232 20204
rect 44284 19378 44312 21286
rect 44376 21146 44404 21354
rect 44364 21140 44416 21146
rect 44364 21082 44416 21088
rect 44048 19332 44128 19360
rect 44272 19372 44324 19378
rect 43996 19314 44048 19320
rect 44272 19314 44324 19320
rect 43904 18216 43956 18222
rect 43904 18158 43956 18164
rect 43812 15496 43864 15502
rect 43812 15438 43864 15444
rect 43812 14952 43864 14958
rect 43812 14894 43864 14900
rect 43824 14618 43852 14894
rect 43812 14612 43864 14618
rect 43812 14554 43864 14560
rect 43732 6886 43852 6914
rect 42340 6860 42392 6866
rect 42340 6802 42392 6808
rect 42352 6186 42380 6802
rect 42340 6180 42392 6186
rect 42340 6122 42392 6128
rect 41696 4548 41748 4554
rect 41696 4490 41748 4496
rect 42248 4548 42300 4554
rect 42248 4490 42300 4496
rect 41788 3936 41840 3942
rect 41788 3878 41840 3884
rect 41604 2916 41656 2922
rect 41604 2858 41656 2864
rect 41800 2514 41828 3878
rect 42260 3466 42288 4490
rect 42432 4140 42484 4146
rect 42432 4082 42484 4088
rect 42444 3738 42472 4082
rect 42432 3732 42484 3738
rect 42432 3674 42484 3680
rect 42340 3664 42392 3670
rect 42340 3606 42392 3612
rect 42248 3460 42300 3466
rect 42248 3402 42300 3408
rect 42260 3126 42288 3402
rect 42248 3120 42300 3126
rect 42248 3062 42300 3068
rect 42352 2530 42380 3606
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42444 3058 42472 3470
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42536 2650 42564 6886
rect 42616 6656 42668 6662
rect 42616 6598 42668 6604
rect 42628 6254 42656 6598
rect 43824 6458 43852 6886
rect 43812 6452 43864 6458
rect 43812 6394 43864 6400
rect 42616 6248 42668 6254
rect 42616 6190 42668 6196
rect 42616 3936 42668 3942
rect 42616 3878 42668 3884
rect 42628 3126 42656 3878
rect 42616 3120 42668 3126
rect 42616 3062 42668 3068
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 42524 2644 42576 2650
rect 42524 2586 42576 2592
rect 40592 2508 40644 2514
rect 40592 2450 40644 2456
rect 41788 2508 41840 2514
rect 42352 2502 42564 2530
rect 41788 2450 41840 2456
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 41248 800 41276 2382
rect 42536 800 42564 2502
rect 43180 800 43208 2926
rect 43916 2922 43944 18158
rect 44008 17882 44036 19314
rect 43996 17876 44048 17882
rect 43996 17818 44048 17824
rect 44652 17814 44680 22066
rect 44732 21344 44784 21350
rect 44732 21286 44784 21292
rect 44744 21010 44772 21286
rect 44732 21004 44784 21010
rect 44732 20946 44784 20952
rect 44640 17808 44692 17814
rect 44640 17750 44692 17756
rect 44088 17604 44140 17610
rect 44088 17546 44140 17552
rect 44100 16726 44128 17546
rect 44272 17264 44324 17270
rect 44272 17206 44324 17212
rect 44088 16720 44140 16726
rect 44088 16662 44140 16668
rect 44284 16182 44312 17206
rect 44272 16176 44324 16182
rect 44272 16118 44324 16124
rect 44180 16040 44232 16046
rect 44180 15982 44232 15988
rect 44192 15706 44220 15982
rect 44180 15700 44232 15706
rect 44180 15642 44232 15648
rect 43996 15496 44048 15502
rect 43996 15438 44048 15444
rect 44008 14414 44036 15438
rect 43996 14408 44048 14414
rect 43996 14350 44048 14356
rect 44008 13938 44036 14350
rect 43996 13932 44048 13938
rect 43996 13874 44048 13880
rect 44836 8634 44864 24822
rect 44928 23798 44956 25842
rect 45008 25288 45060 25294
rect 45008 25230 45060 25236
rect 44916 23792 44968 23798
rect 44916 23734 44968 23740
rect 45020 23118 45048 25230
rect 45008 23112 45060 23118
rect 45008 23054 45060 23060
rect 45020 19446 45048 23054
rect 45192 22568 45244 22574
rect 45192 22510 45244 22516
rect 45100 22432 45152 22438
rect 45100 22374 45152 22380
rect 45112 21962 45140 22374
rect 45204 22234 45232 22510
rect 45192 22228 45244 22234
rect 45192 22170 45244 22176
rect 45100 21956 45152 21962
rect 45100 21898 45152 21904
rect 45284 21412 45336 21418
rect 45284 21354 45336 21360
rect 45296 20942 45324 21354
rect 45388 21162 45416 26206
rect 45468 25696 45520 25702
rect 45468 25638 45520 25644
rect 45480 25362 45508 25638
rect 45468 25356 45520 25362
rect 45468 25298 45520 25304
rect 45664 22438 45692 26551
rect 45848 25430 45876 38898
rect 46216 37806 46244 44338
rect 46308 43994 46336 44814
rect 46296 43988 46348 43994
rect 46296 43930 46348 43936
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 46296 38344 46348 38350
rect 46296 38286 46348 38292
rect 46308 37942 46336 38286
rect 46296 37936 46348 37942
rect 46296 37878 46348 37884
rect 46204 37800 46256 37806
rect 46204 37742 46256 37748
rect 46110 31376 46166 31385
rect 46110 31311 46166 31320
rect 46018 30016 46074 30025
rect 46018 29951 46074 29960
rect 45836 25424 45888 25430
rect 45836 25366 45888 25372
rect 46032 24410 46060 29951
rect 46020 24404 46072 24410
rect 46020 24346 46072 24352
rect 45744 23520 45796 23526
rect 45744 23462 45796 23468
rect 45756 23186 45784 23462
rect 45744 23180 45796 23186
rect 45744 23122 45796 23128
rect 45836 22704 45888 22710
rect 45836 22646 45888 22652
rect 45652 22432 45704 22438
rect 45652 22374 45704 22380
rect 45848 22234 45876 22646
rect 45928 22500 45980 22506
rect 45928 22442 45980 22448
rect 45468 22228 45520 22234
rect 45468 22170 45520 22176
rect 45652 22228 45704 22234
rect 45652 22170 45704 22176
rect 45836 22228 45888 22234
rect 45836 22170 45888 22176
rect 45480 22098 45508 22170
rect 45468 22092 45520 22098
rect 45468 22034 45520 22040
rect 45560 22024 45612 22030
rect 45560 21966 45612 21972
rect 45468 21616 45520 21622
rect 45572 21570 45600 21966
rect 45664 21894 45692 22170
rect 45940 22166 45968 22442
rect 45928 22160 45980 22166
rect 45928 22102 45980 22108
rect 45940 21978 45968 22102
rect 45848 21950 45968 21978
rect 46020 21956 46072 21962
rect 45652 21888 45704 21894
rect 45652 21830 45704 21836
rect 45520 21564 45600 21570
rect 45468 21558 45600 21564
rect 45480 21542 45600 21558
rect 45848 21554 45876 21950
rect 46020 21898 46072 21904
rect 46032 21690 46060 21898
rect 46020 21684 46072 21690
rect 46020 21626 46072 21632
rect 46124 21570 46152 31311
rect 46400 26234 46428 46951
rect 46664 46504 46716 46510
rect 46664 46446 46716 46452
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46492 45082 46520 45834
rect 46676 45558 46704 46446
rect 46664 45552 46716 45558
rect 46664 45494 46716 45500
rect 46768 45490 46796 47382
rect 46860 46510 46888 47631
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 48044 47184 48096 47190
rect 48044 47126 48096 47132
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47768 46368 47820 46374
rect 47964 46345 47992 46514
rect 47768 46310 47820 46316
rect 47950 46336 48006 46345
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 46756 45484 46808 45490
rect 46756 45426 46808 45432
rect 47308 45280 47360 45286
rect 47308 45222 47360 45228
rect 46480 45076 46532 45082
rect 46480 45018 46532 45024
rect 46664 44736 46716 44742
rect 46664 44678 46716 44684
rect 46676 41138 46704 44678
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 46952 43858 46980 44134
rect 46940 43852 46992 43858
rect 46940 43794 46992 43800
rect 46940 43104 46992 43110
rect 46940 43046 46992 43052
rect 46952 42770 46980 43046
rect 46940 42764 46992 42770
rect 46940 42706 46992 42712
rect 46940 41540 46992 41546
rect 46940 41482 46992 41488
rect 46952 41274 46980 41482
rect 46940 41268 46992 41274
rect 46940 41210 46992 41216
rect 46664 41132 46716 41138
rect 46664 41074 46716 41080
rect 46478 39536 46534 39545
rect 46478 39471 46534 39480
rect 46492 35894 46520 39471
rect 46676 38894 46704 41074
rect 46848 39364 46900 39370
rect 46848 39306 46900 39312
rect 46860 39098 46888 39306
rect 46848 39092 46900 39098
rect 46848 39034 46900 39040
rect 46664 38888 46716 38894
rect 46664 38830 46716 38836
rect 46756 38548 46808 38554
rect 46756 38490 46808 38496
rect 46768 37874 46796 38490
rect 46848 38276 46900 38282
rect 46848 38218 46900 38224
rect 46860 38010 46888 38218
rect 46848 38004 46900 38010
rect 46848 37946 46900 37952
rect 46756 37868 46808 37874
rect 46756 37810 46808 37816
rect 47032 37392 47084 37398
rect 47032 37334 47084 37340
rect 46492 35866 46612 35894
rect 46308 26206 46428 26234
rect 46204 25696 46256 25702
rect 46204 25638 46256 25644
rect 46216 24886 46244 25638
rect 46204 24880 46256 24886
rect 46204 24822 46256 24828
rect 46202 22536 46258 22545
rect 46202 22471 46258 22480
rect 45388 21134 45508 21162
rect 45284 20936 45336 20942
rect 45284 20878 45336 20884
rect 45376 20800 45428 20806
rect 45376 20742 45428 20748
rect 45388 20534 45416 20742
rect 45376 20528 45428 20534
rect 45376 20470 45428 20476
rect 45008 19440 45060 19446
rect 45008 19382 45060 19388
rect 45376 18692 45428 18698
rect 45376 18634 45428 18640
rect 45388 18290 45416 18634
rect 45376 18284 45428 18290
rect 45376 18226 45428 18232
rect 45376 17672 45428 17678
rect 45376 17614 45428 17620
rect 45284 17604 45336 17610
rect 45284 17546 45336 17552
rect 45296 17134 45324 17546
rect 45284 17128 45336 17134
rect 45284 17070 45336 17076
rect 45388 16522 45416 17614
rect 45376 16516 45428 16522
rect 45376 16458 45428 16464
rect 45100 14952 45152 14958
rect 45100 14894 45152 14900
rect 44824 8628 44876 8634
rect 44824 8570 44876 8576
rect 44836 8294 44864 8570
rect 44824 8288 44876 8294
rect 44824 8230 44876 8236
rect 44180 6384 44232 6390
rect 44180 6326 44232 6332
rect 44192 5710 44220 6326
rect 44180 5704 44232 5710
rect 44180 5646 44232 5652
rect 43904 2916 43956 2922
rect 43904 2858 43956 2864
rect 44192 2446 44220 5646
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 44180 2440 44232 2446
rect 44180 2382 44232 2388
rect 43824 800 43852 2382
rect 45112 800 45140 14894
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 45204 3058 45232 3470
rect 45480 3398 45508 21134
rect 45572 20806 45600 21542
rect 45836 21548 45888 21554
rect 45836 21490 45888 21496
rect 45940 21542 46152 21570
rect 46216 21554 46244 22471
rect 46308 22001 46336 26206
rect 46584 24886 46612 35866
rect 46848 33516 46900 33522
rect 46848 33458 46900 33464
rect 46664 33448 46716 33454
rect 46860 33425 46888 33458
rect 46664 33390 46716 33396
rect 46846 33416 46902 33425
rect 46676 31754 46704 33390
rect 46846 33351 46902 33360
rect 46940 32836 46992 32842
rect 46940 32778 46992 32784
rect 46952 32570 46980 32778
rect 46940 32564 46992 32570
rect 46940 32506 46992 32512
rect 46756 31884 46808 31890
rect 46756 31826 46808 31832
rect 46664 31748 46716 31754
rect 46664 31690 46716 31696
rect 46572 24880 46624 24886
rect 46572 24822 46624 24828
rect 46572 24744 46624 24750
rect 46572 24686 46624 24692
rect 46388 24676 46440 24682
rect 46388 24618 46440 24624
rect 46400 23905 46428 24618
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46386 23896 46442 23905
rect 46584 23866 46612 24686
rect 46386 23831 46442 23840
rect 46572 23860 46624 23866
rect 46572 23802 46624 23808
rect 46572 23520 46624 23526
rect 46572 23462 46624 23468
rect 46388 23180 46440 23186
rect 46388 23122 46440 23128
rect 46400 22778 46428 23122
rect 46388 22772 46440 22778
rect 46388 22714 46440 22720
rect 46400 22574 46428 22714
rect 46388 22568 46440 22574
rect 46388 22510 46440 22516
rect 46294 21992 46350 22001
rect 46294 21927 46350 21936
rect 46296 21888 46348 21894
rect 46296 21830 46348 21836
rect 46308 21554 46336 21830
rect 46204 21548 46256 21554
rect 45560 20800 45612 20806
rect 45560 20742 45612 20748
rect 45652 19508 45704 19514
rect 45652 19450 45704 19456
rect 45560 18624 45612 18630
rect 45560 18566 45612 18572
rect 45572 18426 45600 18566
rect 45560 18420 45612 18426
rect 45560 18362 45612 18368
rect 45560 18080 45612 18086
rect 45560 18022 45612 18028
rect 45572 17270 45600 18022
rect 45664 17678 45692 19450
rect 45744 19372 45796 19378
rect 45744 19314 45796 19320
rect 45756 18465 45784 19314
rect 45848 18970 45876 21490
rect 45940 19718 45968 21542
rect 46204 21490 46256 21496
rect 46296 21548 46348 21554
rect 46296 21490 46348 21496
rect 46112 21480 46164 21486
rect 46112 21422 46164 21428
rect 46020 20800 46072 20806
rect 46020 20742 46072 20748
rect 45928 19712 45980 19718
rect 45928 19654 45980 19660
rect 45836 18964 45888 18970
rect 45836 18906 45888 18912
rect 45836 18760 45888 18766
rect 45836 18702 45888 18708
rect 45742 18456 45798 18465
rect 45742 18391 45798 18400
rect 45848 18290 45876 18702
rect 45836 18284 45888 18290
rect 45836 18226 45888 18232
rect 45652 17672 45704 17678
rect 45652 17614 45704 17620
rect 45560 17264 45612 17270
rect 45560 17206 45612 17212
rect 45664 16658 45692 17614
rect 45744 17332 45796 17338
rect 45744 17274 45796 17280
rect 45756 17134 45784 17274
rect 45744 17128 45796 17134
rect 45744 17070 45796 17076
rect 45652 16652 45704 16658
rect 45652 16594 45704 16600
rect 45836 16040 45888 16046
rect 45836 15982 45888 15988
rect 45558 15736 45614 15745
rect 45558 15671 45614 15680
rect 45572 15638 45600 15671
rect 45560 15632 45612 15638
rect 45560 15574 45612 15580
rect 45560 8492 45612 8498
rect 45560 8434 45612 8440
rect 45572 7698 45600 8434
rect 45652 8288 45704 8294
rect 45652 8230 45704 8236
rect 45664 7886 45692 8230
rect 45652 7880 45704 7886
rect 45652 7822 45704 7828
rect 45572 7670 45692 7698
rect 45664 7478 45692 7670
rect 45652 7472 45704 7478
rect 45652 7414 45704 7420
rect 45560 7336 45612 7342
rect 45560 7278 45612 7284
rect 45572 6662 45600 7278
rect 45560 6656 45612 6662
rect 45560 6598 45612 6604
rect 45664 4758 45692 7414
rect 45652 4752 45704 4758
rect 45652 4694 45704 4700
rect 45744 4480 45796 4486
rect 45744 4422 45796 4428
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45756 3126 45784 4422
rect 45848 3505 45876 15982
rect 45928 7812 45980 7818
rect 45928 7754 45980 7760
rect 45940 7546 45968 7754
rect 45928 7540 45980 7546
rect 45928 7482 45980 7488
rect 46032 6798 46060 20742
rect 46124 19990 46152 21422
rect 46400 20398 46428 22510
rect 46480 22092 46532 22098
rect 46480 22034 46532 22040
rect 46492 20602 46520 22034
rect 46584 21622 46612 23462
rect 46572 21616 46624 21622
rect 46572 21558 46624 21564
rect 46480 20596 46532 20602
rect 46480 20538 46532 20544
rect 46572 20460 46624 20466
rect 46572 20402 46624 20408
rect 46388 20392 46440 20398
rect 46388 20334 46440 20340
rect 46112 19984 46164 19990
rect 46112 19926 46164 19932
rect 46584 19922 46612 20402
rect 46572 19916 46624 19922
rect 46572 19858 46624 19864
rect 46296 19168 46348 19174
rect 46296 19110 46348 19116
rect 46308 18834 46336 19110
rect 46112 18828 46164 18834
rect 46112 18770 46164 18776
rect 46296 18828 46348 18834
rect 46296 18770 46348 18776
rect 46124 18290 46152 18770
rect 46112 18284 46164 18290
rect 46112 18226 46164 18232
rect 46204 18216 46256 18222
rect 46204 18158 46256 18164
rect 46216 6914 46244 18158
rect 46572 16720 46624 16726
rect 46572 16662 46624 16668
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 46308 12850 46336 13262
rect 46296 12844 46348 12850
rect 46296 12786 46348 12792
rect 46480 10464 46532 10470
rect 46480 10406 46532 10412
rect 46492 10130 46520 10406
rect 46480 10124 46532 10130
rect 46480 10066 46532 10072
rect 46584 7954 46612 16662
rect 46676 9450 46704 31690
rect 46768 24970 46796 31826
rect 46846 28656 46902 28665
rect 46846 28591 46902 28600
rect 46860 28218 46888 28591
rect 46940 28552 46992 28558
rect 46940 28494 46992 28500
rect 46848 28212 46900 28218
rect 46848 28154 46900 28160
rect 46952 27606 46980 28494
rect 47044 28082 47072 37334
rect 47124 35488 47176 35494
rect 47124 35430 47176 35436
rect 47136 34066 47164 35430
rect 47216 34400 47268 34406
rect 47216 34342 47268 34348
rect 47124 34060 47176 34066
rect 47124 34002 47176 34008
rect 47228 33930 47256 34342
rect 47216 33924 47268 33930
rect 47216 33866 47268 33872
rect 47216 29708 47268 29714
rect 47216 29650 47268 29656
rect 47032 28076 47084 28082
rect 47032 28018 47084 28024
rect 46940 27600 46992 27606
rect 46940 27542 46992 27548
rect 46846 25936 46902 25945
rect 46846 25871 46902 25880
rect 46860 25362 46888 25871
rect 46848 25356 46900 25362
rect 46848 25298 46900 25304
rect 47030 25256 47086 25265
rect 47030 25191 47086 25200
rect 46768 24942 46888 24970
rect 46756 24880 46808 24886
rect 46756 24822 46808 24828
rect 46768 22098 46796 24822
rect 46756 22092 46808 22098
rect 46756 22034 46808 22040
rect 46860 20482 46888 24942
rect 47044 24886 47072 25191
rect 47032 24880 47084 24886
rect 47032 24822 47084 24828
rect 47032 23724 47084 23730
rect 47032 23666 47084 23672
rect 47044 23225 47072 23666
rect 47030 23216 47086 23225
rect 47030 23151 47086 23160
rect 47228 22438 47256 29650
rect 47320 23118 47348 45222
rect 47492 45008 47544 45014
rect 47492 44950 47544 44956
rect 47504 42226 47532 44950
rect 47676 44804 47728 44810
rect 47676 44746 47728 44752
rect 47688 44538 47716 44746
rect 47676 44532 47728 44538
rect 47676 44474 47728 44480
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47492 42220 47544 42226
rect 47492 42162 47544 42168
rect 47400 34060 47452 34066
rect 47400 34002 47452 34008
rect 47412 31890 47440 34002
rect 47400 31884 47452 31890
rect 47400 31826 47452 31832
rect 47400 29640 47452 29646
rect 47400 29582 47452 29588
rect 47412 29345 47440 29582
rect 47398 29336 47454 29345
rect 47398 29271 47454 29280
rect 47400 28076 47452 28082
rect 47400 28018 47452 28024
rect 47308 23112 47360 23118
rect 47308 23054 47360 23060
rect 47216 22432 47268 22438
rect 47216 22374 47268 22380
rect 47228 21350 47256 22374
rect 47216 21344 47268 21350
rect 47216 21286 47268 21292
rect 46768 20454 46888 20482
rect 46768 19446 46796 20454
rect 46756 19440 46808 19446
rect 46756 19382 46808 19388
rect 46940 19168 46992 19174
rect 46940 19110 46992 19116
rect 46756 18896 46808 18902
rect 46756 18838 46808 18844
rect 46768 10985 46796 18838
rect 46952 18834 46980 19110
rect 46940 18828 46992 18834
rect 46940 18770 46992 18776
rect 47412 18290 47440 28018
rect 47504 24818 47532 42162
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 40730 47716 41618
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47780 35894 47808 46310
rect 47950 46271 48006 46280
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47860 38956 47912 38962
rect 47860 38898 47912 38904
rect 47872 38865 47900 38898
rect 47858 38856 47914 38865
rect 47858 38791 47914 38800
rect 47780 35866 47992 35894
rect 47860 34944 47912 34950
rect 47860 34886 47912 34892
rect 47768 34604 47820 34610
rect 47768 34546 47820 34552
rect 47780 33658 47808 34546
rect 47768 33652 47820 33658
rect 47768 33594 47820 33600
rect 47872 33318 47900 34886
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 47964 33130 47992 35866
rect 47872 33102 47992 33130
rect 48056 33130 48084 47126
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48134 41576 48190 41585
rect 48134 41511 48136 41520
rect 48188 41511 48190 41520
rect 48136 41482 48188 41488
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48136 38276 48188 38282
rect 48136 38218 48188 38224
rect 48148 38185 48176 38218
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48136 35692 48188 35698
rect 48136 35634 48188 35640
rect 48148 34785 48176 35634
rect 48228 35080 48280 35086
rect 48228 35022 48280 35028
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48240 34105 48268 35022
rect 48226 34096 48282 34105
rect 48226 34031 48282 34040
rect 48056 33102 48268 33130
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27538 47716 27814
rect 47676 27532 47728 27538
rect 47676 27474 47728 27480
rect 47768 25288 47820 25294
rect 47768 25230 47820 25236
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47504 21078 47532 24754
rect 47780 24342 47808 25230
rect 47768 24336 47820 24342
rect 47768 24278 47820 24284
rect 47584 23724 47636 23730
rect 47584 23666 47636 23672
rect 47596 21146 47624 23666
rect 47584 21140 47636 21146
rect 47584 21082 47636 21088
rect 47492 21072 47544 21078
rect 47492 21014 47544 21020
rect 47504 19378 47532 21014
rect 47492 19372 47544 19378
rect 47492 19314 47544 19320
rect 47400 18284 47452 18290
rect 47400 18226 47452 18232
rect 47032 18080 47084 18086
rect 47032 18022 47084 18028
rect 47044 17746 47072 18022
rect 47032 17740 47084 17746
rect 47032 17682 47084 17688
rect 47596 17202 47624 21082
rect 47676 19780 47728 19786
rect 47676 19722 47728 19728
rect 47688 19514 47716 19722
rect 47676 19508 47728 19514
rect 47676 19450 47728 19456
rect 47872 18698 47900 33102
rect 48044 33040 48096 33046
rect 48044 32982 48096 32988
rect 48056 32570 48084 32982
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48044 32564 48096 32570
rect 48044 32506 48096 32512
rect 47952 32428 48004 32434
rect 47952 32370 48004 32376
rect 47964 32065 47992 32370
rect 47950 32056 48006 32065
rect 48240 32026 48268 33102
rect 47950 31991 48006 32000
rect 48228 32020 48280 32026
rect 48228 31962 48280 31968
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48044 23656 48096 23662
rect 48044 23598 48096 23604
rect 47952 23044 48004 23050
rect 47952 22986 48004 22992
rect 47964 21865 47992 22986
rect 48056 22778 48084 23598
rect 48044 22772 48096 22778
rect 48044 22714 48096 22720
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48136 19780 48188 19786
rect 48136 19722 48188 19728
rect 48148 19145 48176 19722
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 47860 18692 47912 18698
rect 47860 18634 47912 18640
rect 48044 18216 48096 18222
rect 48044 18158 48096 18164
rect 47676 18080 47728 18086
rect 47676 18022 47728 18028
rect 47688 17610 47716 18022
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 47584 17196 47636 17202
rect 47584 17138 47636 17144
rect 47596 12434 47624 17138
rect 47676 16992 47728 16998
rect 47676 16934 47728 16940
rect 47688 16522 47716 16934
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47780 16114 47808 16594
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47676 13728 47728 13734
rect 47676 13670 47728 13676
rect 47688 13394 47716 13670
rect 47676 13388 47728 13394
rect 47676 13330 47728 13336
rect 47504 12406 47624 12434
rect 46754 10976 46810 10985
rect 46754 10911 46810 10920
rect 47504 10674 47532 12406
rect 47676 11144 47728 11150
rect 47676 11086 47728 11092
rect 47492 10668 47544 10674
rect 47492 10610 47544 10616
rect 46664 9444 46716 9450
rect 46664 9386 46716 9392
rect 46846 8256 46902 8265
rect 46846 8191 46902 8200
rect 46860 8090 46888 8191
rect 46848 8084 46900 8090
rect 46848 8026 46900 8032
rect 46572 7948 46624 7954
rect 46572 7890 46624 7896
rect 46584 7478 46612 7890
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 46572 7472 46624 7478
rect 46572 7414 46624 7420
rect 46216 6886 46612 6914
rect 46020 6792 46072 6798
rect 46020 6734 46072 6740
rect 46388 4208 46440 4214
rect 46388 4150 46440 4156
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3602 46336 3878
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 45834 3496 45890 3505
rect 45834 3431 45890 3440
rect 45744 3120 45796 3126
rect 45744 3062 45796 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45468 2304 45520 2310
rect 45468 2246 45520 2252
rect 45480 1970 45508 2246
rect 45468 1964 45520 1970
rect 45468 1906 45520 1912
rect 46400 800 46428 4150
rect 46584 2514 46612 6886
rect 47320 6866 47348 7511
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 47504 4690 47532 10610
rect 47688 10198 47716 11086
rect 47676 10192 47728 10198
rect 47676 10134 47728 10140
rect 47858 9616 47914 9625
rect 47858 9551 47860 9560
rect 47912 9551 47914 9560
rect 47860 9522 47912 9528
rect 47766 8936 47822 8945
rect 47766 8871 47768 8880
rect 47820 8871 47822 8880
rect 47768 8842 47820 8848
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 47964 6225 47992 6258
rect 47950 6216 48006 6225
rect 47950 6151 48006 6160
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 47492 4684 47544 4690
rect 47492 4626 47544 4632
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46756 4208 46808 4214
rect 46860 4185 46888 4558
rect 46756 4150 46808 4156
rect 46846 4176 46902 4185
rect 46662 4040 46718 4049
rect 46662 3975 46718 3984
rect 46676 3942 46704 3975
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 30576 734 30788 762
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46768 105 46796 4150
rect 46846 4111 46902 4120
rect 47780 3505 47808 5170
rect 47766 3496 47822 3505
rect 47766 3431 47822 3440
rect 48056 3194 48084 18158
rect 48228 17604 48280 17610
rect 48228 17546 48280 17552
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48148 16658 48176 17031
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 48240 16425 48268 17546
rect 48226 16416 48282 16425
rect 48226 16351 48282 16360
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 48148 12345 48176 13194
rect 48134 12336 48190 12345
rect 48134 12271 48190 12280
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48134 6831 48190 6840
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 48320 3052 48372 3058
rect 48320 2994 48372 3000
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 46848 2372 46900 2378
rect 46848 2314 46900 2320
rect 46860 1465 46888 2314
rect 46846 1456 46902 1465
rect 46846 1391 46902 1400
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48056 785 48084 2382
rect 48332 800 48360 2994
rect 48976 800 49004 3402
rect 48042 776 48098 785
rect 48042 711 48098 720
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1398 47640 1454 47696
rect 3790 46960 3846 47016
rect 1398 42880 1454 42936
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 2778 46280 2834 46336
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3422 44920 3478 44976
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1582 35400 1638 35456
rect 1582 32680 1638 32736
rect 1858 32000 1914 32056
rect 2778 36760 2834 36816
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 1858 23160 1914 23216
rect 2226 19080 2282 19136
rect 3514 43560 3570 43616
rect 3698 39480 3754 39536
rect 3514 31320 3570 31376
rect 3514 30232 3570 30288
rect 3514 28600 3570 28656
rect 1858 17720 1914 17776
rect 1858 16360 1914 16416
rect 1398 12280 1454 12336
rect 2778 15000 2834 15056
rect 3514 7520 3570 7576
rect 3882 29144 3938 29200
rect 3974 19760 4030 19816
rect 3974 18420 4030 18456
rect 3974 18400 3976 18420
rect 3976 18400 4028 18420
rect 4028 18400 4030 18420
rect 3974 17040 4030 17096
rect 3974 13640 4030 13696
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4066 10240 4122 10296
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 14830 24112 14886 24168
rect 15382 24132 15438 24168
rect 15382 24112 15384 24132
rect 15384 24112 15436 24132
rect 15436 24112 15438 24132
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3440 4122 3496
rect 3238 1400 3294 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19522 46980 19578 47016
rect 19522 46960 19524 46980
rect 19524 46960 19576 46980
rect 19576 46960 19578 46980
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 17130 35572 17132 35592
rect 17132 35572 17184 35592
rect 17184 35572 17186 35592
rect 17130 35536 17186 35572
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 17406 3440 17462 3496
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19798 19388 19800 19408
rect 19800 19388 19852 19408
rect 19852 19388 19854 19408
rect 19798 19352 19854 19388
rect 20166 19624 20222 19680
rect 20350 19624 20406 19680
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20626 19624 20682 19680
rect 27066 46824 27122 46880
rect 22650 35692 22706 35728
rect 22650 35672 22652 35692
rect 22652 35672 22704 35692
rect 22704 35672 22706 35692
rect 24490 34720 24546 34776
rect 20718 19488 20774 19544
rect 20534 19352 20590 19408
rect 22006 19488 22062 19544
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 18694 3712 18750 3768
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19246 2896 19302 2952
rect 20074 3304 20130 3360
rect 20902 3712 20958 3768
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 2870 720 2926 776
rect 23018 3984 23074 4040
rect 20718 2896 20774 2952
rect 24214 31456 24270 31512
rect 24766 31456 24822 31512
rect 24858 19352 24914 19408
rect 24674 3304 24730 3360
rect 24122 2916 24178 2952
rect 24122 2896 24124 2916
rect 24124 2896 24176 2916
rect 24176 2896 24178 2916
rect 25042 20324 25098 20360
rect 25042 20304 25044 20324
rect 25044 20304 25096 20324
rect 25096 20304 25098 20324
rect 25042 3304 25098 3360
rect 26514 34720 26570 34776
rect 26146 31456 26202 31512
rect 25502 20712 25558 20768
rect 25870 20712 25926 20768
rect 25870 19488 25926 19544
rect 26330 20304 26386 20360
rect 25686 19352 25742 19408
rect 28998 35672 29054 35728
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 27618 3576 27674 3632
rect 27618 2916 27674 2952
rect 27618 2896 27620 2916
rect 27620 2896 27672 2916
rect 27672 2896 27674 2916
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34886 30232 34942 30288
rect 33138 29144 33194 29200
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 33414 21020 33416 21040
rect 33416 21020 33468 21040
rect 33468 21020 33470 21040
rect 33414 20984 33470 21020
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35346 21548 35402 21584
rect 35346 21528 35348 21548
rect 35348 21528 35400 21548
rect 35400 21528 35402 21548
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38014 20984 38070 21040
rect 40314 24112 40370 24168
rect 44086 35536 44142 35592
rect 46846 47640 46902 47696
rect 46386 46960 46442 47016
rect 45650 26560 45706 26616
rect 46110 31320 46166 31376
rect 46018 29960 46074 30016
rect 46478 39480 46534 39536
rect 46202 22480 46258 22536
rect 46846 33360 46902 33416
rect 46386 23840 46442 23896
rect 46294 21936 46350 21992
rect 45742 18400 45798 18456
rect 45558 15680 45614 15736
rect 46846 28600 46902 28656
rect 46846 25880 46902 25936
rect 47030 25200 47086 25256
rect 47030 23160 47086 23216
rect 47398 29280 47454 29336
rect 47950 46280 48006 46336
rect 47950 40840 48006 40896
rect 47858 38800 47914 38856
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41540 48190 41576
rect 48134 41520 48136 41540
rect 48136 41520 48188 41540
rect 48188 41520 48190 41540
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48226 34040 48282 34096
rect 48134 32680 48190 32736
rect 47950 32000 48006 32056
rect 48134 27920 48190 27976
rect 48134 24520 48190 24576
rect 47950 21800 48006 21856
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 46754 10920 46810 10976
rect 46846 8200 46902 8256
rect 47306 7520 47362 7576
rect 45834 3440 45890 3496
rect 47858 9580 47914 9616
rect 47858 9560 47860 9580
rect 47860 9560 47912 9580
rect 47912 9560 47914 9580
rect 47766 8900 47822 8936
rect 47766 8880 47768 8900
rect 47768 8880 47820 8900
rect 47820 8880 47822 8900
rect 47950 6160 48006 6216
rect 46662 3984 46718 4040
rect 46846 4120 46902 4176
rect 47766 3440 47822 3496
rect 48134 17040 48190 17096
rect 48226 16360 48282 16416
rect 48134 12280 48190 12336
rect 48134 10240 48190 10296
rect 48134 6840 48190 6896
rect 46846 1400 46902 1456
rect 46754 40 46810 96
rect 48042 720 48098 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47548 800 47638
rect 1393 47635 1459 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3785 47018 3851 47021
rect 0 47016 3851 47018
rect 0 46960 3790 47016
rect 3846 46960 3851 47016
rect 0 46958 3851 46960
rect 0 46868 800 46958
rect 3785 46955 3851 46958
rect 19517 47018 19583 47021
rect 20110 47018 20116 47020
rect 19517 47016 20116 47018
rect 19517 46960 19522 47016
rect 19578 46960 20116 47016
rect 19517 46958 20116 46960
rect 19517 46955 19583 46958
rect 20110 46956 20116 46958
rect 20180 46956 20186 47020
rect 46381 47018 46447 47021
rect 49200 47018 50000 47108
rect 46381 47016 50000 47018
rect 46381 46960 46386 47016
rect 46442 46960 50000 47016
rect 46381 46958 50000 46960
rect 46381 46955 46447 46958
rect 27061 46882 27127 46885
rect 27470 46882 27476 46884
rect 27061 46880 27476 46882
rect 27061 46824 27066 46880
rect 27122 46824 27476 46880
rect 27061 46822 27476 46824
rect 27061 46819 27127 46822
rect 27470 46820 27476 46822
rect 27540 46820 27546 46884
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3417 44978 3483 44981
rect 0 44976 3483 44978
rect 0 44920 3422 44976
rect 3478 44920 3483 44976
rect 0 44918 3483 44920
rect 0 44828 800 44918
rect 3417 44915 3483 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3509 43618 3575 43621
rect 0 43616 3575 43618
rect 0 43560 3514 43616
rect 3570 43560 3575 43616
rect 0 43558 3575 43560
rect 0 43468 800 43558
rect 3509 43555 3575 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3693 39538 3759 39541
rect 0 39536 3759 39538
rect 0 39480 3698 39536
rect 3754 39480 3759 39536
rect 0 39478 3759 39480
rect 0 39388 800 39478
rect 3693 39475 3759 39478
rect 46473 39538 46539 39541
rect 49200 39538 50000 39628
rect 46473 39536 50000 39538
rect 46473 39480 46478 39536
rect 46534 39480 50000 39536
rect 46473 39478 50000 39480
rect 46473 39475 46539 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47853 38858 47919 38861
rect 49200 38858 50000 38948
rect 47853 38856 50000 38858
rect 47853 38800 47858 38856
rect 47914 38800 50000 38856
rect 47853 38798 50000 38800
rect 47853 38795 47919 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 22645 35730 22711 35733
rect 28993 35730 29059 35733
rect 22645 35728 29059 35730
rect 22645 35672 22650 35728
rect 22706 35672 28998 35728
rect 29054 35672 29059 35728
rect 22645 35670 29059 35672
rect 22645 35667 22711 35670
rect 28993 35667 29059 35670
rect 17125 35594 17191 35597
rect 44081 35594 44147 35597
rect 17125 35592 44147 35594
rect 0 35458 800 35548
rect 17125 35536 17130 35592
rect 17186 35536 44086 35592
rect 44142 35536 44147 35592
rect 17125 35534 44147 35536
rect 17125 35531 17191 35534
rect 44081 35531 44147 35534
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 24485 34778 24551 34781
rect 26509 34778 26575 34781
rect 24485 34776 26575 34778
rect 24485 34720 24490 34776
rect 24546 34720 26514 34776
rect 26570 34720 26575 34776
rect 24485 34718 26575 34720
rect 24485 34715 24551 34718
rect 26509 34715 26575 34718
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48221 34098 48287 34101
rect 49200 34098 50000 34188
rect 48221 34096 50000 34098
rect 48221 34040 48226 34096
rect 48282 34040 50000 34096
rect 48221 34038 50000 34040
rect 48221 34035 48287 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 46841 33418 46907 33421
rect 49200 33418 50000 33508
rect 46841 33416 50000 33418
rect 46841 33360 46846 33416
rect 46902 33360 50000 33416
rect 46841 33358 50000 33360
rect 46841 33355 46907 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 47945 32058 48011 32061
rect 49200 32058 50000 32148
rect 47945 32056 50000 32058
rect 47945 32000 47950 32056
rect 48006 32000 50000 32056
rect 47945 31998 50000 32000
rect 47945 31995 48011 31998
rect 49200 31908 50000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 24209 31514 24275 31517
rect 24761 31514 24827 31517
rect 26141 31514 26207 31517
rect 24209 31512 26207 31514
rect 0 31378 800 31468
rect 24209 31456 24214 31512
rect 24270 31456 24766 31512
rect 24822 31456 26146 31512
rect 26202 31456 26207 31512
rect 24209 31454 26207 31456
rect 24209 31451 24275 31454
rect 24761 31451 24827 31454
rect 26141 31451 26207 31454
rect 3509 31378 3575 31381
rect 0 31376 3575 31378
rect 0 31320 3514 31376
rect 3570 31320 3575 31376
rect 0 31318 3575 31320
rect 0 31228 800 31318
rect 3509 31315 3575 31318
rect 46105 31378 46171 31381
rect 49200 31378 50000 31468
rect 46105 31376 50000 31378
rect 46105 31320 46110 31376
rect 46166 31320 50000 31376
rect 46105 31318 50000 31320
rect 46105 31315 46171 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 3509 30290 3575 30293
rect 34881 30290 34947 30293
rect 3509 30288 34947 30290
rect 3509 30232 3514 30288
rect 3570 30232 34886 30288
rect 34942 30232 34947 30288
rect 3509 30230 34947 30232
rect 3509 30227 3575 30230
rect 34881 30227 34947 30230
rect 0 29868 800 30108
rect 46013 30018 46079 30021
rect 49200 30018 50000 30108
rect 46013 30016 50000 30018
rect 46013 29960 46018 30016
rect 46074 29960 50000 30016
rect 46013 29958 50000 29960
rect 46013 29955 46079 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47393 29338 47459 29341
rect 49200 29338 50000 29428
rect 47393 29336 50000 29338
rect 47393 29280 47398 29336
rect 47454 29280 50000 29336
rect 47393 29278 50000 29280
rect 47393 29275 47459 29278
rect 3877 29202 3943 29205
rect 33133 29202 33199 29205
rect 3877 29200 33199 29202
rect 3877 29144 3882 29200
rect 3938 29144 33138 29200
rect 33194 29144 33199 29200
rect 49200 29188 50000 29278
rect 3877 29142 33199 29144
rect 3877 29139 3943 29142
rect 33133 29139 33199 29142
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3509 28658 3575 28661
rect 0 28656 3575 28658
rect 0 28600 3514 28656
rect 3570 28600 3575 28656
rect 0 28598 3575 28600
rect 0 28508 800 28598
rect 3509 28595 3575 28598
rect 46841 28658 46907 28661
rect 49200 28658 50000 28748
rect 46841 28656 50000 28658
rect 46841 28600 46846 28656
rect 46902 28600 50000 28656
rect 46841 28598 50000 28600
rect 46841 28595 46907 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 45645 26618 45711 26621
rect 49200 26618 50000 26708
rect 45645 26616 50000 26618
rect 45645 26560 45650 26616
rect 45706 26560 50000 26616
rect 45645 26558 50000 26560
rect 45645 26555 45711 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 46841 25938 46907 25941
rect 49200 25938 50000 26028
rect 46841 25936 50000 25938
rect 46841 25880 46846 25936
rect 46902 25880 50000 25936
rect 46841 25878 50000 25880
rect 46841 25875 46907 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 47025 25258 47091 25261
rect 49200 25258 50000 25348
rect 47025 25256 50000 25258
rect 47025 25200 47030 25256
rect 47086 25200 50000 25256
rect 47025 25198 50000 25200
rect 47025 25195 47091 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 14825 24170 14891 24173
rect 15377 24170 15443 24173
rect 14825 24168 15443 24170
rect 14825 24112 14830 24168
rect 14886 24112 15382 24168
rect 15438 24112 15443 24168
rect 14825 24110 15443 24112
rect 14825 24107 14891 24110
rect 15377 24107 15443 24110
rect 27470 24108 27476 24172
rect 27540 24170 27546 24172
rect 40309 24170 40375 24173
rect 27540 24168 40375 24170
rect 27540 24112 40314 24168
rect 40370 24112 40375 24168
rect 27540 24110 40375 24112
rect 27540 24108 27546 24110
rect 40309 24107 40375 24110
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46381 23898 46447 23901
rect 49200 23898 50000 23988
rect 46381 23896 50000 23898
rect 46381 23840 46386 23896
rect 46442 23840 50000 23896
rect 46381 23838 50000 23840
rect 46381 23835 46447 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 47025 23218 47091 23221
rect 49200 23218 50000 23308
rect 47025 23216 50000 23218
rect 47025 23160 47030 23216
rect 47086 23160 50000 23216
rect 47025 23158 50000 23160
rect 47025 23155 47091 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46197 22538 46263 22541
rect 49200 22538 50000 22628
rect 46197 22536 50000 22538
rect 46197 22480 46202 22536
rect 46258 22480 50000 22536
rect 46197 22478 50000 22480
rect 46197 22475 46263 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 46289 21994 46355 21997
rect 41370 21992 46355 21994
rect 0 21708 800 21948
rect 41370 21936 46294 21992
rect 46350 21936 46355 21992
rect 41370 21934 46355 21936
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 35341 21586 35407 21589
rect 41370 21586 41430 21934
rect 46289 21931 46355 21934
rect 47945 21858 48011 21861
rect 49200 21858 50000 21948
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 49200 21708 50000 21798
rect 35341 21584 41430 21586
rect 35341 21528 35346 21584
rect 35402 21528 41430 21584
rect 35341 21526 41430 21528
rect 35341 21523 35407 21526
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 33409 21042 33475 21045
rect 38009 21042 38075 21045
rect 33409 21040 38075 21042
rect 33409 20984 33414 21040
rect 33470 20984 38014 21040
rect 38070 20984 38075 21040
rect 49200 21028 50000 21118
rect 33409 20982 38075 20984
rect 33409 20979 33475 20982
rect 38009 20979 38075 20982
rect 25497 20770 25563 20773
rect 25865 20770 25931 20773
rect 25497 20768 25931 20770
rect 25497 20712 25502 20768
rect 25558 20712 25870 20768
rect 25926 20712 25931 20768
rect 25497 20710 25931 20712
rect 25497 20707 25563 20710
rect 25865 20707 25931 20710
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 25037 20362 25103 20365
rect 26325 20362 26391 20365
rect 25037 20360 26391 20362
rect 25037 20304 25042 20360
rect 25098 20304 26330 20360
rect 26386 20304 26391 20360
rect 25037 20302 26391 20304
rect 25037 20299 25103 20302
rect 26325 20299 26391 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19668 800 19758
rect 3969 19755 4035 19758
rect 20161 19682 20227 19685
rect 20345 19682 20411 19685
rect 20621 19682 20687 19685
rect 20161 19680 20687 19682
rect 20161 19624 20166 19680
rect 20222 19624 20350 19680
rect 20406 19624 20626 19680
rect 20682 19624 20687 19680
rect 49200 19668 50000 19908
rect 20161 19622 20687 19624
rect 20161 19619 20227 19622
rect 20345 19619 20411 19622
rect 20621 19619 20687 19622
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 20713 19546 20779 19549
rect 22001 19546 22067 19549
rect 25865 19546 25931 19549
rect 20713 19544 25931 19546
rect 20713 19488 20718 19544
rect 20774 19488 22006 19544
rect 22062 19488 25870 19544
rect 25926 19488 25931 19544
rect 20713 19486 25931 19488
rect 20713 19483 20779 19486
rect 22001 19483 22067 19486
rect 25865 19483 25931 19486
rect 19793 19410 19859 19413
rect 20529 19410 20595 19413
rect 19793 19408 20595 19410
rect 19793 19352 19798 19408
rect 19854 19352 20534 19408
rect 20590 19352 20595 19408
rect 19793 19350 20595 19352
rect 19793 19347 19859 19350
rect 20529 19347 20595 19350
rect 24853 19410 24919 19413
rect 25681 19410 25747 19413
rect 24853 19408 25747 19410
rect 24853 19352 24858 19408
rect 24914 19352 25686 19408
rect 25742 19352 25747 19408
rect 24853 19350 25747 19352
rect 24853 19347 24919 19350
rect 25681 19347 25747 19350
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18308 800 18398
rect 3969 18395 4035 18398
rect 45737 18458 45803 18461
rect 49200 18458 50000 18548
rect 45737 18456 50000 18458
rect 45737 18400 45742 18456
rect 45798 18400 50000 18456
rect 45737 18398 50000 18400
rect 45737 18395 45803 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1853 17778 1919 17781
rect 0 17776 1919 17778
rect 0 17720 1858 17776
rect 1914 17720 1919 17776
rect 0 17718 1919 17720
rect 0 17628 800 17718
rect 1853 17715 1919 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3969 17098 4035 17101
rect 0 17096 4035 17098
rect 0 17040 3974 17096
rect 4030 17040 4035 17096
rect 0 17038 4035 17040
rect 0 16948 800 17038
rect 3969 17035 4035 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 48221 16418 48287 16421
rect 49200 16418 50000 16508
rect 48221 16416 50000 16418
rect 48221 16360 48226 16416
rect 48282 16360 50000 16416
rect 48221 16358 50000 16360
rect 48221 16355 48287 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3969 13698 4035 13701
rect 0 13696 4035 13698
rect 0 13640 3974 13696
rect 4030 13640 4035 13696
rect 0 13638 4035 13640
rect 0 13548 800 13638
rect 3969 13635 4035 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 46749 10978 46815 10981
rect 49200 10978 50000 11068
rect 46749 10976 50000 10978
rect 46749 10920 46754 10976
rect 46810 10920 50000 10976
rect 46749 10918 50000 10920
rect 46749 10915 46815 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 4061 10298 4127 10301
rect 0 10296 4127 10298
rect 0 10240 4066 10296
rect 4122 10240 4127 10296
rect 0 10238 4127 10240
rect 0 10148 800 10238
rect 4061 10235 4127 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 47853 9618 47919 9621
rect 49200 9618 50000 9708
rect 47853 9616 50000 9618
rect 47853 9560 47858 9616
rect 47914 9560 50000 9616
rect 47853 9558 50000 9560
rect 47853 9555 47919 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 46841 8258 46907 8261
rect 49200 8258 50000 8348
rect 46841 8256 50000 8258
rect 46841 8200 46846 8256
rect 46902 8200 50000 8256
rect 46841 8198 50000 8200
rect 46841 8195 46907 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3509 7578 3575 7581
rect 0 7576 3575 7578
rect 0 7520 3514 7576
rect 3570 7520 3575 7576
rect 0 7518 3575 7520
rect 0 7428 800 7518
rect 3509 7515 3575 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6748 800 6838
rect 4061 6835 4127 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 47945 6218 48011 6221
rect 49200 6218 50000 6308
rect 47945 6216 50000 6218
rect 47945 6160 47950 6216
rect 48006 6160 50000 6216
rect 47945 6158 50000 6160
rect 47945 6155 48011 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 23013 4042 23079 4045
rect 46657 4042 46723 4045
rect 23013 4040 46723 4042
rect 23013 3984 23018 4040
rect 23074 3984 46662 4040
rect 46718 3984 46723 4040
rect 49200 4028 50000 4118
rect 23013 3982 46723 3984
rect 23013 3979 23079 3982
rect 46657 3979 46723 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 18689 3770 18755 3773
rect 20897 3770 20963 3773
rect 18689 3768 20963 3770
rect 18689 3712 18694 3768
rect 18750 3712 20902 3768
rect 20958 3712 20963 3768
rect 18689 3710 20963 3712
rect 18689 3707 18755 3710
rect 20897 3707 20963 3710
rect 0 3498 800 3588
rect 20110 3572 20116 3636
rect 20180 3634 20186 3636
rect 27613 3634 27679 3637
rect 20180 3632 27679 3634
rect 20180 3576 27618 3632
rect 27674 3576 27679 3632
rect 20180 3574 27679 3576
rect 20180 3572 20186 3574
rect 27613 3571 27679 3574
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3348 800 3438
rect 4061 3435 4127 3438
rect 17401 3498 17467 3501
rect 45829 3498 45895 3501
rect 17401 3496 45895 3498
rect 17401 3440 17406 3496
rect 17462 3440 45834 3496
rect 45890 3440 45895 3496
rect 17401 3438 45895 3440
rect 17401 3435 17467 3438
rect 45829 3435 45895 3438
rect 47761 3498 47827 3501
rect 49200 3498 50000 3588
rect 47761 3496 50000 3498
rect 47761 3440 47766 3496
rect 47822 3440 50000 3496
rect 47761 3438 50000 3440
rect 47761 3435 47827 3438
rect 20069 3362 20135 3365
rect 24669 3362 24735 3365
rect 25037 3362 25103 3365
rect 20069 3360 25103 3362
rect 20069 3304 20074 3360
rect 20130 3304 24674 3360
rect 24730 3304 25042 3360
rect 25098 3304 25103 3360
rect 49200 3348 50000 3438
rect 20069 3302 25103 3304
rect 20069 3299 20135 3302
rect 24669 3299 24735 3302
rect 25037 3299 25103 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 19241 2954 19307 2957
rect 20713 2954 20779 2957
rect 19241 2952 20779 2954
rect 0 2668 800 2908
rect 19241 2896 19246 2952
rect 19302 2896 20718 2952
rect 20774 2896 20779 2952
rect 19241 2894 20779 2896
rect 19241 2891 19307 2894
rect 20713 2891 20779 2894
rect 24117 2954 24183 2957
rect 27613 2954 27679 2957
rect 24117 2952 27679 2954
rect 24117 2896 24122 2952
rect 24178 2896 27618 2952
rect 27674 2896 27679 2952
rect 24117 2894 27679 2896
rect 24117 2891 24183 2894
rect 27613 2891 27679 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3233 1458 3299 1461
rect 0 1456 3299 1458
rect 0 1400 3238 1456
rect 3294 1400 3299 1456
rect 0 1398 3299 1400
rect 0 1308 800 1398
rect 3233 1395 3299 1398
rect 46841 1458 46907 1461
rect 49200 1458 50000 1548
rect 46841 1456 50000 1458
rect 46841 1400 46846 1456
rect 46902 1400 50000 1456
rect 46841 1398 50000 1400
rect 46841 1395 46907 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 48037 778 48103 781
rect 49200 778 50000 868
rect 48037 776 50000 778
rect 48037 720 48042 776
rect 48098 720 50000 776
rect 48037 718 50000 720
rect 48037 715 48103 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 20116 46956 20180 47020
rect 27476 46820 27540 46884
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 27476 24108 27540 24172
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 20116 3572 20180 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 20115 47020 20181 47021
rect 20115 46956 20116 47020
rect 20180 46956 20181 47020
rect 20115 46955 20181 46956
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 20118 3637 20178 46955
rect 27475 46884 27541 46885
rect 27475 46820 27476 46884
rect 27540 46820 27541 46884
rect 27475 46819 27541 46820
rect 27478 24173 27538 46819
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 27475 24172 27541 24173
rect 27475 24108 27476 24172
rect 27540 24108 27541 24172
rect 27475 24107 27541 24108
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 20115 3636 20181 3637
rect 20115 3572 20116 3636
rect 20180 3572 20181 3636
rect 20115 3571 20181 3572
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform -1 0 44988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 35420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 40848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 38640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_206
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_317
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_324
timestamp 1644511149
transform 1 0 30912 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1644511149
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_88
timestamp 1644511149
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_99
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1644511149
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1644511149
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_179
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_191
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_228
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_234
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_256
timestamp 1644511149
transform 1 0 24656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_264
timestamp 1644511149
transform 1 0 25392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1644511149
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_306
timestamp 1644511149
transform 1 0 29256 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1644511149
transform 1 0 30360 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 1644511149
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_366
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_413
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_422
timestamp 1644511149
transform 1 0 39928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_426
timestamp 1644511149
transform 1 0 40296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_435
timestamp 1644511149
transform 1 0 41124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_442
timestamp 1644511149
transform 1 0 41768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_60
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1644511149
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_116
timestamp 1644511149
transform 1 0 11776 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_162
timestamp 1644511149
transform 1 0 16008 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_171
timestamp 1644511149
transform 1 0 16836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1644511149
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_216
timestamp 1644511149
transform 1 0 20976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1644511149
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_266
timestamp 1644511149
transform 1 0 25576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_278
timestamp 1644511149
transform 1 0 26680 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_286
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_294
timestamp 1644511149
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1644511149
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1644511149
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_428
timestamp 1644511149
transform 1 0 40480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1644511149
transform 1 0 42780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_460
timestamp 1644511149
transform 1 0 43424 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_99
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_122
timestamp 1644511149
transform 1 0 12328 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp 1644511149
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1644511149
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1644511149
transform 1 0 15272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_186
timestamp 1644511149
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1644511149
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1644511149
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_234
timestamp 1644511149
transform 1 0 22632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_238
timestamp 1644511149
transform 1 0 23000 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_247
timestamp 1644511149
transform 1 0 23828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_259
timestamp 1644511149
transform 1 0 24932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_271
timestamp 1644511149
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_285
timestamp 1644511149
transform 1 0 27324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_299
timestamp 1644511149
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_323
timestamp 1644511149
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_406
timestamp 1644511149
transform 1 0 38456 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_412
timestamp 1644511149
transform 1 0 39008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_416
timestamp 1644511149
transform 1 0 39376 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_425
timestamp 1644511149
transform 1 0 40204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_432
timestamp 1644511149
transform 1 0 40848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_439
timestamp 1644511149
transform 1 0 41492 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_452
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_464
timestamp 1644511149
transform 1 0 43792 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_476
timestamp 1644511149
transform 1 0 44896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_484
timestamp 1644511149
transform 1 0 45632 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_499
timestamp 1644511149
transform 1 0 47012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1644511149
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_88
timestamp 1644511149
transform 1 0 9200 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_100
timestamp 1644511149
transform 1 0 10304 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_112
timestamp 1644511149
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_124
timestamp 1644511149
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_157
timestamp 1644511149
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1644511149
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1644511149
transform 1 0 16560 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1644511149
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_227
timestamp 1644511149
transform 1 0 21988 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_231
timestamp 1644511149
transform 1 0 22356 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_235
timestamp 1644511149
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1644511149
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1644511149
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_442
timestamp 1644511149
transform 1 0 41768 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_454
timestamp 1644511149
transform 1 0 42872 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_466
timestamp 1644511149
transform 1 0 43976 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_474
timestamp 1644511149
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_410
timestamp 1644511149
transform 1 0 38824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_418
timestamp 1644511149
transform 1 0 39560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_422
timestamp 1644511149
transform 1 0 39928 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_434
timestamp 1644511149
transform 1 0 41032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1644511149
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_429
timestamp 1644511149
transform 1 0 40572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_438
timestamp 1644511149
transform 1 0 41400 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_450
timestamp 1644511149
transform 1 0 42504 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_462
timestamp 1644511149
transform 1 0 43608 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1644511149
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_435
timestamp 1644511149
transform 1 0 41124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1644511149
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_462
timestamp 1644511149
transform 1 0 43608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_474
timestamp 1644511149
transform 1 0 44712 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_486
timestamp 1644511149
transform 1 0 45816 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_498
timestamp 1644511149
transform 1 0 46920 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_429
timestamp 1644511149
transform 1 0 40572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_434
timestamp 1644511149
transform 1 0 41032 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_449
timestamp 1644511149
transform 1 0 42412 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_461
timestamp 1644511149
transform 1 0 43516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_473
timestamp 1644511149
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_481
timestamp 1644511149
transform 1 0 45356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_495
timestamp 1644511149
transform 1 0 46644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_482
timestamp 1644511149
transform 1 0 45448 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_499
timestamp 1644511149
transform 1 0 47012 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_511
timestamp 1644511149
transform 1 0 48116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_515
timestamp 1644511149
transform 1 0 48484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_477
timestamp 1644511149
transform 1 0 44988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_505
timestamp 1644511149
transform 1 0 47564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_253
timestamp 1644511149
transform 1 0 24380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1644511149
transform 1 0 24748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1644511149
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1644511149
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1644511149
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_274
timestamp 1644511149
transform 1 0 26312 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_286
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1644511149
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1644511149
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_507
timestamp 1644511149
transform 1 0 47748 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_515
timestamp 1644511149
transform 1 0 48484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1644511149
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_259
timestamp 1644511149
transform 1 0 24932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_271
timestamp 1644511149
transform 1 0 26036 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_283
timestamp 1644511149
transform 1 0 27140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_295
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_466
timestamp 1644511149
transform 1 0 43976 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1644511149
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1644511149
transform 1 0 23460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1644511149
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1644511149
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_285
timestamp 1644511149
transform 1 0 27324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_297
timestamp 1644511149
transform 1 0 28428 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_309
timestamp 1644511149
transform 1 0 29532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_321
timestamp 1644511149
transform 1 0 30636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1644511149
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_483
timestamp 1644511149
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_495
timestamp 1644511149
transform 1 0 46644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_204
timestamp 1644511149
transform 1 0 19872 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_216
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_224
timestamp 1644511149
transform 1 0 21712 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1644511149
transform 1 0 23184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_260
timestamp 1644511149
transform 1 0 25024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1644511149
transform 1 0 26036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_296
timestamp 1644511149
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_317
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1644511149
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1644511149
transform 1 0 33396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_465
timestamp 1644511149
transform 1 0 43884 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1644511149
transform 1 0 19504 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_207
timestamp 1644511149
transform 1 0 20148 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_215
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1644511149
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1644511149
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_284
timestamp 1644511149
transform 1 0 27232 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_296
timestamp 1644511149
transform 1 0 28336 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1644511149
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_307
timestamp 1644511149
transform 1 0 29348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_319
timestamp 1644511149
transform 1 0 30452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_327
timestamp 1644511149
transform 1 0 31188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_342
timestamp 1644511149
transform 1 0 32568 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_354
timestamp 1644511149
transform 1 0 33672 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_366
timestamp 1644511149
transform 1 0 34776 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_378
timestamp 1644511149
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1644511149
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_465
timestamp 1644511149
transform 1 0 43884 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_487
timestamp 1644511149
transform 1 0 45908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_499
timestamp 1644511149
transform 1 0 47012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_156
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_179
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1644511149
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_212
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_239
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_261
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_270
timestamp 1644511149
transform 1 0 25944 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_282
timestamp 1644511149
transform 1 0 27048 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_291
timestamp 1644511149
transform 1 0 27876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_302
timestamp 1644511149
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_322
timestamp 1644511149
transform 1 0 30728 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_334
timestamp 1644511149
transform 1 0 31832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_338
timestamp 1644511149
transform 1 0 32200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1644511149
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_486
timestamp 1644511149
transform 1 0 45816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_490
timestamp 1644511149
transform 1 0 46184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1644511149
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_155
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_172
timestamp 1644511149
transform 1 0 16928 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1644511149
transform 1 0 18032 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1644511149
transform 1 0 18400 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1644511149
transform 1 0 20332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1644511149
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_228
timestamp 1644511149
transform 1 0 22080 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_240
timestamp 1644511149
transform 1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_264
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_270
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1644511149
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_290
timestamp 1644511149
transform 1 0 27784 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_296
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_304
timestamp 1644511149
transform 1 0 29072 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_313
timestamp 1644511149
transform 1 0 29900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_320
timestamp 1644511149
transform 1 0 30544 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_457
timestamp 1644511149
transform 1 0 43148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_498
timestamp 1644511149
transform 1 0 46920 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_151
timestamp 1644511149
transform 1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_175
timestamp 1644511149
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1644511149
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_217
timestamp 1644511149
transform 1 0 21068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_225
timestamp 1644511149
transform 1 0 21804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1644511149
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1644511149
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1644511149
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_256
timestamp 1644511149
transform 1 0 24656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_281
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_293
timestamp 1644511149
transform 1 0 28060 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1644511149
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_322
timestamp 1644511149
transform 1 0 30728 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_329
timestamp 1644511149
transform 1 0 31372 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_341
timestamp 1644511149
transform 1 0 32476 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_353
timestamp 1644511149
transform 1 0 33580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1644511149
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_378
timestamp 1644511149
transform 1 0 35880 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_382
timestamp 1644511149
transform 1 0 36248 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_394
timestamp 1644511149
transform 1 0 37352 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_406
timestamp 1644511149
transform 1 0 38456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1644511149
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_463
timestamp 1644511149
transform 1 0 43700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_485
timestamp 1644511149
transform 1 0 45724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1644511149
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_120
timestamp 1644511149
transform 1 0 12144 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_126
timestamp 1644511149
transform 1 0 12696 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_134
timestamp 1644511149
transform 1 0 13432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1644511149
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_151
timestamp 1644511149
transform 1 0 14996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1644511149
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1644511149
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_177
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_199
timestamp 1644511149
transform 1 0 19412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_211
timestamp 1644511149
transform 1 0 20516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_248
timestamp 1644511149
transform 1 0 23920 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_264
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1644511149
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_301
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_306
timestamp 1644511149
transform 1 0 29256 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_310
timestamp 1644511149
transform 1 0 29624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_343
timestamp 1644511149
transform 1 0 32660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_365
timestamp 1644511149
transform 1 0 34684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_375
timestamp 1644511149
transform 1 0 35604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1644511149
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_444
timestamp 1644511149
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_470
timestamp 1644511149
transform 1 0 44344 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_490
timestamp 1644511149
transform 1 0 46184 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_496
timestamp 1644511149
transform 1 0 46736 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1644511149
transform 1 0 15732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1644511149
transform 1 0 16376 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_178
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_182
timestamp 1644511149
transform 1 0 17848 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1644511149
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_215
timestamp 1644511149
transform 1 0 20884 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_223
timestamp 1644511149
transform 1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_272
timestamp 1644511149
transform 1 0 26128 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_278
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_285
timestamp 1644511149
transform 1 0 27324 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_314
timestamp 1644511149
transform 1 0 29992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_323
timestamp 1644511149
transform 1 0 30820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_336
timestamp 1644511149
transform 1 0 32016 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_346
timestamp 1644511149
transform 1 0 32936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_353
timestamp 1644511149
transform 1 0 33580 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1644511149
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_386
timestamp 1644511149
transform 1 0 36616 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_398
timestamp 1644511149
transform 1 0 37720 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_410
timestamp 1644511149
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1644511149
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1644511149
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_151
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_173
timestamp 1644511149
transform 1 0 17020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_185
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_196
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_209
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_230
timestamp 1644511149
transform 1 0 22264 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_234
timestamp 1644511149
transform 1 0 22632 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_242
timestamp 1644511149
transform 1 0 23368 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 1644511149
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1644511149
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_346
timestamp 1644511149
transform 1 0 32936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_371
timestamp 1644511149
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1644511149
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_458
timestamp 1644511149
transform 1 0 43240 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_464
timestamp 1644511149
transform 1 0 43792 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_478
timestamp 1644511149
transform 1 0 45080 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_482
timestamp 1644511149
transform 1 0 45448 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_486
timestamp 1644511149
transform 1 0 45816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_493
timestamp 1644511149
transform 1 0 46460 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_113
timestamp 1644511149
transform 1 0 11500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_118
timestamp 1644511149
transform 1 0 11960 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_125
timestamp 1644511149
transform 1 0 12604 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_144
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_152
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_160
timestamp 1644511149
transform 1 0 15824 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_203
timestamp 1644511149
transform 1 0 19780 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_238
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1644511149
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1644511149
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_281
timestamp 1644511149
transform 1 0 26956 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_293
timestamp 1644511149
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1644511149
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_337
timestamp 1644511149
transform 1 0 32108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_368
timestamp 1644511149
transform 1 0 34960 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_380
timestamp 1644511149
transform 1 0 36064 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_392
timestamp 1644511149
transform 1 0 37168 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_404
timestamp 1644511149
transform 1 0 38272 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1644511149
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_454
timestamp 1644511149
transform 1 0 42872 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_467
timestamp 1644511149
transform 1 0 44068 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_483
timestamp 1644511149
transform 1 0 45540 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_487
timestamp 1644511149
transform 1 0 45908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_141
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_153
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_157
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1644511149
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1644511149
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_182
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_190
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_213
timestamp 1644511149
transform 1 0 20700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1644511149
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_229
timestamp 1644511149
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1644511149
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_244
timestamp 1644511149
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_251
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_284
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_288
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1644511149
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_319
timestamp 1644511149
transform 1 0 30452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_327
timestamp 1644511149
transform 1 0 31188 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 1644511149
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_360
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1644511149
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_463
timestamp 1644511149
transform 1 0 43700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_105
timestamp 1644511149
transform 1 0 10764 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1644511149
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_152
timestamp 1644511149
transform 1 0 15088 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_158
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_162
timestamp 1644511149
transform 1 0 16008 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_201
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1644511149
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1644511149
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_259
timestamp 1644511149
transform 1 0 24932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_263
timestamp 1644511149
transform 1 0 25300 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_271
timestamp 1644511149
transform 1 0 26036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_284
timestamp 1644511149
transform 1 0 27232 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1644511149
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_313
timestamp 1644511149
transform 1 0 29900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_325
timestamp 1644511149
transform 1 0 31004 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_380
timestamp 1644511149
transform 1 0 36064 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_404
timestamp 1644511149
transform 1 0 38272 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1644511149
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_448
timestamp 1644511149
transform 1 0 42320 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_459
timestamp 1644511149
transform 1 0 43332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_466
timestamp 1644511149
transform 1 0 43976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1644511149
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_480
timestamp 1644511149
transform 1 0 45264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1644511149
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_120
timestamp 1644511149
transform 1 0 12144 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_128
timestamp 1644511149
transform 1 0 12880 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_132
timestamp 1644511149
transform 1 0 13248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_140
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1644511149
transform 1 0 17296 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_180
timestamp 1644511149
transform 1 0 17664 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_185
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1644511149
transform 1 0 19136 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1644511149
transform 1 0 20240 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_233
timestamp 1644511149
transform 1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_245
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1644511149
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_291
timestamp 1644511149
transform 1 0 27876 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_318
timestamp 1644511149
transform 1 0 30360 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1644511149
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_347
timestamp 1644511149
transform 1 0 33028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_351
timestamp 1644511149
transform 1 0 33396 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_380
timestamp 1644511149
transform 1 0 36064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_384
timestamp 1644511149
transform 1 0 36432 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1644511149
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_455
timestamp 1644511149
transform 1 0 42964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_463
timestamp 1644511149
transform 1 0 43700 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_467
timestamp 1644511149
transform 1 0 44068 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_471
timestamp 1644511149
transform 1 0 44436 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_475
timestamp 1644511149
transform 1 0 44804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_486
timestamp 1644511149
transform 1 0 45816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_510
timestamp 1644511149
transform 1 0 48024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_174
timestamp 1644511149
transform 1 0 17112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_179
timestamp 1644511149
transform 1 0 17572 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1644511149
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_204
timestamp 1644511149
transform 1 0 19872 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_216
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_228
timestamp 1644511149
transform 1 0 22080 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_256
timestamp 1644511149
transform 1 0 24656 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_283
timestamp 1644511149
transform 1 0 27140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_287
timestamp 1644511149
transform 1 0 27508 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_297
timestamp 1644511149
transform 1 0 28428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_312
timestamp 1644511149
transform 1 0 29808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_344
timestamp 1644511149
transform 1 0 32752 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_358
timestamp 1644511149
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1644511149
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_371
timestamp 1644511149
transform 1 0 35236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_375
timestamp 1644511149
transform 1 0 35604 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_387
timestamp 1644511149
transform 1 0 36708 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_412
timestamp 1644511149
transform 1 0 39008 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_426
timestamp 1644511149
transform 1 0 40296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_452
timestamp 1644511149
transform 1 0 42688 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_464
timestamp 1644511149
transform 1 0 43792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_468
timestamp 1644511149
transform 1 0 44160 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1644511149
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_487
timestamp 1644511149
transform 1 0 45908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_120
timestamp 1644511149
transform 1 0 12144 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_132
timestamp 1644511149
transform 1 0 13248 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_138
timestamp 1644511149
transform 1 0 13800 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_150
timestamp 1644511149
transform 1 0 14904 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_159
timestamp 1644511149
transform 1 0 15732 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_172
timestamp 1644511149
transform 1 0 16928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_207
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_245
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_252
timestamp 1644511149
transform 1 0 24288 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_259
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_267
timestamp 1644511149
transform 1 0 25668 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_272
timestamp 1644511149
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1644511149
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_294
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_306
timestamp 1644511149
transform 1 0 29256 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_318
timestamp 1644511149
transform 1 0 30360 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1644511149
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_340
timestamp 1644511149
transform 1 0 32384 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_352
timestamp 1644511149
transform 1 0 33488 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_360
timestamp 1644511149
transform 1 0 34224 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_371
timestamp 1644511149
transform 1 0 35236 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_383
timestamp 1644511149
transform 1 0 36340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_424
timestamp 1644511149
transform 1 0 40112 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_434
timestamp 1644511149
transform 1 0 41032 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_440
timestamp 1644511149
transform 1 0 41584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1644511149
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_465
timestamp 1644511149
transform 1 0 43884 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_471
timestamp 1644511149
transform 1 0 44436 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_475
timestamp 1644511149
transform 1 0 44804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_511
timestamp 1644511149
transform 1 0 48116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_515
timestamp 1644511149
transform 1 0 48484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_125
timestamp 1644511149
transform 1 0 12604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1644511149
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_159
timestamp 1644511149
transform 1 0 15732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1644511149
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1644511149
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_207
timestamp 1644511149
transform 1 0 20148 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_217
timestamp 1644511149
transform 1 0 21068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_225
timestamp 1644511149
transform 1 0 21804 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_232
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_238
timestamp 1644511149
transform 1 0 23000 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_242
timestamp 1644511149
transform 1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1644511149
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_275
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 1644511149
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_313
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_327
timestamp 1644511149
transform 1 0 31188 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_334
timestamp 1644511149
transform 1 0 31832 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_346
timestamp 1644511149
transform 1 0 32936 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1644511149
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_368
timestamp 1644511149
transform 1 0 34960 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_380
timestamp 1644511149
transform 1 0 36064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_388
timestamp 1644511149
transform 1 0 36800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_394
timestamp 1644511149
transform 1 0 37352 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_406
timestamp 1644511149
transform 1 0 38456 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_416
timestamp 1644511149
transform 1 0 39376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_443
timestamp 1644511149
transform 1 0 41860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_449
timestamp 1644511149
transform 1 0 42412 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_455
timestamp 1644511149
transform 1 0 42964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_462
timestamp 1644511149
transform 1 0 43608 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1644511149
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_507
timestamp 1644511149
transform 1 0 47748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_117
timestamp 1644511149
transform 1 0 11868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 1644511149
transform 1 0 12788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1644511149
transform 1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1644511149
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_153
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_177
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_189
timestamp 1644511149
transform 1 0 18492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_197
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_257
timestamp 1644511149
transform 1 0 24748 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_265
timestamp 1644511149
transform 1 0 25484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_288
timestamp 1644511149
transform 1 0 27600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_321
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_327
timestamp 1644511149
transform 1 0 31188 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_342
timestamp 1644511149
transform 1 0 32568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_350
timestamp 1644511149
transform 1 0 33304 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_374
timestamp 1644511149
transform 1 0 35512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_381
timestamp 1644511149
transform 1 0 36156 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1644511149
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_398
timestamp 1644511149
transform 1 0 37720 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_410
timestamp 1644511149
transform 1 0 38824 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_456
timestamp 1644511149
transform 1 0 43056 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_468
timestamp 1644511149
transform 1 0 44160 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_480
timestamp 1644511149
transform 1 0 45264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_484
timestamp 1644511149
transform 1 0 45632 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_488
timestamp 1644511149
transform 1 0 46000 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_496
timestamp 1644511149
transform 1 0 46736 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_115
timestamp 1644511149
transform 1 0 11684 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_147
timestamp 1644511149
transform 1 0 14628 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_171
timestamp 1644511149
transform 1 0 16836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_175
timestamp 1644511149
transform 1 0 17204 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1644511149
transform 1 0 17664 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_206
timestamp 1644511149
transform 1 0 20056 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_212
timestamp 1644511149
transform 1 0 20608 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_217
timestamp 1644511149
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_225
timestamp 1644511149
transform 1 0 21804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1644511149
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1644511149
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_261
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_266
timestamp 1644511149
transform 1 0 25576 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1644511149
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_312
timestamp 1644511149
transform 1 0 29808 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_318
timestamp 1644511149
transform 1 0 30360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_339
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_350
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_356
timestamp 1644511149
transform 1 0 33856 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_369
timestamp 1644511149
transform 1 0 35052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_391
timestamp 1644511149
transform 1 0 37076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1644511149
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_442
timestamp 1644511149
transform 1 0 41768 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_454
timestamp 1644511149
transform 1 0 42872 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_466
timestamp 1644511149
transform 1 0 43976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_474
timestamp 1644511149
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_120
timestamp 1644511149
transform 1 0 12144 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_145
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1644511149
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1644511149
transform 1 0 16928 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_179
timestamp 1644511149
transform 1 0 17572 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1644511149
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_258
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_264
timestamp 1644511149
transform 1 0 25392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_268
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_291
timestamp 1644511149
transform 1 0 27876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_299
timestamp 1644511149
transform 1 0 28612 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_311
timestamp 1644511149
transform 1 0 29716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_323
timestamp 1644511149
transform 1 0 30820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1644511149
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_348
timestamp 1644511149
transform 1 0 33120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_355
timestamp 1644511149
transform 1 0 33764 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_370
timestamp 1644511149
transform 1 0 35144 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_382
timestamp 1644511149
transform 1 0 36248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1644511149
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_414
timestamp 1644511149
transform 1 0 39192 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_422
timestamp 1644511149
transform 1 0 39928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_426
timestamp 1644511149
transform 1 0 40296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_438
timestamp 1644511149
transform 1 0 41400 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1644511149
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1644511149
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_117
timestamp 1644511149
transform 1 0 11868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_128
timestamp 1644511149
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1644511149
transform 1 0 14352 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_156
timestamp 1644511149
transform 1 0 15456 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_185
timestamp 1644511149
transform 1 0 18124 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_201
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_215
timestamp 1644511149
transform 1 0 20884 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_226
timestamp 1644511149
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_238
timestamp 1644511149
transform 1 0 23000 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_312
timestamp 1644511149
transform 1 0 29808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_324
timestamp 1644511149
transform 1 0 30912 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_336
timestamp 1644511149
transform 1 0 32016 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1644511149
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_395
timestamp 1644511149
transform 1 0 37444 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_402
timestamp 1644511149
transform 1 0 38088 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_414
timestamp 1644511149
transform 1 0 39192 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_443
timestamp 1644511149
transform 1 0 41860 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_455
timestamp 1644511149
transform 1 0 42964 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_467
timestamp 1644511149
transform 1 0 44068 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_508
timestamp 1644511149
transform 1 0 47840 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_126
timestamp 1644511149
transform 1 0 12696 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_138
timestamp 1644511149
transform 1 0 13800 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_150
timestamp 1644511149
transform 1 0 14904 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1644511149
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_190
timestamp 1644511149
transform 1 0 18584 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_196
timestamp 1644511149
transform 1 0 19136 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_200
timestamp 1644511149
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_209
timestamp 1644511149
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1644511149
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_264
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_316
timestamp 1644511149
transform 1 0 30176 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1644511149
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_357
timestamp 1644511149
transform 1 0 33948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_368
timestamp 1644511149
transform 1 0 34960 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_374
timestamp 1644511149
transform 1 0 35512 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_378
timestamp 1644511149
transform 1 0 35880 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1644511149
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_479
timestamp 1644511149
transform 1 0 45172 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_491
timestamp 1644511149
transform 1 0 46276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_170
timestamp 1644511149
transform 1 0 16744 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_182
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_188
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_217
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_229
timestamp 1644511149
transform 1 0 22172 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_237
timestamp 1644511149
transform 1 0 22908 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_269
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_279
timestamp 1644511149
transform 1 0 26772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_283
timestamp 1644511149
transform 1 0 27140 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1644511149
transform 1 0 27600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_295
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_316
timestamp 1644511149
transform 1 0 30176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_328
timestamp 1644511149
transform 1 0 31280 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_340
timestamp 1644511149
transform 1 0 32384 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_349
timestamp 1644511149
transform 1 0 33212 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_355
timestamp 1644511149
transform 1 0 33764 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_385
timestamp 1644511149
transform 1 0 36524 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_393
timestamp 1644511149
transform 1 0 37260 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1644511149
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_153
timestamp 1644511149
transform 1 0 15180 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_157
timestamp 1644511149
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_195
timestamp 1644511149
transform 1 0 19044 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_201
timestamp 1644511149
transform 1 0 19596 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_208
timestamp 1644511149
transform 1 0 20240 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_230
timestamp 1644511149
transform 1 0 22264 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_239
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_250
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_259
timestamp 1644511149
transform 1 0 24932 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1644511149
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1644511149
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_311
timestamp 1644511149
transform 1 0 29716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_315
timestamp 1644511149
transform 1 0 30084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_322
timestamp 1644511149
transform 1 0 30728 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_359
timestamp 1644511149
transform 1 0 34132 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_368
timestamp 1644511149
transform 1 0 34960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_375
timestamp 1644511149
transform 1 0 35604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1644511149
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_149
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_173
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_185
timestamp 1644511149
transform 1 0 18124 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1644511149
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_203
timestamp 1644511149
transform 1 0 19780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_220
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_232
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_244
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1644511149
transform 1 0 24840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_270
timestamp 1644511149
transform 1 0 25944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_278
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_296
timestamp 1644511149
transform 1 0 28336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_343
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_349
timestamp 1644511149
transform 1 0 33212 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_353
timestamp 1644511149
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1644511149
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_177
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_187
timestamp 1644511149
transform 1 0 18308 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_199
timestamp 1644511149
transform 1 0 19412 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_211
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_230
timestamp 1644511149
transform 1 0 22264 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_242
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_248
timestamp 1644511149
transform 1 0 23920 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_256
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_268
timestamp 1644511149
transform 1 0 25760 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_290
timestamp 1644511149
transform 1 0 27784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_298
timestamp 1644511149
transform 1 0 28520 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_313
timestamp 1644511149
transform 1 0 29900 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_324
timestamp 1644511149
transform 1 0 30912 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_356
timestamp 1644511149
transform 1 0 33856 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_367
timestamp 1644511149
transform 1 0 34868 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_374
timestamp 1644511149
transform 1 0 35512 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_386
timestamp 1644511149
transform 1 0 36616 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1644511149
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_182
timestamp 1644511149
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1644511149
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_217
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_230
timestamp 1644511149
transform 1 0 22264 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1644511149
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_317
timestamp 1644511149
transform 1 0 30268 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_327
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_339
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_343
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_347
timestamp 1644511149
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1644511149
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_385
timestamp 1644511149
transform 1 0 36524 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_397
timestamp 1644511149
transform 1 0 37628 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_409
timestamp 1644511149
transform 1 0 38732 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_417
timestamp 1644511149
transform 1 0 39468 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_507
timestamp 1644511149
transform 1 0 47748 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_515
timestamp 1644511149
transform 1 0 48484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_177
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_189
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_197
timestamp 1644511149
transform 1 0 19228 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_254
timestamp 1644511149
transform 1 0 24472 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_264
timestamp 1644511149
transform 1 0 25392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_284
timestamp 1644511149
transform 1 0 27232 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_296
timestamp 1644511149
transform 1 0 28336 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_304
timestamp 1644511149
transform 1 0 29072 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_316
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_328
timestamp 1644511149
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_364
timestamp 1644511149
transform 1 0 34592 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_376
timestamp 1644511149
transform 1 0 35696 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_161
timestamp 1644511149
transform 1 0 15916 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_183
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_190
timestamp 1644511149
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_205
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_217
timestamp 1644511149
transform 1 0 21068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_228
timestamp 1644511149
transform 1 0 22080 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_236
timestamp 1644511149
transform 1 0 22816 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_240
timestamp 1644511149
transform 1 0 23184 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_263
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_267
timestamp 1644511149
transform 1 0 25668 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_316
timestamp 1644511149
transform 1 0 30176 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_323
timestamp 1644511149
transform 1 0 30820 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_335
timestamp 1644511149
transform 1 0 31924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_347
timestamp 1644511149
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1644511149
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_368
timestamp 1644511149
transform 1 0 34960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_380
timestamp 1644511149
transform 1 0 36064 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_392
timestamp 1644511149
transform 1 0 37168 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_404
timestamp 1644511149
transform 1 0 38272 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_416
timestamp 1644511149
transform 1 0 39376 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_157
timestamp 1644511149
transform 1 0 15548 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1644511149
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_180
timestamp 1644511149
transform 1 0 17664 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1644511149
transform 1 0 19136 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_208
timestamp 1644511149
transform 1 0 20240 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_212
timestamp 1644511149
transform 1 0 20608 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_245
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_263
timestamp 1644511149
transform 1 0 25300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_285
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_303
timestamp 1644511149
transform 1 0 28980 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_327
timestamp 1644511149
transform 1 0 31188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_348
timestamp 1644511149
transform 1 0 33120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_360
timestamp 1644511149
transform 1 0 34224 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_382
timestamp 1644511149
transform 1 0 36248 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1644511149
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_163
timestamp 1644511149
transform 1 0 16100 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_171
timestamp 1644511149
transform 1 0 16836 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_178
timestamp 1644511149
transform 1 0 17480 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_185
timestamp 1644511149
transform 1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1644511149
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_200
timestamp 1644511149
transform 1 0 19504 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_208
timestamp 1644511149
transform 1 0 20240 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_218
timestamp 1644511149
transform 1 0 21160 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_230
timestamp 1644511149
transform 1 0 22264 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_274
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_281
timestamp 1644511149
transform 1 0 26956 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_288
timestamp 1644511149
transform 1 0 27600 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_313
timestamp 1644511149
transform 1 0 29900 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_319
timestamp 1644511149
transform 1 0 30452 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_327
timestamp 1644511149
transform 1 0 31188 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_355
timestamp 1644511149
transform 1 0 33764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_26
timestamp 1644511149
transform 1 0 3496 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_38
timestamp 1644511149
transform 1 0 4600 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1644511149
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_150
timestamp 1644511149
transform 1 0 14904 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_157
timestamp 1644511149
transform 1 0 15548 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_165
timestamp 1644511149
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_177
timestamp 1644511149
transform 1 0 17388 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_201
timestamp 1644511149
transform 1 0 19596 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_209
timestamp 1644511149
transform 1 0 20332 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1644511149
transform 1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_236
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_247
timestamp 1644511149
transform 1 0 23828 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1644511149
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_264
timestamp 1644511149
transform 1 0 25392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1644511149
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_285
timestamp 1644511149
transform 1 0 27324 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_298
timestamp 1644511149
transform 1 0 28520 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_307
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_346
timestamp 1644511149
transform 1 0 32936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_358
timestamp 1644511149
transform 1 0 34040 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_370
timestamp 1644511149
transform 1 0 35144 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1644511149
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1644511149
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_50
timestamp 1644511149
transform 1 0 5704 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_62
timestamp 1644511149
transform 1 0 6808 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_74
timestamp 1644511149
transform 1 0 7912 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1644511149
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_161
timestamp 1644511149
transform 1 0 15916 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_170
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_178
timestamp 1644511149
transform 1 0 17480 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1644511149
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_205
timestamp 1644511149
transform 1 0 19964 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_226
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_232
timestamp 1644511149
transform 1 0 22448 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_236
timestamp 1644511149
transform 1 0 22816 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1644511149
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_262
timestamp 1644511149
transform 1 0 25208 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_272
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_280
timestamp 1644511149
transform 1 0 26864 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_318
timestamp 1644511149
transform 1 0 30360 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_325
timestamp 1644511149
transform 1 0 31004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_342
timestamp 1644511149
transform 1 0 32568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1644511149
transform 1 0 33212 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_361
timestamp 1644511149
transform 1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_506
timestamp 1644511149
transform 1 0 47656 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_514
timestamp 1644511149
transform 1 0 48392 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_8
timestamp 1644511149
transform 1 0 1840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_33
timestamp 1644511149
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1644511149
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1644511149
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_157
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_182
timestamp 1644511149
transform 1 0 17848 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_194
timestamp 1644511149
transform 1 0 18952 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_206
timestamp 1644511149
transform 1 0 20056 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_218
timestamp 1644511149
transform 1 0 21160 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_248
timestamp 1644511149
transform 1 0 23920 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1644511149
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_290
timestamp 1644511149
transform 1 0 27784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_298
timestamp 1644511149
transform 1 0 28520 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_311
timestamp 1644511149
transform 1 0 29716 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_325
timestamp 1644511149
transform 1 0 31004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1644511149
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_357
timestamp 1644511149
transform 1 0 33948 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_369
timestamp 1644511149
transform 1 0 35052 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_381
timestamp 1644511149
transform 1 0 36156 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_389
timestamp 1644511149
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1644511149
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_14
timestamp 1644511149
transform 1 0 2392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1644511149
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_151
timestamp 1644511149
transform 1 0 14996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1644511149
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_169
timestamp 1644511149
transform 1 0 16652 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_173
timestamp 1644511149
transform 1 0 17020 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_180
timestamp 1644511149
transform 1 0 17664 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1644511149
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_202
timestamp 1644511149
transform 1 0 19688 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_214
timestamp 1644511149
transform 1 0 20792 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_219
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_223
timestamp 1644511149
transform 1 0 21620 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_228
timestamp 1644511149
transform 1 0 22080 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_236
timestamp 1644511149
transform 1 0 22816 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_240
timestamp 1644511149
transform 1 0 23184 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_260
timestamp 1644511149
transform 1 0 25024 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_284
timestamp 1644511149
transform 1 0 27232 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_292
timestamp 1644511149
transform 1 0 27968 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_297
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1644511149
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_322
timestamp 1644511149
transform 1 0 30728 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_332
timestamp 1644511149
transform 1 0 31648 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_341
timestamp 1644511149
transform 1 0 32476 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_353
timestamp 1644511149
transform 1 0 33580 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1644511149
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_483
timestamp 1644511149
transform 1 0 45540 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_487
timestamp 1644511149
transform 1 0 45908 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_148
timestamp 1644511149
transform 1 0 14720 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 1644511149
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1644511149
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_189
timestamp 1644511149
transform 1 0 18492 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_215
timestamp 1644511149
transform 1 0 20884 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_235
timestamp 1644511149
transform 1 0 22724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1644511149
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_255
timestamp 1644511149
transform 1 0 24564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_267
timestamp 1644511149
transform 1 0 25668 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_274
timestamp 1644511149
transform 1 0 26312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_288
timestamp 1644511149
transform 1 0 27600 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_296
timestamp 1644511149
transform 1 0 28336 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_304
timestamp 1644511149
transform 1 0 29072 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_316
timestamp 1644511149
transform 1 0 30176 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_328
timestamp 1644511149
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_340
timestamp 1644511149
transform 1 0 32384 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_347
timestamp 1644511149
transform 1 0 33028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_359
timestamp 1644511149
transform 1 0 34132 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_371
timestamp 1644511149
transform 1 0 35236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1644511149
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_493
timestamp 1644511149
transform 1 0 46460 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_511
timestamp 1644511149
transform 1 0 48116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_515
timestamp 1644511149
transform 1 0 48484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_162
timestamp 1644511149
transform 1 0 16008 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_173
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_58_190
timestamp 1644511149
transform 1 0 18584 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_225
timestamp 1644511149
transform 1 0 21804 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_236
timestamp 1644511149
transform 1 0 22816 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_257
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_269
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_284
timestamp 1644511149
transform 1 0 27232 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_296
timestamp 1644511149
transform 1 0 28336 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_319
timestamp 1644511149
transform 1 0 30452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_344
timestamp 1644511149
transform 1 0 32752 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_356
timestamp 1644511149
transform 1 0 33856 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_153
timestamp 1644511149
transform 1 0 15180 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_157
timestamp 1644511149
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1644511149
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_197
timestamp 1644511149
transform 1 0 19228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp 1644511149
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_231
timestamp 1644511149
transform 1 0 22356 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_244
timestamp 1644511149
transform 1 0 23552 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_252
timestamp 1644511149
transform 1 0 24288 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_260
timestamp 1644511149
transform 1 0 25024 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_265
timestamp 1644511149
transform 1 0 25484 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1644511149
transform 1 0 27416 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_298
timestamp 1644511149
transform 1 0 28520 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_308
timestamp 1644511149
transform 1 0 29440 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 1644511149
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1644511149
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_163
timestamp 1644511149
transform 1 0 16100 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_175
timestamp 1644511149
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_190
timestamp 1644511149
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_215
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_228
timestamp 1644511149
transform 1 0 22080 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1644511149
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_257
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_261
timestamp 1644511149
transform 1 0 25116 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_287
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_298
timestamp 1644511149
transform 1 0 28520 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1644511149
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_313
timestamp 1644511149
transform 1 0 29900 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_162
timestamp 1644511149
transform 1 0 16008 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_176
timestamp 1644511149
transform 1 0 17296 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_184
timestamp 1644511149
transform 1 0 18032 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_189
timestamp 1644511149
transform 1 0 18492 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_201
timestamp 1644511149
transform 1 0 19596 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_213
timestamp 1644511149
transform 1 0 20700 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_221
timestamp 1644511149
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_233
timestamp 1644511149
transform 1 0 22540 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_241
timestamp 1644511149
transform 1 0 23276 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_253
timestamp 1644511149
transform 1 0 24380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_262
timestamp 1644511149
transform 1 0 25208 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_270
timestamp 1644511149
transform 1 0 25944 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_292
timestamp 1644511149
transform 1 0 27968 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_298
timestamp 1644511149
transform 1 0 28520 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_319
timestamp 1644511149
transform 1 0 30452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_331
timestamp 1644511149
transform 1 0 31556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1644511149
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_147
timestamp 1644511149
transform 1 0 14628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1644511149
transform 1 0 16560 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_180
timestamp 1644511149
transform 1 0 17664 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_204
timestamp 1644511149
transform 1 0 19872 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_216
timestamp 1644511149
transform 1 0 20976 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_228
timestamp 1644511149
transform 1 0 22080 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_240
timestamp 1644511149
transform 1 0 23184 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1644511149
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_262
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_274
timestamp 1644511149
transform 1 0 26312 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_291
timestamp 1644511149
transform 1 0 27876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_303
timestamp 1644511149
transform 1 0 28980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_157
timestamp 1644511149
transform 1 0 15548 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1644511149
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_175
timestamp 1644511149
transform 1 0 17204 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1644511149
transform 1 0 19136 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1644511149
transform 1 0 20240 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_270
timestamp 1644511149
transform 1 0 25944 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1644511149
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_288
timestamp 1644511149
transform 1 0 27600 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_297
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1644511149
transform 1 0 29256 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1644511149
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1644511149
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_211
timestamp 1644511149
transform 1 0 20516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_219
timestamp 1644511149
transform 1 0 21252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_246
timestamp 1644511149
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_256
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_260
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_264
timestamp 1644511149
transform 1 0 25392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_268
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_272
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_298
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1644511149
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_465
timestamp 1644511149
transform 1 0 43884 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_471
timestamp 1644511149
transform 1 0 44436 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_199
timestamp 1644511149
transform 1 0 19412 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_228
timestamp 1644511149
transform 1 0 22080 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_240
timestamp 1644511149
transform 1 0 23184 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_247
timestamp 1644511149
transform 1 0 23828 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_255
timestamp 1644511149
transform 1 0 24564 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_289
timestamp 1644511149
transform 1 0 27692 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_481
timestamp 1644511149
transform 1 0 45356 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_493
timestamp 1644511149
transform 1 0 46460 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_499
timestamp 1644511149
transform 1 0 47012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_173
timestamp 1644511149
transform 1 0 17020 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_213
timestamp 1644511149
transform 1 0 20700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_225
timestamp 1644511149
transform 1 0 21804 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_237
timestamp 1644511149
transform 1 0 22908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1644511149
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_449
timestamp 1644511149
transform 1 0 42412 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_459
timestamp 1644511149
transform 1 0 43332 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_472
timestamp 1644511149
transform 1 0 44528 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_486
timestamp 1644511149
transform 1 0 45816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_490
timestamp 1644511149
transform 1 0 46184 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_213
timestamp 1644511149
transform 1 0 20700 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_221
timestamp 1644511149
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_231
timestamp 1644511149
transform 1 0 22356 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_252
timestamp 1644511149
transform 1 0 24288 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_264
timestamp 1644511149
transform 1 0 25392 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_480
timestamp 1644511149
transform 1 0 45264 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_492
timestamp 1644511149
transform 1 0 46368 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_499
timestamp 1644511149
transform 1 0 47012 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_239
timestamp 1644511149
transform 1 0 23092 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_243
timestamp 1644511149
transform 1 0 23460 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_262
timestamp 1644511149
transform 1 0 25208 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_274
timestamp 1644511149
transform 1 0 26312 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_286
timestamp 1644511149
transform 1 0 27416 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_298
timestamp 1644511149
transform 1 0 28520 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_306
timestamp 1644511149
transform 1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1644511149
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_493
timestamp 1644511149
transform 1 0 46460 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_498
timestamp 1644511149
transform 1 0 46920 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_296
timestamp 1644511149
transform 1 0 28336 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_407
timestamp 1644511149
transform 1 0 38548 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_411
timestamp 1644511149
transform 1 0 38916 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_428
timestamp 1644511149
transform 1 0 40480 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_440
timestamp 1644511149
transform 1 0 41584 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_14
timestamp 1644511149
transform 1 0 2392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1644511149
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_461
timestamp 1644511149
transform 1 0 43516 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_465
timestamp 1644511149
transform 1 0 43884 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_28
timestamp 1644511149
transform 1 0 3680 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_40
timestamp 1644511149
transform 1 0 4784 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1644511149
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_140
timestamp 1644511149
transform 1 0 13984 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_152
timestamp 1644511149
transform 1 0 15088 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1644511149
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_216
timestamp 1644511149
transform 1 0 20976 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_267
timestamp 1644511149
transform 1 0 25668 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_274
timestamp 1644511149
transform 1 0 26312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_452
timestamp 1644511149
transform 1 0 42688 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_459
timestamp 1644511149
transform 1 0 43332 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_467
timestamp 1644511149
transform 1 0 44068 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_492
timestamp 1644511149
transform 1 0 46368 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_7
timestamp 1644511149
transform 1 0 1748 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1644511149
transform 1 0 2116 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1644511149
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_35
timestamp 1644511149
transform 1 0 4324 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_39
timestamp 1644511149
transform 1 0 4692 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_48
timestamp 1644511149
transform 1 0 5520 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_60
timestamp 1644511149
transform 1 0 6624 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_72
timestamp 1644511149
transform 1 0 7728 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_125
timestamp 1644511149
transform 1 0 12604 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_132
timestamp 1644511149
transform 1 0 13248 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_205
timestamp 1644511149
transform 1 0 19964 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_234
timestamp 1644511149
transform 1 0 22632 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_246
timestamp 1644511149
transform 1 0 23736 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_259
timestamp 1644511149
transform 1 0 24932 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_284
timestamp 1644511149
transform 1 0 27232 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_296
timestamp 1644511149
transform 1 0 28336 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_336
timestamp 1644511149
transform 1 0 32016 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_348
timestamp 1644511149
transform 1 0 33120 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1644511149
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_458
timestamp 1644511149
transform 1 0 43240 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_464
timestamp 1644511149
transform 1 0 43792 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_7
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_19
timestamp 1644511149
transform 1 0 2852 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_228
timestamp 1644511149
transform 1 0 22080 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_240
timestamp 1644511149
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_252
timestamp 1644511149
transform 1 0 24288 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_358
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_370
timestamp 1644511149
transform 1 0 35144 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_382
timestamp 1644511149
transform 1 0 36248 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_390
timestamp 1644511149
transform 1 0 36984 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1644511149
transform 1 0 6900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1644511149
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_145
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_203
timestamp 1644511149
transform 1 0 19780 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_211
timestamp 1644511149
transform 1 0 20516 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_228
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_240
timestamp 1644511149
transform 1 0 23184 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_259
timestamp 1644511149
transform 1 0 24932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_271
timestamp 1644511149
transform 1 0 26036 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_279
timestamp 1644511149
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_323
timestamp 1644511149
transform 1 0 30820 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_328
timestamp 1644511149
transform 1 0 31280 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_444
timestamp 1644511149
transform 1 0 41952 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0597_
timestamp 1644511149
transform 1 0 32568 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29716 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29256 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0601_
timestamp 1644511149
transform 1 0 32016 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0603_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0604_
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0605_
timestamp 1644511149
transform 1 0 18032 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0606_
timestamp 1644511149
transform 1 0 26956 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0607_
timestamp 1644511149
transform 1 0 23276 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0608_
timestamp 1644511149
transform 1 0 23092 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0609_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0611_
timestamp 1644511149
transform 1 0 20608 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0612_
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0615_
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1644511149
transform 1 0 28060 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32660 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0618_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0620_
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0621_
timestamp 1644511149
transform 1 0 19320 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0622_
timestamp 1644511149
transform 1 0 25944 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0623_
timestamp 1644511149
transform 1 0 24656 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0624_
timestamp 1644511149
transform 1 0 25300 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0625_
timestamp 1644511149
transform 1 0 14536 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0626_
timestamp 1644511149
transform 1 0 19504 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0627_
timestamp 1644511149
transform 1 0 20424 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0628_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32660 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0630_
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34224 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1644511149
transform 1 0 33304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0633_
timestamp 1644511149
transform 1 0 34500 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0634_
timestamp 1644511149
transform 1 0 32568 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1644511149
transform 1 0 35604 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33856 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35328 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1644511149
transform 1 0 35880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0639_
timestamp 1644511149
transform 1 0 34500 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0641_
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0642_
timestamp 1644511149
transform 1 0 32936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0643_
timestamp 1644511149
transform 1 0 33488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0644_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0646_
timestamp 1644511149
transform 1 0 30912 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1644511149
transform 1 0 31556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0648_
timestamp 1644511149
transform 1 0 31280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0651_
timestamp 1644511149
transform 1 0 27232 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1644511149
transform 1 0 23092 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1644511149
transform 1 0 20516 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0656_
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0657_
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1644511149
transform 1 0 22172 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0660_
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 1644511149
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 18308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0665_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1644511149
transform 1 0 17112 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0670_
timestamp 1644511149
transform 1 0 12880 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1644511149
transform 1 0 13892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11960 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0674_
timestamp 1644511149
transform 1 0 12328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0677_
timestamp 1644511149
transform 1 0 12052 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1644511149
transform 1 0 16744 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0680_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1644511149
transform 1 0 13156 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0682_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0683_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0684_
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1644511149
transform 1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0687_
timestamp 1644511149
transform 1 0 15364 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0688_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0690_
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0692_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 14352 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0694_
timestamp 1644511149
transform 1 0 12788 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0695_
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1644511149
transform 1 0 21988 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0698_
timestamp 1644511149
transform 1 0 20700 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0701_
timestamp 1644511149
transform 1 0 20700 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0702_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1644511149
transform 1 0 19872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0704_
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0707_
timestamp 1644511149
transform 1 0 20976 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0710_
timestamp 1644511149
transform 1 0 26312 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0711_
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0712_
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0713_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0714_
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0716_
timestamp 1644511149
transform 1 0 24656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0717_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0719_
timestamp 1644511149
transform 1 0 25392 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1644511149
transform 1 0 26036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0721_
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0722_
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 1644511149
transform 1 0 25760 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1644511149
transform 1 0 25208 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0728_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1644511149
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 29624 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0733_
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0735_
timestamp 1644511149
transform 1 0 26772 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0738_
timestamp 1644511149
transform 1 0 27232 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0739_
timestamp 1644511149
transform 1 0 28704 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0740_
timestamp 1644511149
transform 1 0 25024 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0743_
timestamp 1644511149
transform 1 0 22632 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0744_
timestamp 1644511149
transform 1 0 24472 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0746_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0748_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0749_
timestamp 1644511149
transform 1 0 28152 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0750_
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0751_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0752_
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0755_
timestamp 1644511149
transform 1 0 23552 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0756_
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0757_
timestamp 1644511149
transform 1 0 26220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0758_
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0759_
timestamp 1644511149
transform 1 0 19688 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23920 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0761_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0762_
timestamp 1644511149
transform 1 0 19872 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0763_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19872 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _0764_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0765_
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0766_
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0767_
timestamp 1644511149
transform 1 0 24196 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1644511149
transform 1 0 17204 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1644511149
transform 1 0 16376 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0771_
timestamp 1644511149
transform 1 0 23552 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0773_
timestamp 1644511149
transform 1 0 21528 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0774_
timestamp 1644511149
transform 1 0 21620 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0775_
timestamp 1644511149
transform 1 0 22632 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0776_
timestamp 1644511149
transform 1 0 27968 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0777_
timestamp 1644511149
transform 1 0 24932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0778_
timestamp 1644511149
transform 1 0 20516 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0779_
timestamp 1644511149
transform 1 0 20240 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0780_
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1644511149
transform 1 0 20792 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0783_
timestamp 1644511149
transform 1 0 20056 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0784_
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1644511149
transform 1 0 23184 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0786_
timestamp 1644511149
transform 1 0 23920 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0787_
timestamp 1644511149
transform 1 0 21528 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0788_
timestamp 1644511149
transform 1 0 22172 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0789_
timestamp 1644511149
transform 1 0 20332 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0790_
timestamp 1644511149
transform 1 0 22724 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _0791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0792_
timestamp 1644511149
transform 1 0 23276 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1644511149
transform 1 0 23184 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0795_
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1644511149
transform 1 0 28152 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0797_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0798_
timestamp 1644511149
transform 1 0 17112 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0799_
timestamp 1644511149
transform 1 0 20056 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1644511149
transform 1 0 23552 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0801_
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23644 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0803_
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0805_
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0806_
timestamp 1644511149
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0807_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0808_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0809_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0810_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0811_
timestamp 1644511149
transform 1 0 22632 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0812_
timestamp 1644511149
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0813_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0814_
timestamp 1644511149
transform 1 0 27416 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0815_
timestamp 1644511149
transform 1 0 27876 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0816_
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1644511149
transform 1 0 27968 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0818_
timestamp 1644511149
transform 1 0 27232 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0819_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0820_
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1644511149
transform 1 0 26956 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0822_
timestamp 1644511149
transform 1 0 25944 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0823_
timestamp 1644511149
transform 1 0 25760 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0824_
timestamp 1644511149
transform 1 0 25668 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0825_
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0826_
timestamp 1644511149
transform 1 0 25760 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0827_
timestamp 1644511149
transform 1 0 17020 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1644511149
transform 1 0 16192 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0829_
timestamp 1644511149
transform 1 0 30084 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29348 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1644511149
transform 1 0 15640 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0832_
timestamp 1644511149
transform 1 0 17848 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0833_
timestamp 1644511149
transform 1 0 23368 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0834_
timestamp 1644511149
transform 1 0 23184 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0837_
timestamp 1644511149
transform 1 0 17020 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0838_
timestamp 1644511149
transform 1 0 17112 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0839_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0840_
timestamp 1644511149
transform 1 0 15364 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0841_
timestamp 1644511149
transform 1 0 16192 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0842_
timestamp 1644511149
transform 1 0 17204 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0843_
timestamp 1644511149
transform 1 0 17572 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1644511149
transform 1 0 15364 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0845_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1644511149
transform 1 0 15548 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0847_
timestamp 1644511149
transform 1 0 14628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0848_
timestamp 1644511149
transform 1 0 14444 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0849_
timestamp 1644511149
transform 1 0 16376 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0850_
timestamp 1644511149
transform 1 0 15088 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0851_
timestamp 1644511149
transform 1 0 14260 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0852_
timestamp 1644511149
transform 1 0 15272 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0853_
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0854_
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0855_
timestamp 1644511149
transform 1 0 17848 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0856_
timestamp 1644511149
transform 1 0 17756 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0857_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0858_
timestamp 1644511149
transform 1 0 18952 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0859_
timestamp 1644511149
transform 1 0 18216 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0861_
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 1644511149
transform 1 0 30728 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31096 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0864_
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1644511149
transform 1 0 28888 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0866_
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0867_
timestamp 1644511149
transform 1 0 27140 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0868_
timestamp 1644511149
transform 1 0 29900 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0869_
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0870_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0872_
timestamp 1644511149
transform 1 0 29808 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1644511149
transform 1 0 29992 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0874_
timestamp 1644511149
transform 1 0 30544 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0875_
timestamp 1644511149
transform 1 0 29256 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0876_
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0877_
timestamp 1644511149
transform 1 0 30544 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0878_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0879_
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0880_
timestamp 1644511149
transform 1 0 29256 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0881_
timestamp 1644511149
transform 1 0 30176 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1644511149
transform 1 0 28060 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0883_
timestamp 1644511149
transform 1 0 28704 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1644511149
transform 1 0 27968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0887_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0889_
timestamp 1644511149
transform 1 0 36984 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0890_
timestamp 1644511149
transform 1 0 36156 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 43976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 43700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 46736 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 38640 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 25392 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0902_
timestamp 1644511149
transform 1 0 37168 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 12972 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37628 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 45632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 24472 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0914_
timestamp 1644511149
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32476 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 32292 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 35788 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0921_
timestamp 1644511149
transform 1 0 16928 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 15732 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0927_
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 19320 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 15088 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 17572 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 15272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0933_
timestamp 1644511149
transform 1 0 22264 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 31280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 17296 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 37444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0939_
timestamp 1644511149
transform 1 0 32936 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 37812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0945_
timestamp 1644511149
transform 1 0 44068 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0946_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0952_
timestamp 1644511149
transform 1 0 44252 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0958_
timestamp 1644511149
transform 1 0 43700 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 31096 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 44896 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 39192 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0964_
timestamp 1644511149
transform 1 0 42504 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 24656 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 5244 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0970_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44252 0 -1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0976_
timestamp 1644511149
transform 1 0 33856 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0977_
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 11960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 11868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0983_
timestamp 1644511149
transform 1 0 33396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 37168 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 32752 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 23552 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 46736 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0989_
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 43056 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0995_
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 20056 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1001_
timestamp 1644511149
transform 1 0 22172 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1644511149
transform 1 0 27048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1644511149
transform 1 0 27508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform 1 0 33856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45080 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1015_
timestamp 1644511149
transform 1 0 45264 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1016_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1021_
timestamp 1644511149
transform 1 0 45264 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1644511149
transform 1 0 44528 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1023_
timestamp 1644511149
transform 1 0 45172 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1024_
timestamp 1644511149
transform 1 0 40480 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1644511149
transform 1 0 40664 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1026_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1644511149
transform 1 0 39744 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1029_
timestamp 1644511149
transform 1 0 39928 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1644511149
transform 1 0 40204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21712 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _1032_
timestamp 1644511149
transform 1 0 42504 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1644511149
transform 1 0 43332 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1644511149
transform 1 0 42780 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1035_
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1036_
timestamp 1644511149
transform 1 0 43700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1644511149
transform 1 0 45540 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1644511149
transform 1 0 27508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 1644511149
transform 1 0 28428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1040_
timestamp 1644511149
transform 1 0 28336 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1042_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1043_
timestamp 1644511149
transform 1 0 44068 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1044_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1045_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1644511149
transform 1 0 42688 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1047_
timestamp 1644511149
transform 1 0 42688 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42688 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1049_
timestamp 1644511149
transform 1 0 42964 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1644511149
transform 1 0 42412 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1052_
timestamp 1644511149
transform 1 0 42504 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 1644511149
transform 1 0 43608 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1644511149
transform 1 0 43792 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43884 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1056_
timestamp 1644511149
transform 1 0 43424 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1057_
timestamp 1644511149
transform 1 0 43424 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1058_
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1060_
timestamp 1644511149
transform 1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1061_
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1064_
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1065_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 1644511149
transform 1 0 30360 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1644511149
transform 1 0 32200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1644511149
transform 1 0 42320 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1071_
timestamp 1644511149
transform 1 0 38732 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1072_
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1073_
timestamp 1644511149
transform 1 0 32384 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1644511149
transform 1 0 33304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1075_
timestamp 1644511149
transform 1 0 27600 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1644511149
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1077_
timestamp 1644511149
transform 1 0 1840 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1079_
timestamp 1644511149
transform 1 0 45172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1644511149
transform 1 0 45172 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1081_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform 1 0 34960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1083_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1085_
timestamp 1644511149
transform 1 0 40848 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1644511149
transform 1 0 41216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1087_
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1089_
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 31096 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1093_
timestamp 1644511149
transform 1 0 27692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1644511149
transform 1 0 32752 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 30544 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 32936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1099_
timestamp 1644511149
transform 1 0 18768 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 18216 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1644511149
transform 1 0 18308 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 15272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1644511149
transform 1 0 15732 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1644511149
transform 1 0 25668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1644511149
transform 1 0 18308 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 27324 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1111_
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 27784 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1644511149
transform 1 0 28980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1117_
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1644511149
transform 1 0 22632 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1644511149
transform 1 0 20976 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1644511149
transform 1 0 20148 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1644511149
transform 1 0 22908 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1123_
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1644511149
transform 1 0 25484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1129_
timestamp 1644511149
transform 1 0 28612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1130_
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1644511149
transform 1 0 23920 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1132_
timestamp 1644511149
transform 1 0 26772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1133_
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1134_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1135_
timestamp 1644511149
transform 1 0 23552 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1136_
timestamp 1644511149
transform 1 0 20976 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1137_
timestamp 1644511149
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1138_
timestamp 1644511149
transform 1 0 14536 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1644511149
transform 1 0 17848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1140_
timestamp 1644511149
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1141_
timestamp 1644511149
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1143_
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1144_
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1145_
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1146_
timestamp 1644511149
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1147_
timestamp 1644511149
transform 1 0 11776 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1644511149
transform 1 0 11960 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1149_
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1150_
timestamp 1644511149
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1644511149
transform 1 0 15732 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1152_
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1153_
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1154_
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1155_
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1156_
timestamp 1644511149
transform 1 0 27784 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1157_
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1158_
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1159_
timestamp 1644511149
transform 1 0 30820 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1160_
timestamp 1644511149
transform 1 0 33672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1162_
timestamp 1644511149
transform 1 0 33580 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1163_
timestamp 1644511149
transform 1 0 32292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1644511149
transform 1 0 33580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1644511149
transform 1 0 31924 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1644511149
transform 1 0 29348 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1644511149
transform 1 0 26956 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1644511149
transform 1 0 17296 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1644511149
transform 1 0 14260 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1644511149
transform 1 0 14168 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1644511149
transform 1 0 14720 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1644511149
transform 1 0 16100 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1644511149
transform 1 0 22080 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1182_
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1644511149
transform 1 0 25392 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1644511149
transform 1 0 26680 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1644511149
transform 1 0 28612 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1644511149
transform 1 0 21896 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1644511149
transform 1 0 24656 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 1644511149
transform 1 0 19504 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1644511149
transform 1 0 22448 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1644511149
transform 1 0 19964 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1644511149
transform 1 0 19504 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1644511149
transform 1 0 20056 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1644511149
transform 1 0 22632 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1644511149
transform 1 0 17204 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1198_
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1199_
timestamp 1644511149
transform 1 0 28520 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1200_
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1644511149
transform 1 0 23736 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1202_
timestamp 1644511149
transform 1 0 25024 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1203_
timestamp 1644511149
transform 1 0 26404 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1644511149
transform 1 0 24104 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1644511149
transform 1 0 16928 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1210_
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1644511149
transform 1 0 15364 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1644511149
transform 1 0 13156 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1214_
timestamp 1644511149
transform 1 0 11500 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1215_
timestamp 1644511149
transform 1 0 12512 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 1644511149
transform 1 0 11776 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 1644511149
transform 1 0 14996 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1644511149
transform 1 0 16100 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1644511149
transform 1 0 17296 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1222_
timestamp 1644511149
transform 1 0 27968 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1223_
timestamp 1644511149
transform 1 0 30452 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 1644511149
transform 1 0 30912 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 1644511149
transform 1 0 33672 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1226_
timestamp 1644511149
transform 1 0 35144 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 1644511149
transform 1 0 32292 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1230_
timestamp 1644511149
transform 1 0 24472 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1231__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1232__82
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1233__83
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1234__84
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1235__85
timestamp 1644511149
transform 1 0 47472 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1236__86
timestamp 1644511149
transform 1 0 20700 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1237__87
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1238__88
timestamp 1644511149
transform 1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1239__89
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1240__90
timestamp 1644511149
transform 1 0 26036 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1241__91
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1242__92
timestamp 1644511149
transform 1 0 1840 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1243__93
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1244__94
timestamp 1644511149
transform 1 0 4416 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1245__95
timestamp 1644511149
transform 1 0 1564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1246__96
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1247__97
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1248__98
timestamp 1644511149
transform 1 0 46644 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1249__99
timestamp 1644511149
transform 1 0 44528 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1250__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1251__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1252__102
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1253__103
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1254__104
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1255__105
timestamp 1644511149
transform 1 0 46184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1256__106
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1257__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1258__108
timestamp 1644511149
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1259__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1260__110
timestamp 1644511149
transform 1 0 47564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1261__111
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1262__112
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1263__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1264__114
timestamp 1644511149
transform 1 0 45632 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1265__115
timestamp 1644511149
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1266__116
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1267__117
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1268__118
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1269__119
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1270__120
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1271__121
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1272__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1273__123
timestamp 1644511149
transform 1 0 45632 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1274__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1275__125
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1276__126
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1277__127
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1278__128
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1279__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1280__130
timestamp 1644511149
transform 1 0 47472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1281__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1282__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1283__133
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1284__134
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1285__135
timestamp 1644511149
transform 1 0 43608 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 29716 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 43608 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 43976 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 45264 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 46276 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 38548 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 20700 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 25300 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1315_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1316_
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1317_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1318_
timestamp 1644511149
transform 1 0 37076 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1319_
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1320_
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1321_
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1322_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1323_
timestamp 1644511149
transform 1 0 30360 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1324_
timestamp 1644511149
transform 1 0 23552 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1325_
timestamp 1644511149
transform 1 0 16100 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1326_
timestamp 1644511149
transform 1 0 32292 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1327_
timestamp 1644511149
transform 1 0 21160 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1328_
timestamp 1644511149
transform 1 0 20148 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1329_
timestamp 1644511149
transform 1 0 16376 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1330_
timestamp 1644511149
transform 1 0 11684 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1331_
timestamp 1644511149
transform 1 0 17480 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1332_
timestamp 1644511149
transform 1 0 14260 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1333_
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1334_
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1335_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1336_
timestamp 1644511149
transform 1 0 11684 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1337_
timestamp 1644511149
transform 1 0 16192 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1338_
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1339_
timestamp 1644511149
transform 1 0 18768 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1340_
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1341_
timestamp 1644511149
transform 1 0 15088 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1342_
timestamp 1644511149
transform 1 0 26772 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1343_
timestamp 1644511149
transform 1 0 39928 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1344_
timestamp 1644511149
transform 1 0 31188 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1345_
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1346_
timestamp 1644511149
transform 1 0 37444 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 32660 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 22724 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 1840 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 24564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1372_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1373_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1374_
timestamp 1644511149
transform 1 0 45172 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1375_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1376_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1377_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1378_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1379_
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1380_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1381_
timestamp 1644511149
transform 1 0 44436 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 24288 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 21712 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 27232 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 47288 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 41492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1644511149
transform 1 0 46736 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform 1 0 47840 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1644511149
transform 1 0 12328 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 46460 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 47656 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1644511149
transform 1 0 31004 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 43700 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 11684 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46184 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 45540 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1644511149
transform 1 0 46736 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 40848 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 39192 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 41216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 14352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 15640 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 17204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 20424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27416 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2208 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45816 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 34868 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 41216 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 31188 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 27416 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45448 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35328 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46460 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 32752 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 34868 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 44988 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45264 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 39928 0 1 22848
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
