magic
tech sky130A
magscale 1 2
timestamp 1654519508
<< viali >>
rect 3065 47209 3099 47243
rect 48145 47141 48179 47175
rect 2053 47073 2087 47107
rect 9597 47073 9631 47107
rect 28733 47073 28767 47107
rect 43177 47073 43211 47107
rect 47041 47073 47075 47107
rect 1777 47005 1811 47039
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6377 47005 6411 47039
rect 7297 47005 7331 47039
rect 9413 47005 9447 47039
rect 11621 47005 11655 47039
rect 12357 47005 12391 47039
rect 13093 47005 13127 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 18245 47005 18279 47039
rect 20085 47005 20119 47039
rect 20361 47005 20395 47039
rect 24869 47005 24903 47039
rect 25513 47005 25547 47039
rect 28549 47005 28583 47039
rect 29745 47005 29779 47039
rect 31309 47005 31343 47039
rect 38301 47005 38335 47039
rect 40509 47005 40543 47039
rect 41889 47005 41923 47039
rect 42533 47005 42567 47039
rect 45201 47005 45235 47039
rect 47961 47005 47995 47039
rect 2789 46937 2823 46971
rect 4077 46937 4111 46971
rect 4997 46937 5031 46971
rect 6653 46937 6687 46971
rect 11805 46937 11839 46971
rect 12541 46937 12575 46971
rect 13461 46937 13495 46971
rect 14565 46937 14599 46971
rect 14749 46937 14783 46971
rect 18521 46937 18555 46971
rect 31125 46937 31159 46971
rect 40325 46937 40359 46971
rect 42717 46937 42751 46971
rect 45385 46937 45419 46971
rect 7481 46869 7515 46903
rect 29929 46869 29963 46903
rect 1869 46597 1903 46631
rect 47041 46597 47075 46631
rect 24593 46529 24627 46563
rect 38025 46529 38059 46563
rect 47961 46529 47995 46563
rect 3341 46461 3375 46495
rect 3525 46461 3559 46495
rect 4169 46461 4203 46495
rect 13093 46461 13127 46495
rect 13553 46461 13587 46495
rect 13737 46461 13771 46495
rect 14197 46461 14231 46495
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 32505 46461 32539 46495
rect 32689 46461 32723 46495
rect 33517 46461 33551 46495
rect 38209 46461 38243 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 2145 46325 2179 46359
rect 2881 46325 2915 46359
rect 10701 46325 10735 46359
rect 22017 46325 22051 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 3893 46121 3927 46155
rect 4629 46121 4663 46155
rect 19625 46121 19659 46155
rect 20177 46121 20211 46155
rect 24685 46121 24719 46155
rect 32689 46121 32723 46155
rect 33425 46121 33459 46155
rect 38209 46121 38243 46155
rect 10425 45985 10459 46019
rect 11069 45985 11103 46019
rect 20729 45985 20763 46019
rect 21281 45985 21315 46019
rect 25237 45985 25271 46019
rect 25789 45985 25823 46019
rect 41061 45985 41095 46019
rect 42533 45985 42567 46019
rect 48145 45985 48179 46019
rect 2789 45917 2823 45951
rect 3801 45917 3835 45951
rect 20085 45917 20119 45951
rect 24593 45917 24627 45951
rect 33333 45917 33367 45951
rect 38117 45917 38151 45951
rect 44005 45917 44039 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 10609 45849 10643 45883
rect 20913 45849 20947 45883
rect 25421 45849 25455 45883
rect 41245 45849 41279 45883
rect 44189 45849 44223 45883
rect 46489 45849 46523 45883
rect 2881 45781 2915 45815
rect 45753 45781 45787 45815
rect 10609 45577 10643 45611
rect 13737 45577 13771 45611
rect 20821 45577 20855 45611
rect 25421 45577 25455 45611
rect 41429 45577 41463 45611
rect 2145 45509 2179 45543
rect 42717 45509 42751 45543
rect 47961 45509 47995 45543
rect 10517 45441 10551 45475
rect 13645 45441 13679 45475
rect 20729 45441 20763 45475
rect 25329 45441 25363 45475
rect 41337 45441 41371 45475
rect 42625 45441 42659 45475
rect 43913 45441 43947 45475
rect 1961 45373 1995 45407
rect 2973 45373 3007 45407
rect 38669 45373 38703 45407
rect 38853 45373 38887 45407
rect 39865 45373 39899 45407
rect 43453 45373 43487 45407
rect 44649 45373 44683 45407
rect 44833 45373 44867 45407
rect 46029 45373 46063 45407
rect 44097 45237 44131 45271
rect 48053 45237 48087 45271
rect 38853 45033 38887 45067
rect 40417 45033 40451 45067
rect 45109 45033 45143 45067
rect 45753 45033 45787 45067
rect 44373 44965 44407 44999
rect 46305 44897 46339 44931
rect 48145 44897 48179 44931
rect 29561 44829 29595 44863
rect 38761 44829 38795 44863
rect 40325 44829 40359 44863
rect 44281 44829 44315 44863
rect 45017 44829 45051 44863
rect 45661 44829 45695 44863
rect 46489 44761 46523 44795
rect 29653 44693 29687 44727
rect 46305 44489 46339 44523
rect 47685 44489 47719 44523
rect 45109 44353 45143 44387
rect 45753 44353 45787 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 46949 44149 46983 44183
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 1409 43265 1443 43299
rect 47041 43265 47075 43299
rect 1685 43197 1719 43231
rect 47777 43197 47811 43231
rect 46305 42653 46339 42687
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47041 42177 47075 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 2237 41225 2271 41259
rect 46949 41225 46983 41259
rect 2145 41089 2179 41123
rect 46857 41089 46891 41123
rect 47961 41089 47995 41123
rect 48053 40885 48087 40919
rect 47685 40681 47719 40715
rect 1409 40477 1443 40511
rect 1593 40341 1627 40375
rect 47777 39797 47811 39831
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 46489 39321 46523 39355
rect 26157 39049 26191 39083
rect 46949 39049 46983 39083
rect 25973 38913 26007 38947
rect 26985 38913 27019 38947
rect 46857 38913 46891 38947
rect 47685 38913 47719 38947
rect 27353 38845 27387 38879
rect 47869 38845 47903 38879
rect 26157 38301 26191 38335
rect 47685 38301 47719 38335
rect 27445 38165 27479 38199
rect 25789 37825 25823 37859
rect 26985 37825 27019 37859
rect 47593 37825 47627 37859
rect 26065 37757 26099 37791
rect 27353 37757 27387 37791
rect 47685 37621 47719 37655
rect 48145 37281 48179 37315
rect 26157 37213 26191 37247
rect 46305 37213 46339 37247
rect 26893 37145 26927 37179
rect 46489 37145 46523 37179
rect 26249 36805 26283 36839
rect 26065 36737 26099 36771
rect 27353 36737 27387 36771
rect 27445 36669 27479 36703
rect 27537 36669 27571 36703
rect 26433 36533 26467 36567
rect 26985 36533 27019 36567
rect 28089 36533 28123 36567
rect 26985 36329 27019 36363
rect 2789 36193 2823 36227
rect 26709 36193 26743 36227
rect 1409 36125 1443 36159
rect 23673 36125 23707 36159
rect 25697 36125 25731 36159
rect 26617 36125 26651 36159
rect 1593 36057 1627 36091
rect 23489 35989 23523 36023
rect 25789 35989 25823 36023
rect 24225 35785 24259 35819
rect 2053 35649 2087 35683
rect 27169 35649 27203 35683
rect 22477 35581 22511 35615
rect 22753 35581 22787 35615
rect 24685 35581 24719 35615
rect 24961 35581 24995 35615
rect 27445 35581 27479 35615
rect 29653 35581 29687 35615
rect 29929 35581 29963 35615
rect 31401 35581 31435 35615
rect 26433 35445 26467 35479
rect 26985 35445 27019 35479
rect 27353 35445 27387 35479
rect 2237 35241 2271 35275
rect 22845 35241 22879 35275
rect 25881 35241 25915 35275
rect 29653 35241 29687 35275
rect 30205 35241 30239 35275
rect 30573 35241 30607 35275
rect 30849 35241 30883 35275
rect 27261 35105 27295 35139
rect 30297 35105 30331 35139
rect 1593 35037 1627 35071
rect 2145 35037 2179 35071
rect 22753 35037 22787 35071
rect 24501 35037 24535 35071
rect 26065 35037 26099 35071
rect 26157 35037 26191 35071
rect 26249 35037 26283 35071
rect 26341 35037 26375 35071
rect 29834 35037 29868 35071
rect 30757 35037 30791 35071
rect 31585 35037 31619 35071
rect 48145 35037 48179 35071
rect 27537 34969 27571 35003
rect 1409 34901 1443 34935
rect 24685 34901 24719 34935
rect 29009 34901 29043 34935
rect 29837 34901 29871 34935
rect 31677 34901 31711 34935
rect 47961 34901 47995 34935
rect 26985 34697 27019 34731
rect 28825 34697 28859 34731
rect 30113 34697 30147 34731
rect 27261 34629 27295 34663
rect 30665 34629 30699 34663
rect 20729 34561 20763 34595
rect 21833 34561 21867 34595
rect 24777 34561 24811 34595
rect 26985 34561 27019 34595
rect 28733 34561 28767 34595
rect 30021 34561 30055 34595
rect 30205 34561 30239 34595
rect 30849 34561 30883 34595
rect 48145 34561 48179 34595
rect 24869 34493 24903 34527
rect 27077 34425 27111 34459
rect 20913 34357 20947 34391
rect 22096 34357 22130 34391
rect 23581 34357 23615 34391
rect 31033 34357 31067 34391
rect 47961 34357 47995 34391
rect 22661 34153 22695 34187
rect 23213 34153 23247 34187
rect 26617 34153 26651 34187
rect 29745 34153 29779 34187
rect 48053 34153 48087 34187
rect 22293 34017 22327 34051
rect 24409 34017 24443 34051
rect 26801 34017 26835 34051
rect 28733 34017 28767 34051
rect 30297 34017 30331 34051
rect 31125 34017 31159 34051
rect 20821 33949 20855 33983
rect 21925 33949 21959 33983
rect 22097 33943 22131 33977
rect 22204 33949 22238 33983
rect 22477 33949 22511 33983
rect 23121 33949 23155 33983
rect 26617 33949 26651 33983
rect 26893 33949 26927 33983
rect 28457 33949 28491 33983
rect 28549 33949 28583 33983
rect 29929 33949 29963 33983
rect 30021 33949 30055 33983
rect 33333 33949 33367 33983
rect 33517 33949 33551 33983
rect 47869 33949 47903 33983
rect 24685 33881 24719 33915
rect 30389 33881 30423 33915
rect 31401 33881 31435 33915
rect 20913 33813 20947 33847
rect 26157 33813 26191 33847
rect 27077 33813 27111 33847
rect 28733 33813 28767 33847
rect 32873 33813 32907 33847
rect 33517 33813 33551 33847
rect 25053 33609 25087 33643
rect 27353 33609 27387 33643
rect 28549 33609 28583 33643
rect 29837 33609 29871 33643
rect 31585 33609 31619 33643
rect 35909 33609 35943 33643
rect 16037 33541 16071 33575
rect 25789 33541 25823 33575
rect 29377 33541 29411 33575
rect 1685 33473 1719 33507
rect 2697 33473 2731 33507
rect 19533 33473 19567 33507
rect 24869 33473 24903 33507
rect 25973 33473 26007 33507
rect 26985 33473 27019 33507
rect 27169 33473 27203 33507
rect 27813 33473 27847 33507
rect 27997 33473 28031 33507
rect 28365 33473 28399 33507
rect 29009 33473 29043 33507
rect 29193 33473 29227 33507
rect 30021 33473 30055 33507
rect 30849 33473 30883 33507
rect 31033 33473 31067 33507
rect 31125 33473 31159 33507
rect 31401 33473 31435 33507
rect 32137 33473 32171 33507
rect 32413 33473 32447 33507
rect 33057 33473 33091 33507
rect 33241 33473 33275 33507
rect 47041 33473 47075 33507
rect 47593 33473 47627 33507
rect 1409 33405 1443 33439
rect 14197 33405 14231 33439
rect 14381 33405 14415 33439
rect 19809 33405 19843 33439
rect 24409 33405 24443 33439
rect 24777 33405 24811 33439
rect 28089 33405 28123 33439
rect 28181 33405 28215 33439
rect 31217 33405 31251 33439
rect 32321 33405 32355 33439
rect 34161 33405 34195 33439
rect 34437 33405 34471 33439
rect 48053 33405 48087 33439
rect 33425 33337 33459 33371
rect 2789 33269 2823 33303
rect 3157 33269 3191 33303
rect 21281 33269 21315 33303
rect 26157 33269 26191 33303
rect 26985 33269 27019 33303
rect 32137 33269 32171 33303
rect 32597 33269 32631 33303
rect 33057 33269 33091 33303
rect 46857 33269 46891 33303
rect 47869 33269 47903 33303
rect 22937 33065 22971 33099
rect 25145 33065 25179 33099
rect 26065 33065 26099 33099
rect 27997 33065 28031 33099
rect 30573 33065 30607 33099
rect 32781 33065 32815 33099
rect 32873 33065 32907 33099
rect 34161 33065 34195 33099
rect 35357 33065 35391 33099
rect 27353 32997 27387 33031
rect 1409 32929 1443 32963
rect 11713 32929 11747 32963
rect 14197 32929 14231 32963
rect 16037 32929 16071 32963
rect 25881 32929 25915 32963
rect 26893 32929 26927 32963
rect 32965 32929 32999 32963
rect 33701 32929 33735 32963
rect 47133 32929 47167 32963
rect 47409 32929 47443 32963
rect 3985 32861 4019 32895
rect 11621 32861 11655 32895
rect 13369 32861 13403 32895
rect 21373 32861 21407 32895
rect 21741 32861 21775 32895
rect 22201 32861 22235 32895
rect 22385 32861 22419 32895
rect 22477 32861 22511 32895
rect 22615 32861 22649 32895
rect 22753 32861 22787 32895
rect 24961 32861 24995 32895
rect 25237 32861 25271 32895
rect 26065 32861 26099 32895
rect 26985 32861 27019 32895
rect 28733 32861 28767 32895
rect 29561 32861 29595 32895
rect 30757 32861 30791 32895
rect 30849 32861 30883 32895
rect 31033 32861 31067 32895
rect 31125 32861 31159 32895
rect 32689 32861 32723 32895
rect 33425 32861 33459 32895
rect 33609 32861 33643 32895
rect 33793 32861 33827 32895
rect 33977 32861 34011 32895
rect 35265 32861 35299 32895
rect 46581 32861 46615 32895
rect 1593 32793 1627 32827
rect 3249 32793 3283 32827
rect 13461 32793 13495 32827
rect 14381 32793 14415 32827
rect 21557 32793 21591 32827
rect 25789 32793 25823 32827
rect 27813 32793 27847 32827
rect 28013 32793 28047 32827
rect 47225 32793 47259 32827
rect 3801 32725 3835 32759
rect 11989 32725 12023 32759
rect 24777 32725 24811 32759
rect 26249 32725 26283 32759
rect 28181 32725 28215 32759
rect 28917 32725 28951 32759
rect 29745 32725 29779 32759
rect 14289 32521 14323 32555
rect 22385 32521 22419 32555
rect 23397 32521 23431 32555
rect 30205 32521 30239 32555
rect 33609 32521 33643 32555
rect 37657 32521 37691 32555
rect 2697 32453 2731 32487
rect 11805 32453 11839 32487
rect 25329 32453 25363 32487
rect 28641 32453 28675 32487
rect 29477 32453 29511 32487
rect 29285 32419 29319 32453
rect 14197 32385 14231 32419
rect 22017 32385 22051 32419
rect 22845 32385 22879 32419
rect 25605 32385 25639 32419
rect 30119 32385 30153 32419
rect 30297 32385 30331 32419
rect 31217 32385 31251 32419
rect 32321 32385 32355 32419
rect 33241 32385 33275 32419
rect 33425 32385 33459 32419
rect 36645 32385 36679 32419
rect 46489 32385 46523 32419
rect 47593 32385 47627 32419
rect 2513 32317 2547 32351
rect 3249 32317 3283 32351
rect 11529 32317 11563 32351
rect 22109 32317 22143 32351
rect 23121 32317 23155 32351
rect 25513 32317 25547 32351
rect 28825 32317 28859 32351
rect 29653 32317 29687 32351
rect 32413 32317 32447 32351
rect 37749 32317 37783 32351
rect 37841 32317 37875 32351
rect 46213 32317 46247 32351
rect 25789 32249 25823 32283
rect 31401 32249 31435 32283
rect 37289 32249 37323 32283
rect 2053 32181 2087 32215
rect 13277 32181 13311 32215
rect 23213 32181 23247 32215
rect 25605 32181 25639 32215
rect 32689 32181 32723 32215
rect 36461 32181 36495 32215
rect 47685 32181 47719 32215
rect 1409 31977 1443 32011
rect 12081 31977 12115 32011
rect 12725 31977 12759 32011
rect 27997 31909 28031 31943
rect 28733 31909 28767 31943
rect 33057 31909 33091 31943
rect 9413 31841 9447 31875
rect 9597 31841 9631 31875
rect 9873 31841 9907 31875
rect 15117 31841 15151 31875
rect 31861 31841 31895 31875
rect 35909 31841 35943 31875
rect 36185 31841 36219 31875
rect 37657 31841 37691 31875
rect 46305 31841 46339 31875
rect 46489 31841 46523 31875
rect 48145 31841 48179 31875
rect 1593 31773 1627 31807
rect 2789 31773 2823 31807
rect 11989 31773 12023 31807
rect 12173 31773 12207 31807
rect 12633 31773 12667 31807
rect 15025 31773 15059 31807
rect 20269 31773 20303 31807
rect 20361 31773 20395 31807
rect 20913 31773 20947 31807
rect 22017 31773 22051 31807
rect 22293 31773 22327 31807
rect 24869 31773 24903 31807
rect 25145 31773 25179 31807
rect 25697 31773 25731 31807
rect 25881 31773 25915 31807
rect 26111 31773 26145 31807
rect 27813 31773 27847 31807
rect 28549 31773 28583 31807
rect 31769 31773 31803 31807
rect 31953 31773 31987 31807
rect 32413 31773 32447 31807
rect 32561 31773 32595 31807
rect 32878 31773 32912 31807
rect 34713 31773 34747 31807
rect 34805 31773 34839 31807
rect 25053 31705 25087 31739
rect 25973 31705 26007 31739
rect 32689 31705 32723 31739
rect 32781 31705 32815 31739
rect 2881 31637 2915 31671
rect 15393 31637 15427 31671
rect 21005 31637 21039 31671
rect 21833 31637 21867 31671
rect 22201 31637 22235 31671
rect 24685 31637 24719 31671
rect 26249 31637 26283 31671
rect 9781 31433 9815 31467
rect 11621 31433 11655 31467
rect 15393 31433 15427 31467
rect 34897 31433 34931 31467
rect 37381 31433 37415 31467
rect 2145 31365 2179 31399
rect 15945 31365 15979 31399
rect 23489 31365 23523 31399
rect 24501 31365 24535 31399
rect 27905 31365 27939 31399
rect 30113 31365 30147 31399
rect 30329 31365 30363 31399
rect 46029 31365 46063 31399
rect 46121 31365 46155 31399
rect 47041 31365 47075 31399
rect 1961 31297 1995 31331
rect 9689 31297 9723 31331
rect 11529 31297 11563 31331
rect 15853 31297 15887 31331
rect 16773 31297 16807 31331
rect 23305 31297 23339 31331
rect 27721 31297 27755 31331
rect 36369 31297 36403 31331
rect 37289 31297 37323 31331
rect 2973 31229 3007 31263
rect 13645 31229 13679 31263
rect 13921 31229 13955 31263
rect 19165 31229 19199 31263
rect 19441 31229 19475 31263
rect 22017 31229 22051 31263
rect 22293 31229 22327 31263
rect 24225 31229 24259 31263
rect 33149 31229 33183 31263
rect 33425 31229 33459 31263
rect 36277 31229 36311 31263
rect 36737 31229 36771 31263
rect 16865 31093 16899 31127
rect 20913 31093 20947 31127
rect 23673 31093 23707 31127
rect 25973 31093 26007 31127
rect 30297 31093 30331 31127
rect 30481 31093 30515 31127
rect 15209 30889 15243 30923
rect 22109 30889 22143 30923
rect 22937 30889 22971 30923
rect 25789 30889 25823 30923
rect 26433 30889 26467 30923
rect 14105 30821 14139 30855
rect 12541 30753 12575 30787
rect 16037 30753 16071 30787
rect 19257 30753 19291 30787
rect 25605 30753 25639 30787
rect 10977 30685 11011 30719
rect 11713 30685 11747 30719
rect 11897 30685 11931 30719
rect 14381 30685 14415 30719
rect 15117 30685 15151 30719
rect 15301 30685 15335 30719
rect 15761 30685 15795 30719
rect 21833 30685 21867 30719
rect 21925 30685 21959 30719
rect 22753 30685 22787 30719
rect 23029 30685 23063 30719
rect 25513 30685 25547 30719
rect 26341 30685 26375 30719
rect 28273 30685 28307 30719
rect 33425 30685 33459 30719
rect 11069 30617 11103 30651
rect 12725 30617 12759 30651
rect 14473 30617 14507 30651
rect 19533 30617 19567 30651
rect 24685 30617 24719 30651
rect 31309 30617 31343 30651
rect 33609 30617 33643 30651
rect 11805 30549 11839 30583
rect 12817 30549 12851 30583
rect 12909 30549 12943 30583
rect 13093 30549 13127 30583
rect 14289 30549 14323 30583
rect 14657 30549 14691 30583
rect 17509 30549 17543 30583
rect 21005 30549 21039 30583
rect 21465 30549 21499 30583
rect 22569 30549 22603 30583
rect 24777 30549 24811 30583
rect 28365 30549 28399 30583
rect 31401 30549 31435 30583
rect 33793 30549 33827 30583
rect 13277 30345 13311 30379
rect 13829 30345 13863 30379
rect 15853 30345 15887 30379
rect 24501 30345 24535 30379
rect 11805 30277 11839 30311
rect 14841 30277 14875 30311
rect 22845 30277 22879 30311
rect 11529 30209 11563 30243
rect 14013 30209 14047 30243
rect 14749 30209 14783 30243
rect 15853 30209 15887 30243
rect 20913 30209 20947 30243
rect 22109 30209 22143 30243
rect 22293 30209 22327 30243
rect 22661 30209 22695 30243
rect 24498 30209 24532 30243
rect 27353 30209 27387 30243
rect 29837 30209 29871 30243
rect 33333 30209 33367 30243
rect 33517 30209 33551 30243
rect 33885 30209 33919 30243
rect 34529 30209 34563 30243
rect 14197 30141 14231 30175
rect 14289 30141 14323 30175
rect 21005 30141 21039 30175
rect 22385 30141 22419 30175
rect 22477 30141 22511 30175
rect 24961 30141 24995 30175
rect 27629 30141 27663 30175
rect 30113 30141 30147 30175
rect 33609 30141 33643 30175
rect 33701 30141 33735 30175
rect 34069 30141 34103 30175
rect 34805 30141 34839 30175
rect 24317 30073 24351 30107
rect 24869 30073 24903 30107
rect 21097 30005 21131 30039
rect 21281 30005 21315 30039
rect 29101 30005 29135 30039
rect 31585 30005 31619 30039
rect 36277 30005 36311 30039
rect 11805 29801 11839 29835
rect 12449 29801 12483 29835
rect 21465 29801 21499 29835
rect 22017 29801 22051 29835
rect 22661 29801 22695 29835
rect 27813 29801 27847 29835
rect 28825 29801 28859 29835
rect 29009 29801 29043 29835
rect 30849 29801 30883 29835
rect 31769 29801 31803 29835
rect 32505 29801 32539 29835
rect 33793 29801 33827 29835
rect 35173 29801 35207 29835
rect 36185 29801 36219 29835
rect 23121 29733 23155 29767
rect 11621 29665 11655 29699
rect 25697 29665 25731 29699
rect 26617 29665 26651 29699
rect 28641 29665 28675 29699
rect 29561 29665 29595 29699
rect 30941 29665 30975 29699
rect 31953 29665 31987 29699
rect 33517 29665 33551 29699
rect 36093 29665 36127 29699
rect 11437 29597 11471 29631
rect 11805 29597 11839 29631
rect 12357 29597 12391 29631
rect 15669 29597 15703 29631
rect 15761 29597 15795 29631
rect 16221 29597 16255 29631
rect 21646 29597 21680 29631
rect 22109 29597 22143 29631
rect 22569 29597 22603 29631
rect 22937 29597 22971 29631
rect 25513 29597 25547 29631
rect 25789 29597 25823 29631
rect 26249 29597 26283 29631
rect 27169 29597 27203 29631
rect 27262 29597 27296 29631
rect 27675 29597 27709 29631
rect 28825 29597 28859 29631
rect 30849 29597 30883 29631
rect 31677 29597 31711 29631
rect 32413 29597 32447 29631
rect 33595 29597 33629 29631
rect 35081 29597 35115 29631
rect 36185 29597 36219 29631
rect 47317 29597 47351 29631
rect 47593 29597 47627 29631
rect 16497 29529 16531 29563
rect 26433 29529 26467 29563
rect 27445 29529 27479 29563
rect 27537 29529 27571 29563
rect 28549 29529 28583 29563
rect 35909 29529 35943 29563
rect 11529 29461 11563 29495
rect 17969 29461 18003 29495
rect 21649 29461 21683 29495
rect 25329 29461 25363 29495
rect 29791 29461 29825 29495
rect 31217 29461 31251 29495
rect 31953 29461 31987 29495
rect 36369 29461 36403 29495
rect 17049 29257 17083 29291
rect 26157 29257 26191 29291
rect 27169 29257 27203 29291
rect 30665 29257 30699 29291
rect 13553 29189 13587 29223
rect 14657 29189 14691 29223
rect 19993 29189 20027 29223
rect 34805 29189 34839 29223
rect 9137 29121 9171 29155
rect 12725 29121 12759 29155
rect 14473 29121 14507 29155
rect 15577 29121 15611 29155
rect 16957 29121 16991 29155
rect 21833 29121 21867 29155
rect 22017 29121 22051 29155
rect 24409 29121 24443 29155
rect 24593 29121 24627 29155
rect 24685 29121 24719 29155
rect 24961 29121 24995 29155
rect 25605 29121 25639 29155
rect 25881 29121 25915 29155
rect 26985 29121 27019 29155
rect 27721 29121 27755 29155
rect 29929 29121 29963 29155
rect 30113 29121 30147 29155
rect 30205 29121 30239 29155
rect 30481 29121 30515 29155
rect 31125 29121 31159 29155
rect 31401 29121 31435 29155
rect 32229 29121 32263 29155
rect 32597 29121 32631 29155
rect 33241 29121 33275 29155
rect 33425 29121 33459 29155
rect 33517 29121 33551 29155
rect 33793 29121 33827 29155
rect 34437 29121 34471 29155
rect 34621 29121 34655 29155
rect 9321 29053 9355 29087
rect 10517 29053 10551 29087
rect 14289 29053 14323 29087
rect 15669 29053 15703 29087
rect 15945 29053 15979 29087
rect 18153 29053 18187 29087
rect 18337 29053 18371 29087
rect 24777 29053 24811 29087
rect 30297 29053 30331 29087
rect 31309 29053 31343 29087
rect 33609 29053 33643 29087
rect 32781 28985 32815 29019
rect 33977 28985 34011 29019
rect 12909 28917 12943 28951
rect 13645 28917 13679 28951
rect 22201 28917 22235 28951
rect 25145 28917 25179 28951
rect 25697 28917 25731 28951
rect 29009 28917 29043 28951
rect 31125 28917 31159 28951
rect 31585 28917 31619 28951
rect 32321 28917 32355 28951
rect 9781 28713 9815 28747
rect 26157 28713 26191 28747
rect 28457 28713 28491 28747
rect 29745 28713 29779 28747
rect 30849 28713 30883 28747
rect 33057 28713 33091 28747
rect 36553 28713 36587 28747
rect 29929 28645 29963 28679
rect 10885 28577 10919 28611
rect 11345 28577 11379 28611
rect 24685 28577 24719 28611
rect 27169 28577 27203 28611
rect 27629 28577 27663 28611
rect 33517 28577 33551 28611
rect 35081 28577 35115 28611
rect 9689 28509 9723 28543
rect 10977 28509 11011 28543
rect 14657 28509 14691 28543
rect 15393 28509 15427 28543
rect 16129 28509 16163 28543
rect 19349 28509 19383 28543
rect 21557 28509 21591 28543
rect 21925 28509 21959 28543
rect 22753 28509 22787 28543
rect 23029 28509 23063 28543
rect 24409 28509 24443 28543
rect 27261 28509 27295 28543
rect 29561 28509 29595 28543
rect 29653 28509 29687 28543
rect 30665 28509 30699 28543
rect 31861 28509 31895 28543
rect 32045 28509 32079 28543
rect 33241 28509 33275 28543
rect 33425 28509 33459 28543
rect 34805 28509 34839 28543
rect 47685 28509 47719 28543
rect 13369 28441 13403 28475
rect 14105 28441 14139 28475
rect 14381 28441 14415 28475
rect 15117 28441 15151 28475
rect 15485 28441 15519 28475
rect 19625 28441 19659 28475
rect 21741 28441 21775 28475
rect 21833 28441 21867 28475
rect 22937 28441 22971 28475
rect 28089 28441 28123 28475
rect 28273 28441 28307 28475
rect 30481 28441 30515 28475
rect 13461 28373 13495 28407
rect 14289 28373 14323 28407
rect 14473 28373 14507 28407
rect 15301 28373 15335 28407
rect 15669 28373 15703 28407
rect 16313 28373 16347 28407
rect 21097 28373 21131 28407
rect 22109 28373 22143 28407
rect 22569 28373 22603 28407
rect 32229 28373 32263 28407
rect 14473 28169 14507 28203
rect 14565 28169 14599 28203
rect 18429 28169 18463 28203
rect 20545 28169 20579 28203
rect 21189 28169 21223 28203
rect 25697 28169 25731 28203
rect 26341 28169 26375 28203
rect 28549 28169 28583 28203
rect 33885 28169 33919 28203
rect 34621 28169 34655 28203
rect 36001 28169 36035 28203
rect 11805 28101 11839 28135
rect 13553 28101 13587 28135
rect 16957 28101 16991 28135
rect 25605 28101 25639 28135
rect 30665 28101 30699 28135
rect 30849 28101 30883 28135
rect 31401 28101 31435 28135
rect 10885 28033 10919 28067
rect 14657 28033 14691 28067
rect 15301 28033 15335 28067
rect 15485 28033 15519 28067
rect 15577 28033 15611 28067
rect 16681 28033 16715 28067
rect 20453 28033 20487 28067
rect 21097 28033 21131 28067
rect 21281 28033 21315 28067
rect 22017 28033 22051 28067
rect 22201 28033 22235 28067
rect 22293 28033 22327 28067
rect 22753 28033 22787 28067
rect 24685 28033 24719 28067
rect 26249 28033 26283 28067
rect 26433 28033 26467 28067
rect 27445 28033 27479 28067
rect 28371 28033 28405 28067
rect 29101 28033 29135 28067
rect 29745 28033 29779 28067
rect 32321 28033 32355 28067
rect 32505 28033 32539 28067
rect 33793 28033 33827 28067
rect 34437 28033 34471 28067
rect 35265 28033 35299 28067
rect 35909 28033 35943 28067
rect 45753 28033 45787 28067
rect 47593 28033 47627 28067
rect 10977 27965 11011 27999
rect 11529 27965 11563 27999
rect 14197 27965 14231 27999
rect 15117 27965 15151 27999
rect 21833 27965 21867 27999
rect 27629 27965 27663 27999
rect 29837 27965 29871 27999
rect 32597 27965 32631 27999
rect 46581 27965 46615 27999
rect 29193 27897 29227 27931
rect 31585 27897 31619 27931
rect 35357 27897 35391 27931
rect 22937 27829 22971 27863
rect 24869 27829 24903 27863
rect 32137 27829 32171 27863
rect 47685 27829 47719 27863
rect 21649 27625 21683 27659
rect 22477 27625 22511 27659
rect 34970 27625 35004 27659
rect 12173 27557 12207 27591
rect 18061 27557 18095 27591
rect 21925 27557 21959 27591
rect 25973 27557 26007 27591
rect 27261 27557 27295 27591
rect 28365 27557 28399 27591
rect 30665 27557 30699 27591
rect 31217 27557 31251 27591
rect 32597 27557 32631 27591
rect 36461 27557 36495 27591
rect 9413 27489 9447 27523
rect 14565 27489 14599 27523
rect 21005 27489 21039 27523
rect 21557 27489 21591 27523
rect 22569 27489 22603 27523
rect 34713 27489 34747 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 12081 27421 12115 27455
rect 13369 27421 13403 27455
rect 14105 27421 14139 27455
rect 17969 27421 18003 27455
rect 20637 27421 20671 27455
rect 21471 27421 21505 27455
rect 21741 27421 21775 27455
rect 22477 27421 22511 27455
rect 24869 27421 24903 27455
rect 25881 27421 25915 27455
rect 27077 27421 27111 27455
rect 28549 27421 28583 27455
rect 28733 27421 28767 27455
rect 29653 27421 29687 27455
rect 30573 27421 30607 27455
rect 30757 27421 30791 27455
rect 31217 27421 31251 27455
rect 31401 27421 31435 27455
rect 31953 27421 31987 27455
rect 32046 27421 32080 27455
rect 32229 27421 32263 27455
rect 32459 27421 32493 27455
rect 45661 27421 45695 27455
rect 9597 27353 9631 27387
rect 11253 27353 11287 27387
rect 13461 27353 13495 27387
rect 14289 27353 14323 27387
rect 20821 27353 20855 27387
rect 28825 27353 28859 27387
rect 32321 27353 32355 27387
rect 22845 27285 22879 27319
rect 24961 27285 24995 27319
rect 29837 27285 29871 27319
rect 45753 27285 45787 27319
rect 9781 27081 9815 27115
rect 14657 27081 14691 27115
rect 15485 27081 15519 27115
rect 17417 27081 17451 27115
rect 23121 27081 23155 27115
rect 26341 27081 26375 27115
rect 46581 27081 46615 27115
rect 21281 27013 21315 27047
rect 27445 27013 27479 27047
rect 27629 27013 27663 27047
rect 28181 27013 28215 27047
rect 28397 27013 28431 27047
rect 30389 27013 30423 27047
rect 9689 26945 9723 26979
rect 10793 26945 10827 26979
rect 14473 26945 14507 26979
rect 15301 26945 15335 26979
rect 15577 26945 15611 26979
rect 17325 26945 17359 26979
rect 17969 26945 18003 26979
rect 20821 26945 20855 26979
rect 20913 26945 20947 26979
rect 21097 26945 21131 26979
rect 21833 26945 21867 26979
rect 22017 26945 22051 26979
rect 22201 26945 22235 26979
rect 22385 26945 22419 26979
rect 23029 26945 23063 26979
rect 24225 26945 24259 26979
rect 26157 26945 26191 26979
rect 29377 26945 29411 26979
rect 30297 26945 30331 26979
rect 31125 26945 31159 26979
rect 45293 26945 45327 26979
rect 10885 26877 10919 26911
rect 11529 26877 11563 26911
rect 11805 26877 11839 26911
rect 14289 26877 14323 26911
rect 18153 26877 18187 26911
rect 19809 26877 19843 26911
rect 21189 26877 21223 26911
rect 22109 26877 22143 26911
rect 24501 26877 24535 26911
rect 29193 26877 29227 26911
rect 29745 26877 29779 26911
rect 30941 26877 30975 26911
rect 24317 26809 24351 26843
rect 29653 26809 29687 26843
rect 13277 26741 13311 26775
rect 15301 26741 15335 26775
rect 22569 26741 22603 26775
rect 24409 26741 24443 26775
rect 28365 26741 28399 26775
rect 28549 26741 28583 26775
rect 31309 26741 31343 26775
rect 47777 26741 47811 26775
rect 11069 26537 11103 26571
rect 11897 26537 11931 26571
rect 17417 26537 17451 26571
rect 17969 26537 18003 26571
rect 19704 26537 19738 26571
rect 21189 26537 21223 26571
rect 22201 26537 22235 26571
rect 24777 26537 24811 26571
rect 26525 26537 26559 26571
rect 27445 26537 27479 26571
rect 45661 26537 45695 26571
rect 13093 26469 13127 26503
rect 14657 26469 14691 26503
rect 21741 26469 21775 26503
rect 23857 26469 23891 26503
rect 25053 26469 25087 26503
rect 27629 26469 27663 26503
rect 29745 26469 29779 26503
rect 31769 26469 31803 26503
rect 15209 26401 15243 26435
rect 19441 26401 19475 26435
rect 22293 26401 22327 26435
rect 32321 26401 32355 26435
rect 33793 26401 33827 26435
rect 11069 26333 11103 26367
rect 11253 26333 11287 26367
rect 11805 26333 11839 26367
rect 12909 26333 12943 26367
rect 15669 26333 15703 26367
rect 17877 26333 17911 26367
rect 22017 26333 22051 26367
rect 22109 26333 22143 26367
rect 22385 26333 22419 26367
rect 24685 26333 24719 26367
rect 24869 26333 24903 26367
rect 26433 26333 26467 26367
rect 27077 26333 27111 26367
rect 27445 26333 27479 26367
rect 28365 26333 28399 26367
rect 29561 26333 29595 26367
rect 31342 26333 31376 26367
rect 31861 26333 31895 26367
rect 32505 26333 32539 26367
rect 32597 26333 32631 26367
rect 32781 26333 32815 26367
rect 32873 26333 32907 26367
rect 33425 26333 33459 26367
rect 33613 26333 33647 26367
rect 33710 26333 33744 26367
rect 33977 26333 34011 26367
rect 43545 26333 43579 26367
rect 44281 26333 44315 26367
rect 45477 26333 45511 26367
rect 46305 26333 46339 26367
rect 14841 26265 14875 26299
rect 15025 26265 15059 26299
rect 15945 26265 15979 26299
rect 23489 26265 23523 26299
rect 23673 26265 23707 26299
rect 24409 26265 24443 26299
rect 28181 26265 28215 26299
rect 34161 26265 34195 26299
rect 46489 26265 46523 26299
rect 48145 26265 48179 26299
rect 14933 26197 14967 26231
rect 31217 26197 31251 26231
rect 31401 26197 31435 26231
rect 13461 25993 13495 26027
rect 15301 25993 15335 26027
rect 16037 25993 16071 26027
rect 18797 25993 18831 26027
rect 20729 25993 20763 26027
rect 26157 25993 26191 26027
rect 26985 25993 27019 26027
rect 27353 25993 27387 26027
rect 28825 25993 28859 26027
rect 11529 25925 11563 25959
rect 13093 25925 13127 25959
rect 13293 25925 13327 25959
rect 45385 25925 45419 25959
rect 10149 25857 10183 25891
rect 11713 25857 11747 25891
rect 11805 25857 11839 25891
rect 12265 25857 12299 25891
rect 14289 25857 14323 25891
rect 15117 25857 15151 25891
rect 15853 25857 15887 25891
rect 17049 25857 17083 25891
rect 18061 25857 18095 25891
rect 18705 25857 18739 25891
rect 20637 25857 20671 25891
rect 23029 25857 23063 25891
rect 23857 25857 23891 25891
rect 23949 25857 23983 25891
rect 24685 25857 24719 25891
rect 24869 25857 24903 25891
rect 25053 25857 25087 25891
rect 25145 25857 25179 25891
rect 25973 25857 26007 25891
rect 26249 25857 26283 25891
rect 28273 25857 28307 25891
rect 28641 25857 28675 25891
rect 29561 25857 29595 25891
rect 30849 25857 30883 25891
rect 30941 25857 30975 25891
rect 31217 25857 31251 25891
rect 32137 25857 32171 25891
rect 34345 25857 34379 25891
rect 47593 25857 47627 25891
rect 24041 25789 24075 25823
rect 27445 25789 27479 25823
rect 27629 25789 27663 25823
rect 29745 25789 29779 25823
rect 30665 25789 30699 25823
rect 32413 25789 32447 25823
rect 34621 25789 34655 25823
rect 45201 25789 45235 25823
rect 46857 25789 46891 25823
rect 11529 25721 11563 25755
rect 12449 25721 12483 25755
rect 14473 25721 14507 25755
rect 23489 25721 23523 25755
rect 24961 25721 24995 25755
rect 33885 25721 33919 25755
rect 10241 25653 10275 25687
rect 13277 25653 13311 25687
rect 17233 25653 17267 25687
rect 18153 25653 18187 25687
rect 22845 25653 22879 25687
rect 25789 25653 25823 25687
rect 28365 25653 28399 25687
rect 31125 25653 31159 25687
rect 36093 25653 36127 25687
rect 47685 25653 47719 25687
rect 14289 25449 14323 25483
rect 15117 25449 15151 25483
rect 15669 25449 15703 25483
rect 17601 25449 17635 25483
rect 23857 25449 23891 25483
rect 26617 25449 26651 25483
rect 28917 25449 28951 25483
rect 31401 25449 31435 25483
rect 32137 25449 32171 25483
rect 32873 25449 32907 25483
rect 34161 25449 34195 25483
rect 34897 25449 34931 25483
rect 44465 25449 44499 25483
rect 32321 25381 32355 25415
rect 9873 25313 9907 25347
rect 22385 25313 22419 25347
rect 31953 25313 31987 25347
rect 33701 25313 33735 25347
rect 46305 25313 46339 25347
rect 47961 25313 47995 25347
rect 12081 25245 12115 25279
rect 14933 25245 14967 25279
rect 15669 25245 15703 25279
rect 15853 25245 15887 25279
rect 17417 25245 17451 25279
rect 22109 25245 22143 25279
rect 24961 25245 24995 25279
rect 25145 25245 25179 25279
rect 25237 25245 25271 25279
rect 26433 25245 26467 25279
rect 28733 25245 28767 25279
rect 29837 25245 29871 25279
rect 29929 25245 29963 25279
rect 30113 25245 30147 25279
rect 30205 25245 30239 25279
rect 31217 25245 31251 25279
rect 32137 25245 32171 25279
rect 32781 25245 32815 25279
rect 33425 25245 33459 25279
rect 33609 25245 33643 25279
rect 33793 25245 33827 25279
rect 33977 25245 34011 25279
rect 34805 25245 34839 25279
rect 45477 25245 45511 25279
rect 46121 25245 46155 25279
rect 1869 25177 1903 25211
rect 10149 25177 10183 25211
rect 12173 25177 12207 25211
rect 14105 25177 14139 25211
rect 14321 25177 14355 25211
rect 31033 25177 31067 25211
rect 31861 25177 31895 25211
rect 1961 25109 1995 25143
rect 11621 25109 11655 25143
rect 14473 25109 14507 25143
rect 24777 25109 24811 25143
rect 29653 25109 29687 25143
rect 45569 25109 45603 25143
rect 28181 24905 28215 24939
rect 29469 24905 29503 24939
rect 31401 24905 31435 24939
rect 11529 24837 11563 24871
rect 11729 24837 11763 24871
rect 29377 24837 29411 24871
rect 31217 24837 31251 24871
rect 12449 24769 12483 24803
rect 18153 24769 18187 24803
rect 18337 24769 18371 24803
rect 18429 24769 18463 24803
rect 21281 24769 21315 24803
rect 22109 24769 22143 24803
rect 24961 24769 24995 24803
rect 25145 24769 25179 24803
rect 25237 24769 25271 24803
rect 28365 24769 28399 24803
rect 30481 24769 30515 24803
rect 31493 24769 31527 24803
rect 33885 24769 33919 24803
rect 40325 24769 40359 24803
rect 44649 24769 44683 24803
rect 45109 24769 45143 24803
rect 45753 24769 45787 24803
rect 46581 24769 46615 24803
rect 47593 24769 47627 24803
rect 47685 24769 47719 24803
rect 8585 24701 8619 24735
rect 8769 24701 8803 24735
rect 9045 24701 9079 24735
rect 13829 24701 13863 24735
rect 14013 24701 14047 24735
rect 14473 24701 14507 24735
rect 19441 24701 19475 24735
rect 19625 24701 19659 24735
rect 22753 24701 22787 24735
rect 23029 24701 23063 24735
rect 28641 24701 28675 24735
rect 30297 24701 30331 24735
rect 30757 24701 30791 24735
rect 34161 24701 34195 24735
rect 11897 24633 11931 24667
rect 22201 24633 22235 24667
rect 24501 24633 24535 24667
rect 24961 24633 24995 24667
rect 44465 24633 44499 24667
rect 11713 24565 11747 24599
rect 12541 24565 12575 24599
rect 18153 24565 18187 24599
rect 28549 24565 28583 24599
rect 30665 24565 30699 24599
rect 31217 24565 31251 24599
rect 35633 24565 35667 24599
rect 40417 24565 40451 24599
rect 45201 24565 45235 24599
rect 10517 24361 10551 24395
rect 12725 24361 12759 24395
rect 14197 24361 14231 24395
rect 23397 24361 23431 24395
rect 28549 24361 28583 24395
rect 30205 24361 30239 24395
rect 34805 24361 34839 24395
rect 11069 24293 11103 24327
rect 12909 24293 12943 24327
rect 11161 24225 11195 24259
rect 15117 24225 15151 24259
rect 15393 24225 15427 24259
rect 20269 24225 20303 24259
rect 22109 24225 22143 24259
rect 26709 24225 26743 24259
rect 28365 24225 28399 24259
rect 31125 24225 31159 24259
rect 40417 24225 40451 24259
rect 40693 24225 40727 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 10698 24157 10732 24191
rect 11805 24157 11839 24191
rect 12081 24157 12115 24191
rect 13369 24157 13403 24191
rect 14105 24157 14139 24191
rect 15025 24157 15059 24191
rect 16037 24157 16071 24191
rect 16957 24157 16991 24191
rect 19257 24157 19291 24191
rect 23305 24157 23339 24191
rect 25421 24157 25455 24191
rect 25789 24157 25823 24191
rect 26617 24157 26651 24191
rect 28273 24157 28307 24191
rect 28542 24157 28576 24191
rect 30113 24157 30147 24191
rect 30297 24157 30331 24191
rect 34713 24157 34747 24191
rect 40233 24157 40267 24191
rect 43361 24157 43395 24191
rect 43545 24157 43579 24191
rect 44005 24157 44039 24191
rect 45201 24157 45235 24191
rect 46305 24157 46339 24191
rect 12541 24089 12575 24123
rect 17233 24089 17267 24123
rect 19349 24089 19383 24123
rect 20453 24089 20487 24123
rect 25605 24089 25639 24123
rect 25697 24089 25731 24123
rect 30757 24089 30791 24123
rect 30941 24089 30975 24123
rect 44281 24089 44315 24123
rect 45753 24089 45787 24123
rect 10701 24021 10735 24055
rect 11621 24021 11655 24055
rect 11989 24021 12023 24055
rect 12741 24021 12775 24055
rect 13461 24021 13495 24055
rect 16037 24021 16071 24055
rect 18705 24021 18739 24055
rect 25973 24021 26007 24055
rect 26985 24021 27019 24055
rect 28733 24021 28767 24055
rect 43545 24021 43579 24055
rect 8953 23817 8987 23851
rect 17877 23817 17911 23851
rect 18639 23817 18673 23851
rect 19993 23817 20027 23851
rect 20637 23817 20671 23851
rect 26341 23817 26375 23851
rect 28457 23817 28491 23851
rect 30573 23817 30607 23851
rect 31217 23817 31251 23851
rect 34069 23817 34103 23851
rect 41521 23817 41555 23851
rect 43177 23817 43211 23851
rect 44189 23817 44223 23851
rect 11529 23749 11563 23783
rect 14105 23749 14139 23783
rect 18429 23749 18463 23783
rect 28089 23749 28123 23783
rect 29653 23749 29687 23783
rect 30389 23749 30423 23783
rect 42809 23749 42843 23783
rect 42993 23749 43027 23783
rect 45201 23749 45235 23783
rect 1409 23681 1443 23715
rect 8861 23681 8895 23715
rect 10977 23681 11011 23715
rect 13921 23681 13955 23715
rect 16681 23681 16715 23715
rect 17785 23681 17819 23715
rect 17969 23681 18003 23715
rect 19901 23681 19935 23715
rect 20545 23681 20579 23715
rect 21833 23681 21867 23715
rect 26157 23681 26191 23715
rect 26433 23681 26467 23715
rect 28273 23681 28307 23715
rect 29561 23681 29595 23715
rect 29745 23681 29779 23715
rect 30205 23681 30239 23715
rect 31033 23681 31067 23715
rect 31309 23681 31343 23715
rect 32689 23681 32723 23715
rect 33885 23681 33919 23715
rect 40141 23681 40175 23715
rect 41153 23681 41187 23715
rect 43821 23681 43855 23715
rect 44925 23681 44959 23715
rect 45937 23681 45971 23715
rect 47593 23681 47627 23715
rect 11989 23613 12023 23647
rect 14381 23613 14415 23647
rect 40233 23613 40267 23647
rect 41061 23613 41095 23647
rect 43729 23613 43763 23647
rect 46305 23613 46339 23647
rect 1593 23545 1627 23579
rect 11805 23545 11839 23579
rect 40509 23545 40543 23579
rect 10793 23477 10827 23511
rect 16773 23477 16807 23511
rect 18613 23477 18647 23511
rect 18797 23477 18831 23511
rect 21925 23477 21959 23511
rect 25973 23477 26007 23511
rect 31033 23477 31067 23511
rect 32781 23477 32815 23511
rect 47685 23477 47719 23511
rect 17785 23273 17819 23307
rect 26801 23273 26835 23307
rect 32965 23273 32999 23307
rect 43729 23273 43763 23307
rect 17141 23205 17175 23239
rect 28273 23205 28307 23239
rect 11713 23137 11747 23171
rect 15393 23137 15427 23171
rect 15669 23137 15703 23171
rect 20361 23137 20395 23171
rect 25053 23137 25087 23171
rect 27721 23137 27755 23171
rect 31217 23137 31251 23171
rect 40785 23137 40819 23171
rect 41429 23137 41463 23171
rect 43453 23137 43487 23171
rect 46305 23137 46339 23171
rect 46489 23137 46523 23171
rect 48145 23137 48179 23171
rect 10793 23069 10827 23103
rect 11437 23069 11471 23103
rect 14289 23069 14323 23103
rect 17693 23069 17727 23103
rect 19257 23069 19291 23103
rect 19441 23069 19475 23103
rect 20085 23069 20119 23103
rect 23397 23069 23431 23103
rect 27629 23069 27663 23103
rect 27813 23069 27847 23103
rect 28549 23069 28583 23103
rect 30205 23069 30239 23103
rect 30481 23069 30515 23103
rect 30573 23069 30607 23103
rect 33425 23069 33459 23103
rect 40325 23069 40359 23103
rect 43545 23069 43579 23103
rect 44189 23069 44223 23103
rect 44373 23069 44407 23103
rect 45385 23069 45419 23103
rect 25329 23001 25363 23035
rect 28273 23001 28307 23035
rect 30389 23001 30423 23035
rect 31493 23001 31527 23035
rect 40969 23001 41003 23035
rect 45661 23001 45695 23035
rect 10793 22933 10827 22967
rect 13185 22933 13219 22967
rect 14473 22933 14507 22967
rect 19625 22933 19659 22967
rect 21833 22933 21867 22967
rect 23489 22933 23523 22967
rect 28457 22933 28491 22967
rect 30757 22933 30791 22967
rect 33517 22933 33551 22967
rect 40141 22933 40175 22967
rect 43085 22933 43119 22967
rect 44281 22933 44315 22967
rect 11713 22729 11747 22763
rect 12541 22729 12575 22763
rect 18981 22729 19015 22763
rect 19257 22729 19291 22763
rect 27721 22729 27755 22763
rect 33885 22729 33919 22763
rect 39865 22729 39899 22763
rect 40693 22729 40727 22763
rect 47777 22729 47811 22763
rect 20821 22661 20855 22695
rect 22017 22661 22051 22695
rect 23673 22661 23707 22695
rect 28917 22661 28951 22695
rect 31033 22661 31067 22695
rect 31217 22661 31251 22695
rect 48145 22661 48179 22695
rect 9965 22593 9999 22627
rect 10793 22593 10827 22627
rect 11529 22593 11563 22627
rect 12449 22593 12483 22627
rect 13645 22593 13679 22627
rect 17417 22593 17451 22627
rect 18889 22593 18923 22627
rect 19073 22593 19107 22627
rect 20729 22593 20763 22627
rect 26985 22593 27019 22627
rect 27629 22593 27663 22627
rect 28733 22593 28767 22627
rect 29009 22593 29043 22627
rect 29101 22593 29135 22627
rect 30021 22593 30055 22627
rect 32137 22593 32171 22627
rect 40233 22593 40267 22627
rect 44925 22593 44959 22627
rect 45385 22593 45419 22627
rect 45569 22593 45603 22627
rect 47869 22593 47903 22627
rect 47961 22593 47995 22627
rect 10057 22525 10091 22559
rect 13829 22525 13863 22559
rect 15485 22525 15519 22559
rect 18705 22525 18739 22559
rect 21833 22525 21867 22559
rect 24133 22525 24167 22559
rect 24317 22525 24351 22559
rect 24593 22525 24627 22559
rect 29745 22525 29779 22559
rect 32413 22525 32447 22559
rect 46213 22525 46247 22559
rect 46489 22525 46523 22559
rect 47593 22525 47627 22559
rect 10333 22389 10367 22423
rect 10885 22389 10919 22423
rect 17509 22389 17543 22423
rect 27077 22389 27111 22423
rect 29285 22389 29319 22423
rect 31401 22389 31435 22423
rect 40325 22389 40359 22423
rect 44741 22389 44775 22423
rect 45753 22389 45787 22423
rect 10498 22185 10532 22219
rect 16852 22185 16886 22219
rect 25776 22185 25810 22219
rect 43085 22185 43119 22219
rect 12725 22117 12759 22151
rect 10241 22049 10275 22083
rect 11989 22049 12023 22083
rect 13461 22049 13495 22083
rect 16129 22049 16163 22083
rect 20913 22049 20947 22083
rect 23305 22049 23339 22083
rect 27261 22049 27295 22083
rect 29009 22049 29043 22083
rect 45753 22049 45787 22083
rect 46949 22049 46983 22083
rect 8953 21981 8987 22015
rect 9597 21981 9631 22015
rect 12541 21981 12575 22015
rect 13369 21981 13403 22015
rect 14289 21981 14323 22015
rect 16589 21981 16623 22015
rect 19533 21981 19567 22015
rect 20821 21981 20855 22015
rect 23213 21981 23247 22015
rect 25513 21981 25547 22015
rect 28181 21981 28215 22015
rect 28641 21981 28675 22015
rect 31953 21981 31987 22015
rect 34897 21981 34931 22015
rect 40141 21981 40175 22015
rect 40325 21981 40359 22015
rect 43361 21981 43395 22015
rect 45109 21981 45143 22015
rect 45293 21981 45327 22015
rect 14473 21913 14507 21947
rect 19257 21913 19291 21947
rect 19441 21913 19475 21947
rect 28825 21913 28859 21947
rect 40509 21913 40543 21947
rect 43085 21913 43119 21947
rect 45937 21913 45971 21947
rect 9045 21845 9079 21879
rect 9689 21845 9723 21879
rect 18337 21845 18371 21879
rect 19355 21845 19389 21879
rect 27997 21845 28031 21879
rect 31769 21845 31803 21879
rect 34713 21845 34747 21879
rect 43269 21845 43303 21879
rect 45293 21845 45327 21879
rect 14657 21641 14691 21675
rect 16865 21641 16899 21675
rect 29193 21641 29227 21675
rect 33885 21641 33919 21675
rect 48145 21641 48179 21675
rect 8861 21573 8895 21607
rect 20913 21573 20947 21607
rect 23213 21573 23247 21607
rect 27721 21573 27755 21607
rect 34437 21573 34471 21607
rect 34529 21573 34563 21607
rect 42533 21573 42567 21607
rect 43085 21573 43119 21607
rect 8677 21505 8711 21539
rect 14565 21505 14599 21539
rect 16681 21505 16715 21539
rect 17601 21505 17635 21539
rect 18521 21505 18555 21539
rect 18705 21505 18739 21539
rect 22201 21505 22235 21539
rect 27445 21505 27479 21539
rect 33425 21505 33459 21539
rect 42441 21505 42475 21539
rect 42625 21505 42659 21539
rect 44005 21505 44039 21539
rect 44189 21505 44223 21539
rect 44833 21505 44867 21539
rect 45293 21505 45327 21539
rect 46213 21505 46247 21539
rect 46489 21505 46523 21539
rect 47593 21505 47627 21539
rect 9137 21437 9171 21471
rect 17693 21437 17727 21471
rect 17969 21437 18003 21471
rect 22293 21437 22327 21471
rect 23029 21437 23063 21471
rect 23489 21437 23523 21471
rect 47869 21437 47903 21471
rect 34989 21369 35023 21403
rect 43361 21369 43395 21403
rect 44097 21369 44131 21403
rect 18521 21301 18555 21335
rect 21005 21301 21039 21335
rect 22569 21301 22603 21335
rect 33701 21301 33735 21335
rect 43545 21301 43579 21335
rect 44649 21301 44683 21335
rect 45477 21301 45511 21335
rect 45753 21301 45787 21335
rect 47685 21301 47719 21335
rect 16589 21097 16623 21131
rect 23857 21097 23891 21131
rect 26617 21097 26651 21131
rect 27629 21097 27663 21131
rect 14289 21029 14323 21063
rect 35817 21029 35851 21063
rect 8953 20961 8987 20995
rect 9137 20961 9171 20995
rect 22385 20961 22419 20995
rect 31677 20961 31711 20995
rect 43453 20961 43487 20995
rect 44097 20961 44131 20995
rect 45201 20961 45235 20995
rect 46305 20961 46339 20995
rect 48145 20961 48179 20995
rect 14105 20893 14139 20927
rect 14841 20893 14875 20927
rect 16589 20893 16623 20927
rect 17417 20893 17451 20927
rect 19257 20893 19291 20927
rect 21373 20893 21407 20927
rect 21649 20893 21683 20927
rect 22109 20893 22143 20927
rect 26433 20893 26467 20927
rect 27537 20893 27571 20927
rect 30573 20893 30607 20927
rect 43545 20893 43579 20927
rect 45845 20893 45879 20927
rect 10793 20825 10827 20859
rect 31769 20825 31803 20859
rect 32689 20825 32723 20859
rect 35265 20825 35299 20859
rect 35357 20825 35391 20859
rect 46489 20825 46523 20859
rect 14933 20757 14967 20791
rect 17509 20757 17543 20791
rect 19349 20757 19383 20791
rect 30665 20757 30699 20791
rect 45661 20757 45695 20791
rect 19717 20553 19751 20587
rect 22109 20553 22143 20587
rect 22385 20553 22419 20587
rect 22937 20553 22971 20587
rect 33517 20553 33551 20587
rect 44373 20553 44407 20587
rect 47685 20553 47719 20587
rect 18245 20485 18279 20519
rect 21833 20485 21867 20519
rect 32229 20485 32263 20519
rect 32321 20485 32355 20519
rect 45385 20485 45419 20519
rect 11713 20417 11747 20451
rect 11989 20417 12023 20451
rect 12173 20417 12207 20451
rect 12817 20417 12851 20451
rect 17233 20417 17267 20451
rect 17969 20417 18003 20451
rect 21005 20417 21039 20451
rect 22017 20417 22051 20451
rect 22201 20417 22235 20451
rect 22845 20417 22879 20451
rect 24685 20417 24719 20451
rect 26249 20417 26283 20451
rect 26985 20417 27019 20451
rect 31125 20417 31159 20451
rect 40049 20417 40083 20451
rect 42625 20417 42659 20451
rect 42809 20417 42843 20451
rect 43729 20417 43763 20451
rect 45201 20417 45235 20451
rect 47593 20417 47627 20451
rect 13093 20349 13127 20383
rect 13553 20349 13587 20383
rect 13829 20349 13863 20383
rect 28365 20349 28399 20383
rect 28549 20349 28583 20383
rect 28825 20349 28859 20383
rect 32597 20349 32631 20383
rect 40233 20349 40267 20383
rect 41889 20349 41923 20383
rect 43821 20349 43855 20383
rect 45845 20349 45879 20383
rect 11529 20213 11563 20247
rect 15301 20213 15335 20247
rect 17417 20213 17451 20247
rect 21097 20213 21131 20247
rect 24869 20213 24903 20247
rect 26341 20213 26375 20247
rect 27077 20213 27111 20247
rect 31309 20213 31343 20247
rect 31585 20213 31619 20247
rect 42625 20213 42659 20247
rect 40417 20009 40451 20043
rect 44005 20009 44039 20043
rect 12909 19941 12943 19975
rect 14105 19941 14139 19975
rect 14657 19941 14691 19975
rect 15669 19941 15703 19975
rect 20637 19941 20671 19975
rect 22845 19941 22879 19975
rect 43453 19941 43487 19975
rect 11437 19873 11471 19907
rect 15209 19873 15243 19907
rect 20361 19873 20395 19907
rect 21097 19873 21131 19907
rect 21373 19873 21407 19907
rect 25053 19873 25087 19907
rect 27077 19873 27111 19907
rect 28181 19873 28215 19907
rect 30665 19873 30699 19907
rect 32321 19873 32355 19907
rect 45753 19873 45787 19907
rect 45937 19873 45971 19907
rect 46213 19873 46247 19907
rect 2053 19805 2087 19839
rect 10609 19805 10643 19839
rect 10701 19805 10735 19839
rect 11161 19805 11195 19839
rect 13369 19805 13403 19839
rect 14289 19805 14323 19839
rect 15301 19805 15335 19839
rect 16957 19805 16991 19839
rect 18245 19805 18279 19839
rect 20269 19805 20303 19839
rect 24593 19805 24627 19839
rect 28365 19805 28399 19839
rect 30481 19805 30515 19839
rect 40325 19805 40359 19839
rect 42809 19805 42843 19839
rect 42993 19805 43027 19839
rect 43269 19805 43303 19839
rect 43453 19805 43487 19839
rect 44005 19805 44039 19839
rect 44189 19805 44223 19839
rect 45293 19805 45327 19839
rect 13461 19737 13495 19771
rect 25329 19737 25363 19771
rect 14381 19669 14415 19703
rect 14473 19669 14507 19703
rect 17049 19669 17083 19703
rect 18337 19669 18371 19703
rect 24409 19669 24443 19703
rect 28549 19669 28583 19703
rect 45109 19669 45143 19703
rect 15301 19465 15335 19499
rect 21005 19465 21039 19499
rect 22293 19465 22327 19499
rect 28365 19465 28399 19499
rect 28917 19465 28951 19499
rect 32137 19465 32171 19499
rect 43269 19465 43303 19499
rect 43821 19465 43855 19499
rect 14105 19397 14139 19431
rect 14933 19397 14967 19431
rect 15133 19397 15167 19431
rect 19901 19397 19935 19431
rect 20637 19397 20671 19431
rect 20837 19397 20871 19431
rect 27997 19397 28031 19431
rect 29745 19397 29779 19431
rect 47777 19397 47811 19431
rect 1777 19329 1811 19363
rect 13093 19329 13127 19363
rect 13185 19329 13219 19363
rect 14197 19329 14231 19363
rect 14289 19329 14323 19363
rect 17233 19329 17267 19363
rect 20085 19329 20119 19363
rect 20177 19329 20211 19363
rect 22201 19329 22235 19363
rect 24593 19329 24627 19363
rect 25421 19329 25455 19363
rect 28181 19329 28215 19363
rect 28825 19329 28859 19363
rect 29561 19329 29595 19363
rect 32321 19329 32355 19363
rect 42901 19329 42935 19363
rect 43085 19329 43119 19363
rect 43729 19329 43763 19363
rect 43913 19329 43947 19363
rect 45201 19329 45235 19363
rect 47869 19329 47903 19363
rect 47961 19329 47995 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 17509 19261 17543 19295
rect 18981 19261 19015 19295
rect 24685 19261 24719 19295
rect 30021 19261 30055 19295
rect 45385 19261 45419 19295
rect 45845 19261 45879 19295
rect 48145 19261 48179 19295
rect 13921 19193 13955 19227
rect 24961 19193 24995 19227
rect 47593 19193 47627 19227
rect 14473 19125 14507 19159
rect 15117 19125 15151 19159
rect 19901 19125 19935 19159
rect 20821 19125 20855 19159
rect 25421 19125 25455 19159
rect 2237 18921 2271 18955
rect 43913 18921 43947 18955
rect 18521 18853 18555 18887
rect 26985 18853 27019 18887
rect 28733 18853 28767 18887
rect 14105 18785 14139 18819
rect 18245 18785 18279 18819
rect 25237 18785 25271 18819
rect 25513 18785 25547 18819
rect 30481 18785 30515 18819
rect 45109 18785 45143 18819
rect 48145 18785 48179 18819
rect 2145 18717 2179 18751
rect 13369 18717 13403 18751
rect 13553 18717 13587 18751
rect 16681 18717 16715 18751
rect 18153 18717 18187 18751
rect 20545 18717 20579 18751
rect 20729 18717 20763 18751
rect 21189 18717 21223 18751
rect 23673 18717 23707 18751
rect 23857 18717 23891 18751
rect 24593 18717 24627 18751
rect 27997 18717 28031 18751
rect 28181 18717 28215 18751
rect 28917 18717 28951 18751
rect 29653 18717 29687 18751
rect 40509 18717 40543 18751
rect 40693 18717 40727 18751
rect 42441 18717 42475 18751
rect 42625 18717 42659 18751
rect 43453 18717 43487 18751
rect 44005 18717 44039 18751
rect 44189 18717 44223 18751
rect 44465 18717 44499 18751
rect 45017 18717 45051 18751
rect 45201 18717 45235 18751
rect 45845 18717 45879 18751
rect 46305 18717 46339 18751
rect 13461 18649 13495 18683
rect 14381 18649 14415 18683
rect 16957 18649 16991 18683
rect 20637 18649 20671 18683
rect 21465 18649 21499 18683
rect 24409 18649 24443 18683
rect 28273 18649 28307 18683
rect 29837 18649 29871 18683
rect 46489 18649 46523 18683
rect 15853 18581 15887 18615
rect 22937 18581 22971 18615
rect 23857 18581 23891 18615
rect 24777 18581 24811 18615
rect 40693 18581 40727 18615
rect 42625 18581 42659 18615
rect 1593 18377 1627 18411
rect 32137 18377 32171 18411
rect 47685 18377 47719 18411
rect 14289 18309 14323 18343
rect 15117 18309 15151 18343
rect 18061 18309 18095 18343
rect 18797 18309 18831 18343
rect 21281 18309 21315 18343
rect 22293 18309 22327 18343
rect 25145 18309 25179 18343
rect 45845 18309 45879 18343
rect 1409 18241 1443 18275
rect 14473 18241 14507 18275
rect 14565 18241 14599 18275
rect 15025 18241 15059 18275
rect 16773 18241 16807 18275
rect 17969 18241 18003 18275
rect 18613 18241 18647 18275
rect 21097 18241 21131 18275
rect 22201 18241 22235 18275
rect 24777 18241 24811 18275
rect 24961 18241 24995 18275
rect 27629 18241 27663 18275
rect 28273 18241 28307 18275
rect 30205 18241 30239 18275
rect 30849 18241 30883 18275
rect 32321 18241 32355 18275
rect 40417 18241 40451 18275
rect 40601 18241 40635 18275
rect 41337 18241 41371 18275
rect 42717 18241 42751 18275
rect 46857 18241 46891 18275
rect 47593 18241 47627 18275
rect 2513 18173 2547 18207
rect 2697 18173 2731 18207
rect 2973 18173 3007 18207
rect 20453 18173 20487 18207
rect 41613 18173 41647 18207
rect 42901 18173 42935 18207
rect 43453 18173 43487 18207
rect 44005 18173 44039 18207
rect 44189 18173 44223 18207
rect 29009 18105 29043 18139
rect 14289 18037 14323 18071
rect 16957 18037 16991 18071
rect 30297 18037 30331 18071
rect 31125 18037 31159 18071
rect 31309 18037 31343 18071
rect 40417 18037 40451 18071
rect 41429 18037 41463 18071
rect 41521 18037 41555 18071
rect 46949 18037 46983 18071
rect 2881 17833 2915 17867
rect 21465 17833 21499 17867
rect 24409 17833 24443 17867
rect 45385 17833 45419 17867
rect 41061 17765 41095 17799
rect 42257 17765 42291 17799
rect 44189 17765 44223 17799
rect 30757 17697 30791 17731
rect 40785 17697 40819 17731
rect 41705 17697 41739 17731
rect 46489 17697 46523 17731
rect 2145 17629 2179 17663
rect 2789 17629 2823 17663
rect 14749 17629 14783 17663
rect 14841 17629 14875 17663
rect 16405 17629 16439 17663
rect 24593 17629 24627 17663
rect 27629 17629 27663 17663
rect 27997 17629 28031 17663
rect 28273 17629 28307 17663
rect 28641 17629 28675 17663
rect 30573 17629 30607 17663
rect 41889 17629 41923 17663
rect 42165 17629 42199 17663
rect 43821 17629 43855 17663
rect 43913 17629 43947 17663
rect 44281 17629 44315 17663
rect 45017 17629 45051 17663
rect 46305 17629 46339 17663
rect 16589 17561 16623 17595
rect 18245 17561 18279 17595
rect 21189 17561 21223 17595
rect 28917 17561 28951 17595
rect 32413 17561 32447 17595
rect 42533 17561 42567 17595
rect 45201 17561 45235 17595
rect 48145 17561 48179 17595
rect 2237 17493 2271 17527
rect 15025 17493 15059 17527
rect 41245 17493 41279 17527
rect 16773 17289 16807 17323
rect 24133 17289 24167 17323
rect 25145 17289 25179 17323
rect 1961 17221 1995 17255
rect 23121 17221 23155 17255
rect 24225 17221 24259 17255
rect 45385 17221 45419 17255
rect 47685 17221 47719 17255
rect 14565 17153 14599 17187
rect 15117 17153 15151 17187
rect 16681 17153 16715 17187
rect 20177 17153 20211 17187
rect 22937 17153 22971 17187
rect 23029 17153 23063 17187
rect 24041 17153 24075 17187
rect 25053 17153 25087 17187
rect 25237 17153 25271 17187
rect 25881 17153 25915 17187
rect 27077 17153 27111 17187
rect 27629 17153 27663 17187
rect 42625 17153 42659 17187
rect 47593 17153 47627 17187
rect 1777 17085 1811 17119
rect 2789 17085 2823 17119
rect 42533 17085 42567 17119
rect 45201 17085 45235 17119
rect 46857 17085 46891 17119
rect 22753 17017 22787 17051
rect 23305 17017 23339 17051
rect 23857 17017 23891 17051
rect 24869 17017 24903 17051
rect 42993 17017 43027 17051
rect 14381 16949 14415 16983
rect 15209 16949 15243 16983
rect 20361 16949 20395 16983
rect 24409 16949 24443 16983
rect 25421 16949 25455 16983
rect 26065 16949 26099 16983
rect 2053 16745 2087 16779
rect 27261 16745 27295 16779
rect 47685 16745 47719 16779
rect 23765 16677 23799 16711
rect 24593 16677 24627 16711
rect 14105 16609 14139 16643
rect 17693 16609 17727 16643
rect 17969 16609 18003 16643
rect 23397 16609 23431 16643
rect 24869 16609 24903 16643
rect 25053 16609 25087 16643
rect 26893 16609 26927 16643
rect 45017 16609 45051 16643
rect 45477 16609 45511 16643
rect 17601 16541 17635 16575
rect 18429 16541 18463 16575
rect 19257 16541 19291 16575
rect 21649 16541 21683 16575
rect 24777 16541 24811 16575
rect 24961 16541 24995 16575
rect 27077 16541 27111 16575
rect 44281 16541 44315 16575
rect 14381 16473 14415 16507
rect 44373 16473 44407 16507
rect 45201 16473 45235 16507
rect 15853 16405 15887 16439
rect 18613 16405 18647 16439
rect 19349 16405 19383 16439
rect 21833 16405 21867 16439
rect 23857 16405 23891 16439
rect 23137 16201 23171 16235
rect 23305 16201 23339 16235
rect 23765 16201 23799 16235
rect 26157 16201 26191 16235
rect 18061 16133 18095 16167
rect 22937 16133 22971 16167
rect 24685 16133 24719 16167
rect 13737 16065 13771 16099
rect 14657 16065 14691 16099
rect 15485 16065 15519 16099
rect 15761 16065 15795 16099
rect 15945 16065 15979 16099
rect 20085 16065 20119 16099
rect 20913 16065 20947 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 23949 16065 23983 16099
rect 41245 16065 41279 16099
rect 47777 16065 47811 16099
rect 13829 15997 13863 16031
rect 14105 15997 14139 16031
rect 17785 15997 17819 16031
rect 22109 15997 22143 16031
rect 24409 15997 24443 16031
rect 14749 15861 14783 15895
rect 15301 15861 15335 15895
rect 19533 15861 19567 15895
rect 20085 15861 20119 15895
rect 20913 15861 20947 15895
rect 22385 15861 22419 15895
rect 23121 15861 23155 15895
rect 41337 15861 41371 15895
rect 17785 15657 17819 15691
rect 17969 15657 18003 15691
rect 23581 15657 23615 15691
rect 24409 15657 24443 15691
rect 25329 15657 25363 15691
rect 21373 15589 21407 15623
rect 15025 15521 15059 15555
rect 19625 15521 19659 15555
rect 19901 15521 19935 15555
rect 21833 15521 21867 15555
rect 22109 15521 22143 15555
rect 41245 15521 41279 15555
rect 41429 15521 41463 15555
rect 42901 15521 42935 15555
rect 2053 15453 2087 15487
rect 14749 15453 14783 15487
rect 18429 15453 18463 15487
rect 24409 15453 24443 15487
rect 25237 15453 25271 15487
rect 17601 15385 17635 15419
rect 17817 15385 17851 15419
rect 16497 15317 16531 15351
rect 18613 15317 18647 15351
rect 14933 15113 14967 15147
rect 17433 15113 17467 15147
rect 17601 15113 17635 15147
rect 19809 15113 19843 15147
rect 21189 15113 21223 15147
rect 23029 15113 23063 15147
rect 17233 15045 17267 15079
rect 21833 15045 21867 15079
rect 1777 14977 1811 15011
rect 14749 14977 14783 15011
rect 18061 14977 18095 15011
rect 21097 14977 21131 15011
rect 22017 14977 22051 15011
rect 22109 14977 22143 15011
rect 22937 14977 22971 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 18337 14909 18371 14943
rect 21833 14841 21867 14875
rect 17417 14773 17451 14807
rect 2237 14569 2271 14603
rect 18061 14569 18095 14603
rect 19441 14569 19475 14603
rect 17049 14433 17083 14467
rect 17693 14433 17727 14467
rect 2145 14365 2179 14399
rect 16957 14365 16991 14399
rect 17141 14365 17175 14399
rect 17785 14365 17819 14399
rect 19349 14365 19383 14399
rect 22201 14365 22235 14399
rect 22845 14365 22879 14399
rect 22293 14229 22327 14263
rect 22937 14229 22971 14263
rect 22017 13957 22051 13991
rect 16681 13889 16715 13923
rect 46857 13889 46891 13923
rect 16865 13821 16899 13855
rect 18521 13821 18555 13855
rect 21833 13821 21867 13855
rect 22293 13821 22327 13855
rect 46949 13685 46983 13719
rect 16957 13345 16991 13379
rect 19441 13345 19475 13379
rect 21097 13345 21131 13379
rect 22477 13345 22511 13379
rect 46489 13345 46523 13379
rect 15761 13277 15795 13311
rect 16405 13277 16439 13311
rect 19257 13277 19291 13311
rect 22017 13277 22051 13311
rect 46305 13277 46339 13311
rect 15853 13209 15887 13243
rect 16589 13209 16623 13243
rect 22201 13209 22235 13243
rect 48145 13209 48179 13243
rect 1593 12937 1627 12971
rect 16037 12869 16071 12903
rect 16865 12869 16899 12903
rect 22017 12869 22051 12903
rect 1409 12801 1443 12835
rect 15945 12801 15979 12835
rect 16681 12801 16715 12835
rect 21833 12801 21867 12835
rect 47777 12801 47811 12835
rect 18061 12733 18095 12767
rect 22293 12733 22327 12767
rect 16773 12393 16807 12427
rect 17785 12393 17819 12427
rect 22661 12393 22695 12427
rect 16681 12189 16715 12223
rect 17693 12189 17727 12223
rect 22569 12189 22603 12223
rect 47777 11509 47811 11543
rect 46305 11169 46339 11203
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 46949 10761 46983 10795
rect 46857 10625 46891 10659
rect 47593 10625 47627 10659
rect 46397 10421 46431 10455
rect 47685 10421 47719 10455
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 47869 9537 47903 9571
rect 48053 9401 48087 9435
rect 47777 8857 47811 8891
rect 47869 8789 47903 8823
rect 45109 8449 45143 8483
rect 44925 8245 44959 8279
rect 43637 8041 43671 8075
rect 44097 8041 44131 8075
rect 44465 8041 44499 8075
rect 45569 7905 45603 7939
rect 47593 7905 47627 7939
rect 44005 7837 44039 7871
rect 47317 7837 47351 7871
rect 45201 7769 45235 7803
rect 45293 7769 45327 7803
rect 47961 7497 47995 7531
rect 44833 7429 44867 7463
rect 48145 7361 48179 7395
rect 44741 7293 44775 7327
rect 45569 7293 45603 7327
rect 48053 6409 48087 6443
rect 47961 6273 47995 6307
rect 40233 5661 40267 5695
rect 42809 5661 42843 5695
rect 40325 5525 40359 5559
rect 42625 5525 42659 5559
rect 41061 5321 41095 5355
rect 37473 5253 37507 5287
rect 38393 5253 38427 5287
rect 42625 5253 42659 5287
rect 43545 5253 43579 5287
rect 18705 5185 18739 5219
rect 39681 5185 39715 5219
rect 40509 5185 40543 5219
rect 40969 5185 41003 5219
rect 43821 5185 43855 5219
rect 47869 5185 47903 5219
rect 37381 5117 37415 5151
rect 38669 5117 38703 5151
rect 42533 5117 42567 5151
rect 48053 5049 48087 5083
rect 18797 4981 18831 5015
rect 39773 4981 39807 5015
rect 40325 4981 40359 5015
rect 25605 4641 25639 4675
rect 27261 4641 27295 4675
rect 40325 4641 40359 4675
rect 40509 4641 40543 4675
rect 42165 4641 42199 4675
rect 42901 4641 42935 4675
rect 43913 4641 43947 4675
rect 47593 4641 47627 4675
rect 9505 4573 9539 4607
rect 18061 4573 18095 4607
rect 19349 4573 19383 4607
rect 19441 4573 19475 4607
rect 19993 4573 20027 4607
rect 20637 4573 20671 4607
rect 21373 4573 21407 4607
rect 22017 4573 22051 4607
rect 22661 4573 22695 4607
rect 25421 4573 25455 4607
rect 46673 4573 46707 4607
rect 47317 4573 47351 4607
rect 21465 4505 21499 4539
rect 42993 4505 43027 4539
rect 18153 4437 18187 4471
rect 20085 4437 20119 4471
rect 20729 4437 20763 4471
rect 22109 4437 22143 4471
rect 22753 4437 22787 4471
rect 46765 4437 46799 4471
rect 19809 4233 19843 4267
rect 20453 4233 20487 4267
rect 40969 4233 41003 4267
rect 37473 4165 37507 4199
rect 37565 4165 37599 4199
rect 38485 4165 38519 4199
rect 40601 4165 40635 4199
rect 47777 4165 47811 4199
rect 10149 4097 10183 4131
rect 13737 4097 13771 4131
rect 17233 4097 17267 4131
rect 17877 4097 17911 4131
rect 19073 4097 19107 4131
rect 19717 4097 19751 4131
rect 20361 4097 20395 4131
rect 21005 4097 21039 4131
rect 21833 4097 21867 4131
rect 22477 4097 22511 4131
rect 22569 4097 22603 4131
rect 23121 4097 23155 4131
rect 23765 4097 23799 4131
rect 36737 4097 36771 4131
rect 40785 4097 40819 4131
rect 42993 4097 43027 4131
rect 46765 4097 46799 4131
rect 2053 4029 2087 4063
rect 2237 4029 2271 4063
rect 3065 4029 3099 4063
rect 7389 4029 7423 4063
rect 7573 4029 7607 4063
rect 7849 4029 7883 4063
rect 17325 4029 17359 4063
rect 39497 4029 39531 4063
rect 39681 4029 39715 4063
rect 23213 3961 23247 3995
rect 36553 3961 36587 3995
rect 47961 3961 47995 3995
rect 10241 3893 10275 3927
rect 11713 3893 11747 3927
rect 13829 3893 13863 3927
rect 17969 3893 18003 3927
rect 19165 3893 19199 3927
rect 21097 3893 21131 3927
rect 21925 3893 21959 3927
rect 23857 3893 23891 3927
rect 40141 3893 40175 3927
rect 43085 3893 43119 3927
rect 43821 3893 43855 3927
rect 46305 3893 46339 3927
rect 46949 3893 46983 3927
rect 2973 3689 3007 3723
rect 3985 3689 4019 3723
rect 17049 3689 17083 3723
rect 18613 3689 18647 3723
rect 21557 3689 21591 3723
rect 22201 3689 22235 3723
rect 23765 3689 23799 3723
rect 40233 3689 40267 3723
rect 43177 3689 43211 3723
rect 43545 3689 43579 3723
rect 6469 3553 6503 3587
rect 9321 3553 9355 3587
rect 9781 3553 9815 3587
rect 42165 3553 42199 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 1685 3485 1719 3519
rect 2145 3485 2179 3519
rect 2881 3485 2915 3519
rect 5273 3485 5307 3519
rect 5917 3485 5951 3519
rect 8217 3485 8251 3519
rect 12081 3485 12115 3519
rect 14289 3485 14323 3519
rect 16957 3485 16991 3519
rect 17601 3485 17635 3519
rect 18521 3485 18555 3519
rect 19533 3485 19567 3519
rect 20361 3485 20395 3519
rect 20821 3485 20855 3519
rect 20913 3485 20947 3519
rect 21465 3485 21499 3519
rect 22109 3485 22143 3519
rect 23213 3485 23247 3519
rect 23673 3485 23707 3519
rect 25421 3485 25455 3519
rect 27261 3485 27295 3519
rect 32965 3485 32999 3519
rect 33793 3485 33827 3519
rect 38117 3485 38151 3519
rect 38669 3485 38703 3519
rect 40141 3485 40175 3519
rect 40785 3485 40819 3519
rect 43085 3485 43119 3519
rect 44005 3485 44039 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 5365 3417 5399 3451
rect 6101 3417 6135 3451
rect 9505 3417 9539 3451
rect 25605 3417 25639 3451
rect 33057 3417 33091 3451
rect 40969 3417 41003 3451
rect 48145 3417 48179 3451
rect 2237 3349 2271 3383
rect 8309 3349 8343 3383
rect 12173 3349 12207 3383
rect 17693 3349 17727 3383
rect 19625 3349 19659 3383
rect 38761 3349 38795 3383
rect 44097 3349 44131 3383
rect 45753 3349 45787 3383
rect 36737 3145 36771 3179
rect 40877 3145 40911 3179
rect 41337 3145 41371 3179
rect 48053 3145 48087 3179
rect 1961 3077 1995 3111
rect 8217 3077 8251 3111
rect 11713 3077 11747 3111
rect 14013 3077 14047 3111
rect 17785 3077 17819 3111
rect 18889 3077 18923 3111
rect 33057 3077 33091 3111
rect 38025 3077 38059 3111
rect 42993 3077 43027 3111
rect 45385 3077 45419 3111
rect 1777 3009 1811 3043
rect 6561 3009 6595 3043
rect 7573 3009 7607 3043
rect 11529 3009 11563 3043
rect 13829 3009 13863 3043
rect 16865 3009 16899 3043
rect 17693 3009 17727 3043
rect 18797 3009 18831 3043
rect 22293 3009 22327 3043
rect 22937 3009 22971 3043
rect 25605 3009 25639 3043
rect 27169 3009 27203 3043
rect 36277 3009 36311 3043
rect 37841 3009 37875 3043
rect 41521 3009 41555 3043
rect 42809 3009 42843 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2237 2941 2271 2975
rect 8033 2941 8067 2975
rect 8493 2941 8527 2975
rect 11989 2941 12023 2975
rect 14289 2941 14323 2975
rect 16773 2941 16807 2975
rect 17233 2941 17267 2975
rect 19441 2941 19475 2975
rect 19625 2941 19659 2975
rect 19993 2941 20027 2975
rect 23121 2941 23155 2975
rect 23397 2941 23431 2975
rect 32873 2941 32907 2975
rect 33517 2941 33551 2975
rect 39313 2941 39347 2975
rect 40233 2941 40267 2975
rect 40417 2941 40451 2975
rect 43269 2941 43303 2975
rect 47041 2941 47075 2975
rect 22477 2873 22511 2907
rect 25881 2805 25915 2839
rect 26065 2805 26099 2839
rect 26985 2805 27019 2839
rect 36369 2805 36403 2839
rect 3065 2601 3099 2635
rect 8217 2601 8251 2635
rect 16865 2601 16899 2635
rect 17601 2601 17635 2635
rect 18245 2601 18279 2635
rect 19349 2601 19383 2635
rect 20177 2601 20211 2635
rect 20913 2601 20947 2635
rect 23765 2601 23799 2635
rect 24961 2601 24995 2635
rect 25513 2601 25547 2635
rect 28641 2601 28675 2635
rect 35541 2601 35575 2635
rect 38301 2601 38335 2635
rect 40417 2601 40451 2635
rect 2145 2533 2179 2567
rect 27629 2533 27663 2567
rect 29745 2533 29779 2567
rect 39313 2533 39347 2567
rect 42441 2533 42475 2567
rect 5273 2465 5307 2499
rect 23029 2465 23063 2499
rect 36461 2465 36495 2499
rect 41337 2465 41371 2499
rect 46489 2465 46523 2499
rect 47869 2465 47903 2499
rect 4997 2397 5031 2431
rect 8953 2397 8987 2431
rect 16681 2397 16715 2431
rect 17509 2397 17543 2431
rect 18153 2397 18187 2431
rect 19257 2397 19291 2431
rect 20085 2397 20119 2431
rect 22385 2397 22419 2431
rect 22753 2397 22787 2431
rect 23673 2397 23707 2431
rect 25697 2397 25731 2431
rect 29929 2397 29963 2431
rect 35725 2397 35759 2431
rect 37657 2397 37691 2431
rect 40049 2397 40083 2431
rect 40417 2397 40451 2431
rect 41153 2397 41187 2431
rect 42625 2397 42659 2431
rect 43637 2397 43671 2431
rect 43913 2397 43947 2431
rect 46213 2397 46247 2431
rect 47685 2397 47719 2431
rect 1869 2329 1903 2363
rect 2789 2329 2823 2363
rect 15669 2329 15703 2363
rect 20821 2329 20855 2363
rect 24869 2329 24903 2363
rect 26249 2329 26283 2363
rect 27445 2329 27479 2363
rect 28549 2329 28583 2363
rect 36277 2329 36311 2363
rect 38209 2329 38243 2363
rect 39129 2329 39163 2363
rect 45385 2329 45419 2363
rect 9137 2261 9171 2295
rect 15761 2261 15795 2295
rect 26341 2261 26375 2295
rect 37473 2261 37507 2295
rect 40601 2261 40635 2295
rect 45477 2261 45511 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 3053 47243 3111 47249
rect 3053 47209 3065 47243
rect 3099 47240 3111 47243
rect 34238 47240 34244 47252
rect 3099 47212 34244 47240
rect 3099 47209 3111 47212
rect 3053 47203 3111 47209
rect 34238 47200 34244 47212
rect 34296 47200 34302 47252
rect 39758 47172 39764 47184
rect 6886 47144 39764 47172
rect 2041 47107 2099 47113
rect 2041 47073 2053 47107
rect 2087 47104 2099 47107
rect 6886 47104 6914 47144
rect 39758 47132 39764 47144
rect 39816 47132 39822 47184
rect 48133 47175 48191 47181
rect 48133 47172 48145 47175
rect 39960 47144 48145 47172
rect 2087 47076 6914 47104
rect 9585 47107 9643 47113
rect 2087 47073 2099 47076
rect 2041 47067 2099 47073
rect 9585 47073 9597 47107
rect 9631 47104 9643 47107
rect 28721 47107 28779 47113
rect 9631 47076 26234 47104
rect 9631 47073 9643 47076
rect 9585 47067 9643 47073
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47036 1823 47039
rect 1946 47036 1952 47048
rect 1811 47008 1952 47036
rect 1811 47005 1823 47008
rect 1765 46999 1823 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4706 47036 4712 47048
rect 4667 47008 4712 47036
rect 3789 46999 3847 47005
rect 4706 46996 4712 47008
rect 4764 46996 4770 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 5868 47008 6377 47036
rect 5868 46996 5874 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 7282 47036 7288 47048
rect 7243 47008 7288 47036
rect 6365 46999 6423 47005
rect 7282 46996 7288 47008
rect 7340 46996 7346 47048
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 11606 47036 11612 47048
rect 11567 47008 11612 47036
rect 9401 46999 9459 47005
rect 11606 46996 11612 47008
rect 11664 46996 11670 47048
rect 12250 46996 12256 47048
rect 12308 47036 12314 47048
rect 12345 47039 12403 47045
rect 12345 47036 12357 47039
rect 12308 47008 12357 47036
rect 12308 46996 12314 47008
rect 12345 47005 12357 47008
rect 12391 47005 12403 47039
rect 12345 46999 12403 47005
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12952 47008 13093 47036
rect 12952 46996 12958 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 13081 46999 13139 47005
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16942 47036 16948 47048
rect 16903 47008 16948 47036
rect 16669 46999 16727 47005
rect 16942 46996 16948 47008
rect 17000 46996 17006 47048
rect 18233 47039 18291 47045
rect 18233 47005 18245 47039
rect 18279 47036 18291 47039
rect 18690 47036 18696 47048
rect 18279 47008 18696 47036
rect 18279 47005 18291 47008
rect 18233 46999 18291 47005
rect 18690 46996 18696 47008
rect 18748 46996 18754 47048
rect 19978 46996 19984 47048
rect 20036 47036 20042 47048
rect 20073 47039 20131 47045
rect 20073 47036 20085 47039
rect 20036 47008 20085 47036
rect 20036 46996 20042 47008
rect 20073 47005 20085 47008
rect 20119 47005 20131 47039
rect 20346 47036 20352 47048
rect 20307 47008 20352 47036
rect 20073 46999 20131 47005
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 24854 47036 24860 47048
rect 24815 47008 24860 47036
rect 24854 46996 24860 47008
rect 24912 46996 24918 47048
rect 25498 47036 25504 47048
rect 25459 47008 25504 47036
rect 25498 46996 25504 47008
rect 25556 46996 25562 47048
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 2777 46931 2835 46937
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 2792 46900 2820 46931
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 4982 46968 4988 46980
rect 4943 46940 4988 46968
rect 4982 46928 4988 46940
rect 5040 46928 5046 46980
rect 6638 46968 6644 46980
rect 6599 46940 6644 46968
rect 6638 46928 6644 46940
rect 6696 46928 6702 46980
rect 8202 46968 8208 46980
rect 7484 46940 8208 46968
rect 7484 46909 7512 46940
rect 8202 46928 8208 46940
rect 8260 46928 8266 46980
rect 11698 46928 11704 46980
rect 11756 46968 11762 46980
rect 11793 46971 11851 46977
rect 11793 46968 11805 46971
rect 11756 46940 11805 46968
rect 11756 46928 11762 46940
rect 11793 46937 11805 46940
rect 11839 46937 11851 46971
rect 11793 46931 11851 46937
rect 12434 46928 12440 46980
rect 12492 46968 12498 46980
rect 12529 46971 12587 46977
rect 12529 46968 12541 46971
rect 12492 46940 12541 46968
rect 12492 46928 12498 46940
rect 12529 46937 12541 46940
rect 12575 46937 12587 46971
rect 12529 46931 12587 46937
rect 13354 46928 13360 46980
rect 13412 46968 13418 46980
rect 13449 46971 13507 46977
rect 13449 46968 13461 46971
rect 13412 46940 13461 46968
rect 13412 46928 13418 46940
rect 13449 46937 13461 46940
rect 13495 46937 13507 46971
rect 13449 46931 13507 46937
rect 14553 46971 14611 46977
rect 14553 46937 14565 46971
rect 14599 46937 14611 46971
rect 14553 46931 14611 46937
rect 2648 46872 2820 46900
rect 7469 46903 7527 46909
rect 2648 46860 2654 46872
rect 7469 46869 7481 46903
rect 7515 46869 7527 46903
rect 7469 46863 7527 46869
rect 13538 46860 13544 46912
rect 13596 46900 13602 46912
rect 14568 46900 14596 46931
rect 14642 46928 14648 46980
rect 14700 46968 14706 46980
rect 14737 46971 14795 46977
rect 14737 46968 14749 46971
rect 14700 46940 14749 46968
rect 14700 46928 14706 46940
rect 14737 46937 14749 46940
rect 14783 46937 14795 46971
rect 14737 46931 14795 46937
rect 18509 46971 18567 46977
rect 18509 46937 18521 46971
rect 18555 46968 18567 46971
rect 18874 46968 18880 46980
rect 18555 46940 18880 46968
rect 18555 46937 18567 46940
rect 18509 46931 18567 46937
rect 18874 46928 18880 46940
rect 18932 46928 18938 46980
rect 26206 46968 26234 47076
rect 28721 47073 28733 47107
rect 28767 47104 28779 47107
rect 32398 47104 32404 47116
rect 28767 47076 32404 47104
rect 28767 47073 28779 47076
rect 28721 47067 28779 47073
rect 32398 47064 32404 47076
rect 32456 47064 32462 47116
rect 37642 47064 37648 47116
rect 37700 47104 37706 47116
rect 39960 47104 39988 47144
rect 48133 47141 48145 47144
rect 48179 47141 48191 47175
rect 48133 47135 48191 47141
rect 43162 47104 43168 47116
rect 37700 47076 39988 47104
rect 43123 47076 43168 47104
rect 37700 47064 37706 47076
rect 43162 47064 43168 47076
rect 43220 47064 43226 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28537 47039 28595 47045
rect 28537 47036 28549 47039
rect 28408 47008 28549 47036
rect 28408 46996 28414 47008
rect 28537 47005 28549 47008
rect 28583 47005 28595 47039
rect 28537 46999 28595 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 30926 46996 30932 47048
rect 30984 47036 30990 47048
rect 31297 47039 31355 47045
rect 31297 47036 31309 47039
rect 30984 47008 31309 47036
rect 30984 46996 30990 47008
rect 31297 47005 31309 47008
rect 31343 47005 31355 47039
rect 31297 46999 31355 47005
rect 38010 46996 38016 47048
rect 38068 47036 38074 47048
rect 38289 47039 38347 47045
rect 38289 47036 38301 47039
rect 38068 47008 38301 47036
rect 38068 46996 38074 47008
rect 38289 47005 38301 47008
rect 38335 47005 38347 47039
rect 38289 46999 38347 47005
rect 40126 46996 40132 47048
rect 40184 47036 40190 47048
rect 40497 47039 40555 47045
rect 40497 47036 40509 47039
rect 40184 47008 40509 47036
rect 40184 46996 40190 47008
rect 40497 47005 40509 47008
rect 40543 47005 40555 47039
rect 40497 46999 40555 47005
rect 41877 47039 41935 47045
rect 41877 47005 41889 47039
rect 41923 47036 41935 47039
rect 42521 47039 42579 47045
rect 42521 47036 42533 47039
rect 41923 47008 42533 47036
rect 41923 47005 41935 47008
rect 41877 46999 41935 47005
rect 42521 47005 42533 47008
rect 42567 47005 42579 47039
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 42521 46999 42579 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47949 47039 48007 47045
rect 47949 47036 47961 47039
rect 47728 47008 47961 47036
rect 47728 46996 47734 47008
rect 47949 47005 47961 47008
rect 47995 47005 48007 47039
rect 47949 46999 48007 47005
rect 30190 46968 30196 46980
rect 26206 46940 30196 46968
rect 30190 46928 30196 46940
rect 30248 46928 30254 46980
rect 31018 46928 31024 46980
rect 31076 46968 31082 46980
rect 31113 46971 31171 46977
rect 31113 46968 31125 46971
rect 31076 46940 31125 46968
rect 31076 46928 31082 46940
rect 31113 46937 31125 46940
rect 31159 46937 31171 46971
rect 31113 46931 31171 46937
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 42702 46968 42708 46980
rect 42663 46940 42708 46968
rect 40313 46931 40371 46937
rect 29914 46900 29920 46912
rect 13596 46872 14596 46900
rect 29875 46872 29920 46900
rect 13596 46860 13602 46872
rect 29914 46860 29920 46872
rect 29972 46860 29978 46912
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 42702 46928 42708 46940
rect 42760 46928 42766 46980
rect 45373 46971 45431 46977
rect 45373 46937 45385 46971
rect 45419 46968 45431 46971
rect 45462 46968 45468 46980
rect 45419 46940 45468 46968
rect 45419 46937 45431 46940
rect 45373 46931 45431 46937
rect 45462 46928 45468 46940
rect 45520 46928 45526 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1854 46628 1860 46640
rect 1815 46600 1860 46628
rect 1854 46588 1860 46600
rect 1912 46588 1918 46640
rect 24854 46628 24860 46640
rect 24596 46600 24860 46628
rect 24596 46569 24624 46600
rect 24854 46588 24860 46600
rect 24912 46588 24918 46640
rect 27062 46588 27068 46640
rect 27120 46628 27126 46640
rect 34054 46628 34060 46640
rect 27120 46600 34060 46628
rect 27120 46588 27126 46600
rect 34054 46588 34060 46600
rect 34112 46588 34118 46640
rect 47026 46628 47032 46640
rect 46987 46600 47032 46628
rect 47026 46588 47032 46600
rect 47084 46588 47090 46640
rect 24581 46563 24639 46569
rect 24581 46529 24593 46563
rect 24627 46529 24639 46563
rect 38010 46560 38016 46572
rect 37971 46532 38016 46560
rect 24581 46523 24639 46529
rect 38010 46520 38016 46532
rect 38068 46520 38074 46572
rect 47946 46560 47952 46572
rect 47907 46532 47952 46560
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 3329 46495 3387 46501
rect 3329 46461 3341 46495
rect 3375 46461 3387 46495
rect 3329 46455 3387 46461
rect 3513 46495 3571 46501
rect 3513 46461 3525 46495
rect 3559 46492 3571 46495
rect 3878 46492 3884 46504
rect 3559 46464 3884 46492
rect 3559 46461 3571 46464
rect 3513 46455 3571 46461
rect 3344 46424 3372 46455
rect 3878 46452 3884 46464
rect 3936 46452 3942 46504
rect 3970 46452 3976 46504
rect 4028 46492 4034 46504
rect 4157 46495 4215 46501
rect 4157 46492 4169 46495
rect 4028 46464 4169 46492
rect 4028 46452 4034 46464
rect 4157 46461 4169 46464
rect 4203 46461 4215 46495
rect 4157 46455 4215 46461
rect 13081 46495 13139 46501
rect 13081 46461 13093 46495
rect 13127 46492 13139 46495
rect 13541 46495 13599 46501
rect 13541 46492 13553 46495
rect 13127 46464 13553 46492
rect 13127 46461 13139 46464
rect 13081 46455 13139 46461
rect 13541 46461 13553 46464
rect 13587 46461 13599 46495
rect 13722 46492 13728 46504
rect 13683 46464 13728 46492
rect 13541 46455 13599 46461
rect 13722 46452 13728 46464
rect 13780 46452 13786 46504
rect 14182 46492 14188 46504
rect 14143 46464 14188 46492
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 19426 46492 19432 46504
rect 19387 46464 19432 46492
rect 19426 46452 19432 46464
rect 19484 46452 19490 46504
rect 19613 46495 19671 46501
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 20162 46492 20168 46504
rect 19659 46464 20168 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 20162 46452 20168 46464
rect 20220 46452 20226 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 32490 46492 32496 46504
rect 32451 46464 32496 46492
rect 32490 46452 32496 46464
rect 32548 46452 32554 46504
rect 32677 46495 32735 46501
rect 32677 46461 32689 46495
rect 32723 46492 32735 46495
rect 33410 46492 33416 46504
rect 32723 46464 33416 46492
rect 32723 46461 32735 46464
rect 32677 46455 32735 46461
rect 33410 46452 33416 46464
rect 33468 46452 33474 46504
rect 33505 46495 33563 46501
rect 33505 46461 33517 46495
rect 33551 46461 33563 46495
rect 38194 46492 38200 46504
rect 38155 46464 38200 46492
rect 33505 46455 33563 46461
rect 4614 46424 4620 46436
rect 3344 46396 4620 46424
rect 4614 46384 4620 46396
rect 4672 46384 4678 46436
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 33520 46424 33548 46455
rect 38194 46452 38200 46464
rect 38252 46452 38258 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 42889 46455 42947 46461
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45370 46492 45376 46504
rect 45331 46464 45376 46492
rect 45189 46455 45247 46461
rect 32272 46396 33548 46424
rect 32272 46384 32278 46396
rect 42242 46384 42248 46436
rect 42300 46424 42306 46436
rect 42904 46424 42932 46455
rect 42300 46396 42932 46424
rect 45204 46424 45232 46455
rect 45370 46452 45376 46464
rect 45428 46452 45434 46504
rect 45646 46424 45652 46436
rect 45204 46396 45652 46424
rect 42300 46384 42306 46396
rect 45646 46384 45652 46396
rect 45704 46384 45710 46436
rect 2133 46359 2191 46365
rect 2133 46325 2145 46359
rect 2179 46356 2191 46359
rect 2314 46356 2320 46368
rect 2179 46328 2320 46356
rect 2179 46325 2191 46328
rect 2133 46319 2191 46325
rect 2314 46316 2320 46328
rect 2372 46316 2378 46368
rect 2774 46316 2780 46368
rect 2832 46356 2838 46368
rect 2869 46359 2927 46365
rect 2869 46356 2881 46359
rect 2832 46328 2881 46356
rect 2832 46316 2838 46328
rect 2869 46325 2881 46328
rect 2915 46325 2927 46359
rect 2869 46319 2927 46325
rect 10410 46316 10416 46368
rect 10468 46356 10474 46368
rect 10689 46359 10747 46365
rect 10689 46356 10701 46359
rect 10468 46328 10701 46356
rect 10468 46316 10474 46328
rect 10689 46325 10701 46328
rect 10735 46325 10747 46359
rect 10689 46319 10747 46325
rect 20714 46316 20720 46368
rect 20772 46356 20778 46368
rect 22005 46359 22063 46365
rect 22005 46356 22017 46359
rect 20772 46328 22017 46356
rect 20772 46316 20778 46328
rect 22005 46325 22017 46328
rect 22051 46325 22063 46359
rect 22005 46319 22063 46325
rect 41046 46316 41052 46368
rect 41104 46356 41110 46368
rect 41233 46359 41291 46365
rect 41233 46356 41245 46359
rect 41104 46328 41245 46356
rect 41104 46316 41110 46328
rect 41233 46325 41245 46328
rect 41279 46325 41291 46359
rect 41233 46319 41291 46325
rect 47210 46316 47216 46368
rect 47268 46356 47274 46368
rect 48041 46359 48099 46365
rect 48041 46356 48053 46359
rect 47268 46328 48053 46356
rect 47268 46316 47274 46328
rect 48041 46325 48053 46328
rect 48087 46325 48099 46359
rect 48041 46319 48099 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3878 46152 3884 46164
rect 3839 46124 3884 46152
rect 3878 46112 3884 46124
rect 3936 46112 3942 46164
rect 4614 46152 4620 46164
rect 4575 46124 4620 46152
rect 4614 46112 4620 46124
rect 4672 46112 4678 46164
rect 19426 46112 19432 46164
rect 19484 46152 19490 46164
rect 19613 46155 19671 46161
rect 19613 46152 19625 46155
rect 19484 46124 19625 46152
rect 19484 46112 19490 46124
rect 19613 46121 19625 46124
rect 19659 46121 19671 46155
rect 20162 46152 20168 46164
rect 20123 46124 20168 46152
rect 19613 46115 19671 46121
rect 20162 46112 20168 46124
rect 20220 46112 20226 46164
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 32490 46112 32496 46164
rect 32548 46152 32554 46164
rect 32677 46155 32735 46161
rect 32677 46152 32689 46155
rect 32548 46124 32689 46152
rect 32548 46112 32554 46124
rect 32677 46121 32689 46124
rect 32723 46121 32735 46155
rect 33410 46152 33416 46164
rect 33371 46124 33416 46152
rect 32677 46115 32735 46121
rect 33410 46112 33416 46124
rect 33468 46112 33474 46164
rect 38194 46152 38200 46164
rect 38155 46124 38200 46152
rect 38194 46112 38200 46124
rect 38252 46112 38258 46164
rect 45830 46084 45836 46096
rect 38120 46056 45836 46084
rect 10410 46016 10416 46028
rect 10371 45988 10416 46016
rect 10410 45976 10416 45988
rect 10468 45976 10474 46028
rect 10962 45976 10968 46028
rect 11020 46016 11026 46028
rect 11057 46019 11115 46025
rect 11057 46016 11069 46019
rect 11020 45988 11069 46016
rect 11020 45976 11026 45988
rect 11057 45985 11069 45988
rect 11103 45985 11115 46019
rect 20714 46016 20720 46028
rect 20675 45988 20720 46016
rect 11057 45979 11115 45985
rect 20714 45976 20720 45988
rect 20772 45976 20778 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25225 46019 25283 46025
rect 25225 45985 25237 46019
rect 25271 46016 25283 46019
rect 25498 46016 25504 46028
rect 25271 45988 25504 46016
rect 25271 45985 25283 45988
rect 25225 45979 25283 45985
rect 25498 45976 25504 45988
rect 25556 45976 25562 46028
rect 25774 46016 25780 46028
rect 25735 45988 25780 46016
rect 25774 45976 25780 45988
rect 25832 45976 25838 46028
rect 38120 45960 38148 46056
rect 45830 46044 45836 46056
rect 45888 46044 45894 46096
rect 41046 46016 41052 46028
rect 41007 45988 41052 46016
rect 41046 45976 41052 45988
rect 41104 45976 41110 46028
rect 42518 46016 42524 46028
rect 42479 45988 42524 46016
rect 42518 45976 42524 45988
rect 42576 45976 42582 46028
rect 48130 46016 48136 46028
rect 48091 45988 48136 46016
rect 48130 45976 48136 45988
rect 48188 45976 48194 46028
rect 2777 45951 2835 45957
rect 2777 45917 2789 45951
rect 2823 45917 2835 45951
rect 2777 45911 2835 45917
rect 2792 45880 2820 45911
rect 3050 45908 3056 45960
rect 3108 45948 3114 45960
rect 3789 45951 3847 45957
rect 3789 45948 3801 45951
rect 3108 45920 3801 45948
rect 3108 45908 3114 45920
rect 3789 45917 3801 45920
rect 3835 45917 3847 45951
rect 20070 45948 20076 45960
rect 20031 45920 20076 45948
rect 3789 45911 3847 45917
rect 20070 45908 20076 45920
rect 20128 45908 20134 45960
rect 24581 45951 24639 45957
rect 24581 45917 24593 45951
rect 24627 45948 24639 45951
rect 24854 45948 24860 45960
rect 24627 45920 24860 45948
rect 24627 45917 24639 45920
rect 24581 45911 24639 45917
rect 24854 45908 24860 45920
rect 24912 45908 24918 45960
rect 33321 45951 33379 45957
rect 33321 45917 33333 45951
rect 33367 45948 33379 45951
rect 38102 45948 38108 45960
rect 33367 45920 35894 45948
rect 38015 45920 38108 45948
rect 33367 45917 33379 45920
rect 33321 45911 33379 45917
rect 10594 45880 10600 45892
rect 2792 45852 6914 45880
rect 10555 45852 10600 45880
rect 2866 45812 2872 45824
rect 2827 45784 2872 45812
rect 2866 45772 2872 45784
rect 2924 45772 2930 45824
rect 6886 45812 6914 45852
rect 10594 45840 10600 45852
rect 10652 45840 10658 45892
rect 20898 45880 20904 45892
rect 20859 45852 20904 45880
rect 20898 45840 20904 45852
rect 20956 45840 20962 45892
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 35866 45880 35894 45920
rect 38102 45908 38108 45920
rect 38160 45908 38166 45960
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43993 45951 44051 45957
rect 43993 45948 44005 45951
rect 43864 45920 44005 45948
rect 43864 45908 43870 45920
rect 43993 45917 44005 45920
rect 44039 45917 44051 45951
rect 43993 45911 44051 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 46290 45948 46296 45960
rect 46251 45920 46296 45948
rect 46290 45908 46296 45920
rect 46348 45908 46354 45960
rect 40034 45880 40040 45892
rect 35866 45852 40040 45880
rect 40034 45840 40040 45852
rect 40092 45840 40098 45892
rect 41230 45880 41236 45892
rect 41191 45852 41236 45880
rect 41230 45840 41236 45852
rect 41288 45840 41294 45892
rect 44177 45883 44235 45889
rect 44177 45849 44189 45883
rect 44223 45880 44235 45883
rect 44450 45880 44456 45892
rect 44223 45852 44456 45880
rect 44223 45849 44235 45852
rect 44177 45843 44235 45849
rect 44450 45840 44456 45852
rect 44508 45840 44514 45892
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 10502 45812 10508 45824
rect 6886 45784 10508 45812
rect 10502 45772 10508 45784
rect 10560 45772 10566 45824
rect 45554 45772 45560 45824
rect 45612 45812 45618 45824
rect 45741 45815 45799 45821
rect 45741 45812 45753 45815
rect 45612 45784 45753 45812
rect 45612 45772 45618 45784
rect 45741 45781 45753 45784
rect 45787 45781 45799 45815
rect 45741 45775 45799 45781
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 10594 45608 10600 45620
rect 10555 45580 10600 45608
rect 10594 45568 10600 45580
rect 10652 45568 10658 45620
rect 13722 45608 13728 45620
rect 13683 45580 13728 45608
rect 13722 45568 13728 45580
rect 13780 45568 13786 45620
rect 16114 45568 16120 45620
rect 16172 45608 16178 45620
rect 17402 45608 17408 45620
rect 16172 45580 17408 45608
rect 16172 45568 16178 45580
rect 17402 45568 17408 45580
rect 17460 45568 17466 45620
rect 20809 45611 20867 45617
rect 20809 45577 20821 45611
rect 20855 45608 20867 45611
rect 20898 45608 20904 45620
rect 20855 45580 20904 45608
rect 20855 45577 20867 45580
rect 20809 45571 20867 45577
rect 20898 45568 20904 45580
rect 20956 45568 20962 45620
rect 25406 45608 25412 45620
rect 25367 45580 25412 45608
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 41417 45611 41475 45617
rect 41417 45577 41429 45611
rect 41463 45608 41475 45611
rect 42610 45608 42616 45620
rect 41463 45580 42616 45608
rect 41463 45577 41475 45580
rect 41417 45571 41475 45577
rect 42610 45568 42616 45580
rect 42668 45568 42674 45620
rect 45094 45568 45100 45620
rect 45152 45608 45158 45620
rect 45152 45580 45600 45608
rect 45152 45568 45158 45580
rect 2133 45543 2191 45549
rect 2133 45509 2145 45543
rect 2179 45540 2191 45543
rect 2866 45540 2872 45552
rect 2179 45512 2872 45540
rect 2179 45509 2191 45512
rect 2133 45503 2191 45509
rect 2866 45500 2872 45512
rect 2924 45500 2930 45552
rect 24854 45540 24860 45552
rect 12544 45512 24860 45540
rect 10502 45472 10508 45484
rect 10415 45444 10508 45472
rect 10502 45432 10508 45444
rect 10560 45472 10566 45484
rect 12544 45472 12572 45512
rect 24854 45500 24860 45512
rect 24912 45500 24918 45552
rect 42702 45540 42708 45552
rect 42663 45512 42708 45540
rect 42702 45500 42708 45512
rect 42760 45500 42766 45552
rect 43990 45540 43996 45552
rect 43364 45512 43996 45540
rect 10560 45444 12572 45472
rect 13633 45475 13691 45481
rect 10560 45432 10566 45444
rect 13633 45441 13645 45475
rect 13679 45472 13691 45475
rect 20717 45475 20775 45481
rect 13679 45444 16574 45472
rect 13679 45441 13691 45444
rect 13633 45435 13691 45441
rect 1949 45407 2007 45413
rect 1949 45373 1961 45407
rect 1995 45404 2007 45407
rect 2774 45404 2780 45416
rect 1995 45376 2780 45404
rect 1995 45373 2007 45376
rect 1949 45367 2007 45373
rect 2774 45364 2780 45376
rect 2832 45364 2838 45416
rect 2958 45404 2964 45416
rect 2919 45376 2964 45404
rect 2958 45364 2964 45376
rect 3016 45364 3022 45416
rect 16546 45336 16574 45444
rect 20717 45441 20729 45475
rect 20763 45441 20775 45475
rect 24872 45472 24900 45500
rect 25317 45475 25375 45481
rect 25317 45472 25329 45475
rect 24872 45444 25329 45472
rect 20717 45435 20775 45441
rect 25317 45441 25329 45444
rect 25363 45472 25375 45475
rect 26050 45472 26056 45484
rect 25363 45444 26056 45472
rect 25363 45441 25375 45444
rect 25317 45435 25375 45441
rect 20732 45404 20760 45435
rect 26050 45432 26056 45444
rect 26108 45432 26114 45484
rect 41325 45475 41383 45481
rect 41325 45441 41337 45475
rect 41371 45472 41383 45475
rect 42613 45475 42671 45481
rect 42613 45472 42625 45475
rect 41371 45444 42625 45472
rect 41371 45441 41383 45444
rect 41325 45435 41383 45441
rect 42613 45441 42625 45444
rect 42659 45472 42671 45475
rect 43364 45472 43392 45512
rect 43990 45500 43996 45512
rect 44048 45500 44054 45552
rect 45572 45540 45600 45580
rect 46198 45568 46204 45620
rect 46256 45608 46262 45620
rect 46256 45580 47992 45608
rect 46256 45568 46262 45580
rect 47964 45549 47992 45580
rect 47949 45543 48007 45549
rect 45572 45512 46060 45540
rect 42659 45444 43392 45472
rect 43901 45475 43959 45481
rect 42659 45441 42671 45444
rect 42613 45435 42671 45441
rect 43901 45441 43913 45475
rect 43947 45472 43959 45475
rect 44174 45472 44180 45484
rect 43947 45444 44180 45472
rect 43947 45441 43959 45444
rect 43901 45435 43959 45441
rect 44174 45432 44180 45444
rect 44232 45432 44238 45484
rect 27338 45404 27344 45416
rect 20732 45376 27344 45404
rect 27338 45364 27344 45376
rect 27396 45364 27402 45416
rect 38654 45404 38660 45416
rect 38615 45376 38660 45404
rect 38654 45364 38660 45376
rect 38712 45364 38718 45416
rect 38838 45404 38844 45416
rect 38799 45376 38844 45404
rect 38838 45364 38844 45376
rect 38896 45364 38902 45416
rect 39850 45404 39856 45416
rect 39811 45376 39856 45404
rect 39850 45364 39856 45376
rect 39908 45364 39914 45416
rect 43441 45407 43499 45413
rect 43441 45373 43453 45407
rect 43487 45404 43499 45407
rect 44637 45407 44695 45413
rect 44637 45404 44649 45407
rect 43487 45376 44649 45404
rect 43487 45373 43499 45376
rect 43441 45367 43499 45373
rect 44637 45373 44649 45376
rect 44683 45373 44695 45407
rect 44637 45367 44695 45373
rect 44821 45407 44879 45413
rect 44821 45373 44833 45407
rect 44867 45404 44879 45407
rect 45094 45404 45100 45416
rect 44867 45376 45100 45404
rect 44867 45373 44879 45376
rect 44821 45367 44879 45373
rect 45094 45364 45100 45376
rect 45152 45364 45158 45416
rect 46032 45413 46060 45512
rect 47949 45509 47961 45543
rect 47995 45509 48007 45543
rect 47949 45503 48007 45509
rect 46017 45407 46075 45413
rect 46017 45373 46029 45407
rect 46063 45373 46075 45407
rect 46017 45367 46075 45373
rect 40678 45336 40684 45348
rect 16546 45308 40684 45336
rect 40678 45296 40684 45308
rect 40736 45296 40742 45348
rect 42794 45296 42800 45348
rect 42852 45336 42858 45348
rect 42852 45308 44220 45336
rect 42852 45296 42858 45308
rect 44082 45268 44088 45280
rect 44043 45240 44088 45268
rect 44082 45228 44088 45240
rect 44140 45228 44146 45280
rect 44192 45268 44220 45308
rect 44266 45296 44272 45348
rect 44324 45336 44330 45348
rect 47578 45336 47584 45348
rect 44324 45308 47584 45336
rect 44324 45296 44330 45308
rect 47578 45296 47584 45308
rect 47636 45296 47642 45348
rect 48041 45271 48099 45277
rect 48041 45268 48053 45271
rect 44192 45240 48053 45268
rect 48041 45237 48053 45240
rect 48087 45237 48099 45271
rect 48041 45231 48099 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 38838 45064 38844 45076
rect 38799 45036 38844 45064
rect 38838 45024 38844 45036
rect 38896 45024 38902 45076
rect 40405 45067 40463 45073
rect 40405 45033 40417 45067
rect 40451 45064 40463 45067
rect 41230 45064 41236 45076
rect 40451 45036 41236 45064
rect 40451 45033 40463 45036
rect 40405 45027 40463 45033
rect 41230 45024 41236 45036
rect 41288 45024 41294 45076
rect 45094 45064 45100 45076
rect 45055 45036 45100 45064
rect 45094 45024 45100 45036
rect 45152 45024 45158 45076
rect 45741 45067 45799 45073
rect 45741 45033 45753 45067
rect 45787 45064 45799 45067
rect 46474 45064 46480 45076
rect 45787 45036 46480 45064
rect 45787 45033 45799 45036
rect 45741 45027 45799 45033
rect 46474 45024 46480 45036
rect 46532 45024 46538 45076
rect 44361 44999 44419 45005
rect 44361 44965 44373 44999
rect 44407 44996 44419 44999
rect 45370 44996 45376 45008
rect 44407 44968 45376 44996
rect 44407 44965 44419 44968
rect 44361 44959 44419 44965
rect 45370 44956 45376 44968
rect 45428 44956 45434 45008
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 47026 44928 47032 44940
rect 46339 44900 47032 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 47026 44888 47032 44900
rect 47084 44888 47090 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 28626 44820 28632 44872
rect 28684 44860 28690 44872
rect 29549 44863 29607 44869
rect 29549 44860 29561 44863
rect 28684 44832 29561 44860
rect 28684 44820 28690 44832
rect 29549 44829 29561 44832
rect 29595 44829 29607 44863
rect 29549 44823 29607 44829
rect 38749 44863 38807 44869
rect 38749 44829 38761 44863
rect 38795 44860 38807 44863
rect 40034 44860 40040 44872
rect 38795 44832 40040 44860
rect 38795 44829 38807 44832
rect 38749 44823 38807 44829
rect 40034 44820 40040 44832
rect 40092 44820 40098 44872
rect 40310 44860 40316 44872
rect 40271 44832 40316 44860
rect 40310 44820 40316 44832
rect 40368 44820 40374 44872
rect 44266 44860 44272 44872
rect 44227 44832 44272 44860
rect 44266 44820 44272 44832
rect 44324 44820 44330 44872
rect 45002 44860 45008 44872
rect 44963 44832 45008 44860
rect 45002 44820 45008 44832
rect 45060 44820 45066 44872
rect 45649 44863 45707 44869
rect 45649 44829 45661 44863
rect 45695 44829 45707 44863
rect 45649 44823 45707 44829
rect 29641 44727 29699 44733
rect 29641 44693 29653 44727
rect 29687 44724 29699 44727
rect 38654 44724 38660 44736
rect 29687 44696 38660 44724
rect 29687 44693 29699 44696
rect 29641 44687 29699 44693
rect 38654 44684 38660 44696
rect 38712 44684 38718 44736
rect 45664 44724 45692 44823
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 47670 44792 47676 44804
rect 46523 44764 47676 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 47670 44752 47676 44764
rect 47728 44752 47734 44804
rect 45830 44724 45836 44736
rect 45664 44696 45836 44724
rect 45830 44684 45836 44696
rect 45888 44724 45894 44736
rect 46750 44724 46756 44736
rect 45888 44696 46756 44724
rect 45888 44684 45894 44696
rect 46750 44684 46756 44696
rect 46808 44684 46814 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 45462 44480 45468 44532
rect 45520 44520 45526 44532
rect 46293 44523 46351 44529
rect 46293 44520 46305 44523
rect 45520 44492 46305 44520
rect 45520 44480 45526 44492
rect 46293 44489 46305 44492
rect 46339 44489 46351 44523
rect 47670 44520 47676 44532
rect 47631 44492 47676 44520
rect 46293 44483 46351 44489
rect 47670 44480 47676 44492
rect 47728 44480 47734 44532
rect 40678 44412 40684 44464
rect 40736 44452 40742 44464
rect 40736 44424 46612 44452
rect 40736 44412 40742 44424
rect 46584 44396 46612 44424
rect 20070 44344 20076 44396
rect 20128 44384 20134 44396
rect 45097 44387 45155 44393
rect 20128 44356 26234 44384
rect 20128 44344 20134 44356
rect 26206 44316 26234 44356
rect 45097 44353 45109 44387
rect 45143 44384 45155 44387
rect 45186 44384 45192 44396
rect 45143 44356 45192 44384
rect 45143 44353 45155 44356
rect 45097 44347 45155 44353
rect 45186 44344 45192 44356
rect 45244 44344 45250 44396
rect 45738 44384 45744 44396
rect 45699 44356 45744 44384
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46201 44387 46259 44393
rect 46201 44384 46213 44387
rect 45940 44356 46213 44384
rect 45940 44328 45968 44356
rect 46201 44353 46213 44356
rect 46247 44353 46259 44387
rect 46201 44347 46259 44353
rect 46566 44344 46572 44396
rect 46624 44384 46630 44396
rect 46845 44387 46903 44393
rect 46845 44384 46857 44387
rect 46624 44356 46857 44384
rect 46624 44344 46630 44356
rect 46845 44353 46857 44356
rect 46891 44384 46903 44387
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 46891 44356 47593 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 45922 44316 45928 44328
rect 26206 44288 45928 44316
rect 45922 44276 45928 44288
rect 45980 44276 45986 44328
rect 46934 44180 46940 44192
rect 46895 44152 46940 44180
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 46934 43840 46940 43852
rect 46523 43812 46940 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 46934 43800 46940 43812
rect 46992 43800 46998 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 1670 43228 1676 43240
rect 1631 43200 1676 43228
rect 1670 43188 1676 43200
rect 1728 43188 1734 43240
rect 46290 43188 46296 43240
rect 46348 43228 46354 43240
rect 47765 43231 47823 43237
rect 47765 43228 47777 43231
rect 46348 43200 47777 43228
rect 46348 43188 46354 43200
rect 47765 43197 47777 43200
rect 47811 43197 47823 43231
rect 47765 43191 47823 43197
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46290 42684 46296 42696
rect 46251 42656 46296 42684
rect 46290 42644 46296 42656
rect 46348 42644 46354 42696
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 46290 42168 46296 42220
rect 46348 42208 46354 42220
rect 47029 42211 47087 42217
rect 47029 42208 47041 42211
rect 46348 42180 47041 42208
rect 46348 42168 46354 42180
rect 47029 42177 47041 42180
rect 47075 42177 47087 42211
rect 47578 42208 47584 42220
rect 47539 42180 47584 42208
rect 47029 42171 47087 42177
rect 47578 42168 47584 42180
rect 47636 42168 47642 42220
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46477 41531 46535 41537
rect 46477 41497 46489 41531
rect 46523 41528 46535 41531
rect 46934 41528 46940 41540
rect 46523 41500 46940 41528
rect 46523 41497 46535 41500
rect 46477 41491 46535 41497
rect 46934 41488 46940 41500
rect 46992 41488 46998 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2225 41259 2283 41265
rect 2225 41256 2237 41259
rect 1636 41228 2237 41256
rect 1636 41216 1642 41228
rect 2225 41225 2237 41228
rect 2271 41225 2283 41259
rect 46934 41256 46940 41268
rect 46895 41228 46940 41256
rect 2225 41219 2283 41225
rect 46934 41216 46940 41228
rect 46992 41216 46998 41268
rect 2130 41120 2136 41132
rect 2091 41092 2136 41120
rect 2130 41080 2136 41092
rect 2188 41120 2194 41132
rect 20070 41120 20076 41132
rect 2188 41092 20076 41120
rect 2188 41080 2194 41092
rect 20070 41080 20076 41092
rect 20128 41080 20134 41132
rect 46750 41080 46756 41132
rect 46808 41120 46814 41132
rect 46845 41123 46903 41129
rect 46845 41120 46857 41123
rect 46808 41092 46857 41120
rect 46808 41080 46814 41092
rect 46845 41089 46857 41092
rect 46891 41089 46903 41123
rect 46845 41083 46903 41089
rect 47949 41123 48007 41129
rect 47949 41089 47961 41123
rect 47995 41120 48007 41123
rect 48038 41120 48044 41132
rect 47995 41092 48044 41120
rect 47995 41089 48007 41092
rect 47949 41083 48007 41089
rect 48038 41080 48044 41092
rect 48096 41080 48102 41132
rect 47946 40876 47952 40928
rect 48004 40916 48010 40928
rect 48041 40919 48099 40925
rect 48041 40916 48053 40919
rect 48004 40888 48053 40916
rect 48004 40876 48010 40888
rect 48041 40885 48053 40888
rect 48087 40885 48099 40919
rect 48041 40879 48099 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 1394 40508 1400 40520
rect 1355 40480 1400 40508
rect 1394 40468 1400 40480
rect 1452 40468 1458 40520
rect 1581 40375 1639 40381
rect 1581 40341 1593 40375
rect 1627 40372 1639 40375
rect 1762 40372 1768 40384
rect 1627 40344 1768 40372
rect 1627 40341 1639 40344
rect 1581 40335 1639 40341
rect 1762 40332 1768 40344
rect 1820 40332 1826 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 46934 39352 46940 39364
rect 46523 39324 46940 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 46934 39312 46940 39324
rect 46992 39312 46998 39364
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 3326 39040 3332 39092
rect 3384 39080 3390 39092
rect 7558 39080 7564 39092
rect 3384 39052 7564 39080
rect 3384 39040 3390 39052
rect 7558 39040 7564 39052
rect 7616 39040 7622 39092
rect 26142 39080 26148 39092
rect 26055 39052 26148 39080
rect 26142 39040 26148 39052
rect 26200 39080 26206 39092
rect 46934 39080 46940 39092
rect 26200 39052 27016 39080
rect 46895 39052 46940 39080
rect 26200 39040 26206 39052
rect 25314 38904 25320 38956
rect 25372 38944 25378 38956
rect 25958 38944 25964 38956
rect 25372 38916 25964 38944
rect 25372 38904 25378 38916
rect 25958 38904 25964 38916
rect 26016 38904 26022 38956
rect 26988 38953 27016 39052
rect 46934 39040 46940 39052
rect 46992 39040 46998 39092
rect 26973 38947 27031 38953
rect 26973 38913 26985 38947
rect 27019 38913 27031 38947
rect 26973 38907 27031 38913
rect 46014 38904 46020 38956
rect 46072 38944 46078 38956
rect 46845 38947 46903 38953
rect 46845 38944 46857 38947
rect 46072 38916 46857 38944
rect 46072 38904 46078 38916
rect 46845 38913 46857 38916
rect 46891 38913 46903 38947
rect 47670 38944 47676 38956
rect 47631 38916 47676 38944
rect 46845 38907 46903 38913
rect 47670 38904 47676 38916
rect 47728 38904 47734 38956
rect 8202 38836 8208 38888
rect 8260 38876 8266 38888
rect 27341 38879 27399 38885
rect 27341 38876 27353 38879
rect 8260 38848 27353 38876
rect 8260 38836 8266 38848
rect 27341 38845 27353 38848
rect 27387 38876 27399 38879
rect 38102 38876 38108 38888
rect 27387 38848 38108 38876
rect 27387 38845 27399 38848
rect 27341 38839 27399 38845
rect 38102 38836 38108 38848
rect 38160 38836 38166 38888
rect 47854 38876 47860 38888
rect 45526 38848 47860 38876
rect 25958 38768 25964 38820
rect 26016 38808 26022 38820
rect 45526 38808 45554 38848
rect 47854 38836 47860 38848
rect 47912 38836 47918 38888
rect 26016 38780 45554 38808
rect 26016 38768 26022 38780
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 26142 38332 26148 38344
rect 26103 38304 26148 38332
rect 26142 38292 26148 38304
rect 26200 38292 26206 38344
rect 46934 38292 46940 38344
rect 46992 38332 46998 38344
rect 47673 38335 47731 38341
rect 47673 38332 47685 38335
rect 46992 38304 47685 38332
rect 46992 38292 46998 38304
rect 47673 38301 47685 38304
rect 47719 38301 47731 38335
rect 47673 38295 47731 38301
rect 26326 38156 26332 38208
rect 26384 38196 26390 38208
rect 27433 38199 27491 38205
rect 27433 38196 27445 38199
rect 26384 38168 27445 38196
rect 26384 38156 26390 38168
rect 27433 38165 27445 38168
rect 27479 38196 27491 38199
rect 44266 38196 44272 38208
rect 27479 38168 44272 38196
rect 27479 38165 27491 38168
rect 27433 38159 27491 38165
rect 44266 38156 44272 38168
rect 44324 38156 44330 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 25777 37859 25835 37865
rect 25777 37825 25789 37859
rect 25823 37856 25835 37859
rect 26142 37856 26148 37868
rect 25823 37828 26148 37856
rect 25823 37825 25835 37828
rect 25777 37819 25835 37825
rect 26142 37816 26148 37828
rect 26200 37856 26206 37868
rect 26973 37859 27031 37865
rect 26973 37856 26985 37859
rect 26200 37828 26985 37856
rect 26200 37816 26206 37828
rect 26973 37825 26985 37828
rect 27019 37825 27031 37859
rect 47578 37856 47584 37868
rect 26973 37819 27031 37825
rect 35866 37828 47584 37856
rect 25406 37748 25412 37800
rect 25464 37788 25470 37800
rect 26050 37788 26056 37800
rect 25464 37760 26056 37788
rect 25464 37748 25470 37760
rect 26050 37748 26056 37760
rect 26108 37748 26114 37800
rect 26786 37748 26792 37800
rect 26844 37788 26850 37800
rect 27338 37788 27344 37800
rect 26844 37760 27344 37788
rect 26844 37748 26850 37760
rect 27338 37748 27344 37760
rect 27396 37788 27402 37800
rect 35866 37788 35894 37828
rect 47578 37816 47584 37828
rect 47636 37816 47642 37868
rect 27396 37760 35894 37788
rect 27396 37748 27402 37760
rect 47670 37652 47676 37664
rect 47631 37624 47676 37652
rect 47670 37612 47676 37624
rect 47728 37612 47734 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 26142 37244 26148 37256
rect 26103 37216 26148 37244
rect 26142 37204 26148 37216
rect 26200 37204 26206 37256
rect 46293 37247 46351 37253
rect 46293 37213 46305 37247
rect 46339 37213 46351 37247
rect 46293 37207 46351 37213
rect 26694 37136 26700 37188
rect 26752 37176 26758 37188
rect 26881 37179 26939 37185
rect 26881 37176 26893 37179
rect 26752 37148 26893 37176
rect 26752 37136 26758 37148
rect 26881 37145 26893 37148
rect 26927 37176 26939 37179
rect 40310 37176 40316 37188
rect 26927 37148 40316 37176
rect 26927 37145 26939 37148
rect 26881 37139 26939 37145
rect 40310 37136 40316 37148
rect 40368 37136 40374 37188
rect 46308 37108 46336 37207
rect 46477 37179 46535 37185
rect 46477 37145 46489 37179
rect 46523 37176 46535 37179
rect 47670 37176 47676 37188
rect 46523 37148 47676 37176
rect 46523 37145 46535 37148
rect 46477 37139 46535 37145
rect 47670 37136 47676 37148
rect 47728 37136 47734 37188
rect 46934 37108 46940 37120
rect 46308 37080 46940 37108
rect 46934 37068 46940 37080
rect 46992 37068 46998 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 26237 36839 26295 36845
rect 26237 36805 26249 36839
rect 26283 36836 26295 36839
rect 27522 36836 27528 36848
rect 26283 36808 27528 36836
rect 26283 36805 26295 36808
rect 26237 36799 26295 36805
rect 27522 36796 27528 36808
rect 27580 36796 27586 36848
rect 12434 36728 12440 36780
rect 12492 36768 12498 36780
rect 26053 36771 26111 36777
rect 26053 36768 26065 36771
rect 12492 36740 26065 36768
rect 12492 36728 12498 36740
rect 26053 36737 26065 36740
rect 26099 36737 26111 36771
rect 26053 36731 26111 36737
rect 27341 36771 27399 36777
rect 27341 36737 27353 36771
rect 27387 36768 27399 36771
rect 27387 36740 28120 36768
rect 27387 36737 27399 36740
rect 27341 36731 27399 36737
rect 26970 36660 26976 36712
rect 27028 36700 27034 36712
rect 27433 36703 27491 36709
rect 27433 36700 27445 36703
rect 27028 36672 27445 36700
rect 27028 36660 27034 36672
rect 27433 36669 27445 36672
rect 27479 36669 27491 36703
rect 27433 36663 27491 36669
rect 27522 36660 27528 36712
rect 27580 36700 27586 36712
rect 27580 36672 27625 36700
rect 27580 36660 27586 36672
rect 26418 36564 26424 36576
rect 26379 36536 26424 36564
rect 26418 36524 26424 36536
rect 26476 36524 26482 36576
rect 26510 36524 26516 36576
rect 26568 36564 26574 36576
rect 28092 36573 28120 36740
rect 26973 36567 27031 36573
rect 26973 36564 26985 36567
rect 26568 36536 26985 36564
rect 26568 36524 26574 36536
rect 26973 36533 26985 36536
rect 27019 36533 27031 36567
rect 26973 36527 27031 36533
rect 28077 36567 28135 36573
rect 28077 36533 28089 36567
rect 28123 36564 28135 36567
rect 45554 36564 45560 36576
rect 28123 36536 45560 36564
rect 28123 36533 28135 36536
rect 28077 36527 28135 36533
rect 45554 36524 45560 36536
rect 45612 36524 45618 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 26970 36360 26976 36372
rect 26931 36332 26976 36360
rect 26970 36320 26976 36332
rect 27028 36320 27034 36372
rect 2774 36224 2780 36236
rect 2735 36196 2780 36224
rect 2774 36184 2780 36196
rect 2832 36184 2838 36236
rect 26510 36224 26516 36236
rect 23676 36196 26516 36224
rect 1394 36156 1400 36168
rect 1355 36128 1400 36156
rect 1394 36116 1400 36128
rect 1452 36116 1458 36168
rect 23676 36165 23704 36196
rect 26510 36184 26516 36196
rect 26568 36184 26574 36236
rect 26697 36227 26755 36233
rect 26697 36193 26709 36227
rect 26743 36224 26755 36227
rect 27430 36224 27436 36236
rect 26743 36196 27436 36224
rect 26743 36193 26755 36196
rect 26697 36187 26755 36193
rect 27430 36184 27436 36196
rect 27488 36184 27494 36236
rect 23661 36159 23719 36165
rect 23661 36125 23673 36159
rect 23707 36125 23719 36159
rect 23661 36119 23719 36125
rect 25685 36159 25743 36165
rect 25685 36125 25697 36159
rect 25731 36156 25743 36159
rect 25774 36156 25780 36168
rect 25731 36128 25780 36156
rect 25731 36125 25743 36128
rect 25685 36119 25743 36125
rect 25774 36116 25780 36128
rect 25832 36116 25838 36168
rect 26602 36156 26608 36168
rect 26563 36128 26608 36156
rect 26602 36116 26608 36128
rect 26660 36116 26666 36168
rect 1581 36091 1639 36097
rect 1581 36057 1593 36091
rect 1627 36088 1639 36091
rect 2222 36088 2228 36100
rect 1627 36060 2228 36088
rect 1627 36057 1639 36060
rect 1581 36051 1639 36057
rect 2222 36048 2228 36060
rect 2280 36048 2286 36100
rect 23474 36020 23480 36032
rect 23435 35992 23480 36020
rect 23474 35980 23480 35992
rect 23532 35980 23538 36032
rect 25682 35980 25688 36032
rect 25740 36020 25746 36032
rect 25777 36023 25835 36029
rect 25777 36020 25789 36023
rect 25740 35992 25789 36020
rect 25740 35980 25746 35992
rect 25777 35989 25789 35992
rect 25823 35989 25835 36023
rect 25777 35983 25835 35989
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 24213 35819 24271 35825
rect 24213 35785 24225 35819
rect 24259 35816 24271 35819
rect 26602 35816 26608 35828
rect 24259 35788 26608 35816
rect 24259 35785 24271 35788
rect 24213 35779 24271 35785
rect 26602 35776 26608 35788
rect 26660 35776 26666 35828
rect 22830 35708 22836 35760
rect 22888 35748 22894 35760
rect 22888 35720 23230 35748
rect 22888 35708 22894 35720
rect 25682 35708 25688 35760
rect 25740 35708 25746 35760
rect 30926 35708 30932 35760
rect 30984 35708 30990 35760
rect 1394 35640 1400 35692
rect 1452 35680 1458 35692
rect 2041 35683 2099 35689
rect 2041 35680 2053 35683
rect 1452 35652 2053 35680
rect 1452 35640 1458 35652
rect 2041 35649 2053 35652
rect 2087 35649 2099 35683
rect 2041 35643 2099 35649
rect 26418 35640 26424 35692
rect 26476 35680 26482 35692
rect 27157 35683 27215 35689
rect 27157 35680 27169 35683
rect 26476 35652 27169 35680
rect 26476 35640 26482 35652
rect 27157 35649 27169 35652
rect 27203 35649 27215 35683
rect 27157 35643 27215 35649
rect 22465 35615 22523 35621
rect 22465 35581 22477 35615
rect 22511 35581 22523 35615
rect 22465 35575 22523 35581
rect 22741 35615 22799 35621
rect 22741 35581 22753 35615
rect 22787 35612 22799 35615
rect 23474 35612 23480 35624
rect 22787 35584 23480 35612
rect 22787 35581 22799 35584
rect 22741 35575 22799 35581
rect 22480 35476 22508 35575
rect 23474 35572 23480 35584
rect 23532 35572 23538 35624
rect 24670 35612 24676 35624
rect 24631 35584 24676 35612
rect 24670 35572 24676 35584
rect 24728 35572 24734 35624
rect 24946 35612 24952 35624
rect 24907 35584 24952 35612
rect 24946 35572 24952 35584
rect 25004 35572 25010 35624
rect 27433 35615 27491 35621
rect 27433 35581 27445 35615
rect 27479 35612 27491 35615
rect 28442 35612 28448 35624
rect 27479 35584 28448 35612
rect 27479 35581 27491 35584
rect 27433 35575 27491 35581
rect 28442 35572 28448 35584
rect 28500 35572 28506 35624
rect 29641 35615 29699 35621
rect 29641 35581 29653 35615
rect 29687 35581 29699 35615
rect 29914 35612 29920 35624
rect 29875 35584 29920 35612
rect 29641 35575 29699 35581
rect 23474 35476 23480 35488
rect 22480 35448 23480 35476
rect 23474 35436 23480 35448
rect 23532 35476 23538 35488
rect 24670 35476 24676 35488
rect 23532 35448 24676 35476
rect 23532 35436 23538 35448
rect 24670 35436 24676 35448
rect 24728 35436 24734 35488
rect 26421 35479 26479 35485
rect 26421 35445 26433 35479
rect 26467 35476 26479 35479
rect 26510 35476 26516 35488
rect 26467 35448 26516 35476
rect 26467 35445 26479 35448
rect 26421 35439 26479 35445
rect 26510 35436 26516 35448
rect 26568 35436 26574 35488
rect 26970 35476 26976 35488
rect 26931 35448 26976 35476
rect 26970 35436 26976 35448
rect 27028 35436 27034 35488
rect 27341 35479 27399 35485
rect 27341 35445 27353 35479
rect 27387 35476 27399 35479
rect 27430 35476 27436 35488
rect 27387 35448 27436 35476
rect 27387 35445 27399 35448
rect 27341 35439 27399 35445
rect 27430 35436 27436 35448
rect 27488 35436 27494 35488
rect 29656 35476 29684 35575
rect 29914 35572 29920 35584
rect 29972 35572 29978 35624
rect 30282 35572 30288 35624
rect 30340 35612 30346 35624
rect 31389 35615 31447 35621
rect 31389 35612 31401 35615
rect 30340 35584 31401 35612
rect 30340 35572 30346 35584
rect 31389 35581 31401 35584
rect 31435 35581 31447 35615
rect 31389 35575 31447 35581
rect 31110 35476 31116 35488
rect 29656 35448 31116 35476
rect 31110 35436 31116 35448
rect 31168 35436 31174 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 2222 35272 2228 35284
rect 2183 35244 2228 35272
rect 2222 35232 2228 35244
rect 2280 35232 2286 35284
rect 22830 35272 22836 35284
rect 22791 35244 22836 35272
rect 22830 35232 22836 35244
rect 22888 35232 22894 35284
rect 24946 35232 24952 35284
rect 25004 35272 25010 35284
rect 25869 35275 25927 35281
rect 25869 35272 25881 35275
rect 25004 35244 25881 35272
rect 25004 35232 25010 35244
rect 25869 35241 25881 35244
rect 25915 35241 25927 35275
rect 29641 35275 29699 35281
rect 25869 35235 25927 35241
rect 25976 35244 27292 35272
rect 24670 35164 24676 35216
rect 24728 35204 24734 35216
rect 25976 35204 26004 35244
rect 26418 35204 26424 35216
rect 24728 35176 26004 35204
rect 26068 35176 26424 35204
rect 24728 35164 24734 35176
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35028 1642 35080
rect 2133 35071 2191 35077
rect 2133 35037 2145 35071
rect 2179 35068 2191 35071
rect 2222 35068 2228 35080
rect 2179 35040 2228 35068
rect 2179 35037 2191 35040
rect 2133 35031 2191 35037
rect 2222 35028 2228 35040
rect 2280 35028 2286 35080
rect 22002 35028 22008 35080
rect 22060 35068 22066 35080
rect 22741 35071 22799 35077
rect 22741 35068 22753 35071
rect 22060 35040 22753 35068
rect 22060 35028 22066 35040
rect 22741 35037 22753 35040
rect 22787 35037 22799 35071
rect 24486 35068 24492 35080
rect 24447 35040 24492 35068
rect 22741 35031 22799 35037
rect 24486 35028 24492 35040
rect 24544 35028 24550 35080
rect 26068 35077 26096 35176
rect 26418 35164 26424 35176
rect 26476 35164 26482 35216
rect 27264 35145 27292 35244
rect 29641 35241 29653 35275
rect 29687 35272 29699 35275
rect 29914 35272 29920 35284
rect 29687 35244 29920 35272
rect 29687 35241 29699 35244
rect 29641 35235 29699 35241
rect 29914 35232 29920 35244
rect 29972 35232 29978 35284
rect 30190 35272 30196 35284
rect 30151 35244 30196 35272
rect 30190 35232 30196 35244
rect 30248 35272 30254 35284
rect 30561 35275 30619 35281
rect 30561 35272 30573 35275
rect 30248 35244 30573 35272
rect 30248 35232 30254 35244
rect 30561 35241 30573 35244
rect 30607 35241 30619 35275
rect 30561 35235 30619 35241
rect 30837 35275 30895 35281
rect 30837 35241 30849 35275
rect 30883 35272 30895 35275
rect 30926 35272 30932 35284
rect 30883 35244 30932 35272
rect 30883 35241 30895 35244
rect 30837 35235 30895 35241
rect 30926 35232 30932 35244
rect 30984 35232 30990 35284
rect 27249 35139 27307 35145
rect 27249 35105 27261 35139
rect 27295 35105 27307 35139
rect 27249 35099 27307 35105
rect 29730 35096 29736 35148
rect 29788 35136 29794 35148
rect 30285 35139 30343 35145
rect 30285 35136 30297 35139
rect 29788 35108 30297 35136
rect 29788 35096 29794 35108
rect 30285 35105 30297 35108
rect 30331 35105 30343 35139
rect 30285 35099 30343 35105
rect 26053 35071 26111 35077
rect 26053 35037 26065 35071
rect 26099 35037 26111 35071
rect 26053 35031 26111 35037
rect 26145 35071 26203 35077
rect 26145 35037 26157 35071
rect 26191 35037 26203 35071
rect 26145 35031 26203 35037
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35037 26295 35071
rect 26237 35031 26295 35037
rect 26329 35071 26387 35077
rect 26329 35037 26341 35071
rect 26375 35068 26387 35071
rect 26970 35068 26976 35080
rect 26375 35040 26976 35068
rect 26375 35037 26387 35040
rect 26329 35031 26387 35037
rect 1397 34935 1455 34941
rect 1397 34901 1409 34935
rect 1443 34932 1455 34935
rect 1486 34932 1492 34944
rect 1443 34904 1492 34932
rect 1443 34901 1455 34904
rect 1397 34895 1455 34901
rect 1486 34892 1492 34904
rect 1544 34892 1550 34944
rect 24673 34935 24731 34941
rect 24673 34901 24685 34935
rect 24719 34932 24731 34935
rect 24946 34932 24952 34944
rect 24719 34904 24952 34932
rect 24719 34901 24731 34904
rect 24673 34895 24731 34901
rect 24946 34892 24952 34904
rect 25004 34892 25010 34944
rect 26160 34932 26188 35031
rect 26252 35000 26280 35031
rect 26970 35028 26976 35040
rect 27028 35028 27034 35080
rect 29822 35071 29880 35077
rect 29822 35037 29834 35071
rect 29868 35068 29880 35071
rect 30098 35068 30104 35080
rect 29868 35040 30104 35068
rect 29868 35037 29880 35040
rect 29822 35031 29880 35037
rect 30098 35028 30104 35040
rect 30156 35028 30162 35080
rect 30745 35071 30803 35077
rect 30745 35037 30757 35071
rect 30791 35068 30803 35071
rect 31573 35071 31631 35077
rect 31573 35068 31585 35071
rect 30791 35040 31585 35068
rect 30791 35037 30803 35040
rect 30745 35031 30803 35037
rect 31573 35037 31585 35040
rect 31619 35037 31631 35071
rect 48130 35068 48136 35080
rect 48091 35040 48136 35068
rect 31573 35031 31631 35037
rect 26510 35000 26516 35012
rect 26252 34972 26516 35000
rect 26510 34960 26516 34972
rect 26568 34960 26574 35012
rect 27525 35003 27583 35009
rect 27525 34969 27537 35003
rect 27571 35000 27583 35003
rect 27798 35000 27804 35012
rect 27571 34972 27804 35000
rect 27571 34969 27583 34972
rect 27525 34963 27583 34969
rect 27798 34960 27804 34972
rect 27856 34960 27862 35012
rect 28810 35000 28816 35012
rect 28750 34972 28816 35000
rect 28810 34960 28816 34972
rect 28868 34960 28874 35012
rect 28902 34960 28908 35012
rect 28960 35000 28966 35012
rect 30760 35000 30788 35031
rect 48130 35028 48136 35040
rect 48188 35028 48194 35080
rect 28960 34972 30788 35000
rect 28960 34960 28966 34972
rect 27338 34932 27344 34944
rect 26160 34904 27344 34932
rect 27338 34892 27344 34904
rect 27396 34892 27402 34944
rect 28997 34935 29055 34941
rect 28997 34901 29009 34935
rect 29043 34932 29055 34935
rect 29178 34932 29184 34944
rect 29043 34904 29184 34932
rect 29043 34901 29055 34904
rect 28997 34895 29055 34901
rect 29178 34892 29184 34904
rect 29236 34892 29242 34944
rect 29822 34932 29828 34944
rect 29783 34904 29828 34932
rect 29822 34892 29828 34904
rect 29880 34892 29886 34944
rect 31665 34935 31723 34941
rect 31665 34901 31677 34935
rect 31711 34932 31723 34935
rect 31846 34932 31852 34944
rect 31711 34904 31852 34932
rect 31711 34901 31723 34904
rect 31665 34895 31723 34901
rect 31846 34892 31852 34904
rect 31904 34892 31910 34944
rect 47118 34892 47124 34944
rect 47176 34932 47182 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47176 34904 47961 34932
rect 47176 34892 47182 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 23474 34728 23480 34740
rect 21836 34700 23480 34728
rect 21836 34601 21864 34700
rect 23474 34688 23480 34700
rect 23532 34688 23538 34740
rect 26973 34731 27031 34737
rect 26973 34697 26985 34731
rect 27019 34728 27031 34731
rect 27982 34728 27988 34740
rect 27019 34700 27988 34728
rect 27019 34697 27031 34700
rect 26973 34691 27031 34697
rect 27982 34688 27988 34700
rect 28040 34688 28046 34740
rect 28810 34728 28816 34740
rect 28771 34700 28816 34728
rect 28810 34688 28816 34700
rect 28868 34688 28874 34740
rect 30098 34728 30104 34740
rect 30059 34700 30104 34728
rect 30098 34688 30104 34700
rect 30156 34688 30162 34740
rect 26510 34620 26516 34672
rect 26568 34660 26574 34672
rect 27249 34663 27307 34669
rect 27249 34660 27261 34663
rect 26568 34632 27261 34660
rect 26568 34620 26574 34632
rect 27249 34629 27261 34632
rect 27295 34629 27307 34663
rect 30653 34663 30711 34669
rect 30653 34660 30665 34663
rect 27249 34623 27307 34629
rect 30024 34632 30665 34660
rect 20717 34595 20775 34601
rect 20717 34561 20729 34595
rect 20763 34561 20775 34595
rect 20717 34555 20775 34561
rect 21821 34595 21879 34601
rect 21821 34561 21833 34595
rect 21867 34561 21879 34595
rect 21821 34555 21879 34561
rect 20732 34524 20760 34555
rect 23198 34552 23204 34604
rect 23256 34552 23262 34604
rect 24765 34595 24823 34601
rect 24765 34561 24777 34595
rect 24811 34592 24823 34595
rect 24946 34592 24952 34604
rect 24811 34564 24952 34592
rect 24811 34561 24823 34564
rect 24765 34555 24823 34561
rect 24946 34552 24952 34564
rect 25004 34592 25010 34604
rect 25774 34592 25780 34604
rect 25004 34564 25780 34592
rect 25004 34552 25010 34564
rect 25774 34552 25780 34564
rect 25832 34592 25838 34604
rect 25832 34564 26832 34592
rect 25832 34552 25838 34564
rect 23566 34524 23572 34536
rect 20732 34496 23572 34524
rect 23566 34484 23572 34496
rect 23624 34524 23630 34536
rect 24486 34524 24492 34536
rect 23624 34496 24492 34524
rect 23624 34484 23630 34496
rect 24486 34484 24492 34496
rect 24544 34484 24550 34536
rect 24857 34527 24915 34533
rect 24857 34493 24869 34527
rect 24903 34524 24915 34527
rect 25130 34524 25136 34536
rect 24903 34496 25136 34524
rect 24903 34493 24915 34496
rect 24857 34487 24915 34493
rect 25130 34484 25136 34496
rect 25188 34484 25194 34536
rect 26804 34524 26832 34564
rect 26878 34552 26884 34604
rect 26936 34592 26942 34604
rect 26973 34595 27031 34601
rect 26973 34592 26985 34595
rect 26936 34564 26985 34592
rect 26936 34552 26942 34564
rect 26973 34561 26985 34564
rect 27019 34561 27031 34595
rect 26973 34555 27031 34561
rect 28721 34595 28779 34601
rect 28721 34561 28733 34595
rect 28767 34592 28779 34595
rect 28902 34592 28908 34604
rect 28767 34564 28908 34592
rect 28767 34561 28779 34564
rect 28721 34555 28779 34561
rect 28736 34524 28764 34555
rect 28902 34552 28908 34564
rect 28960 34552 28966 34604
rect 30024 34601 30052 34632
rect 30653 34629 30665 34632
rect 30699 34660 30711 34663
rect 33502 34660 33508 34672
rect 30699 34632 33508 34660
rect 30699 34629 30711 34632
rect 30653 34623 30711 34629
rect 33502 34620 33508 34632
rect 33560 34620 33566 34672
rect 30009 34595 30067 34601
rect 30009 34561 30021 34595
rect 30055 34561 30067 34595
rect 30009 34555 30067 34561
rect 30193 34595 30251 34601
rect 30193 34561 30205 34595
rect 30239 34592 30251 34595
rect 30282 34592 30288 34604
rect 30239 34564 30288 34592
rect 30239 34561 30251 34564
rect 30193 34555 30251 34561
rect 30282 34552 30288 34564
rect 30340 34592 30346 34604
rect 30837 34595 30895 34601
rect 30837 34592 30849 34595
rect 30340 34564 30849 34592
rect 30340 34552 30346 34564
rect 30837 34561 30849 34564
rect 30883 34561 30895 34595
rect 48130 34592 48136 34604
rect 48091 34564 48136 34592
rect 30837 34555 30895 34561
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 26804 34496 28764 34524
rect 27065 34459 27123 34465
rect 27065 34425 27077 34459
rect 27111 34456 27123 34459
rect 27246 34456 27252 34468
rect 27111 34428 27252 34456
rect 27111 34425 27123 34428
rect 27065 34419 27123 34425
rect 27246 34416 27252 34428
rect 27304 34456 27310 34468
rect 29178 34456 29184 34468
rect 27304 34428 29184 34456
rect 27304 34416 27310 34428
rect 29178 34416 29184 34428
rect 29236 34416 29242 34468
rect 20806 34348 20812 34400
rect 20864 34388 20870 34400
rect 20901 34391 20959 34397
rect 20901 34388 20913 34391
rect 20864 34360 20913 34388
rect 20864 34348 20870 34360
rect 20901 34357 20913 34360
rect 20947 34357 20959 34391
rect 20901 34351 20959 34357
rect 22084 34391 22142 34397
rect 22084 34357 22096 34391
rect 22130 34388 22142 34391
rect 22646 34388 22652 34400
rect 22130 34360 22652 34388
rect 22130 34357 22142 34360
rect 22084 34351 22142 34357
rect 22646 34348 22652 34360
rect 22704 34348 22710 34400
rect 22830 34348 22836 34400
rect 22888 34388 22894 34400
rect 23569 34391 23627 34397
rect 23569 34388 23581 34391
rect 22888 34360 23581 34388
rect 22888 34348 22894 34360
rect 23569 34357 23581 34360
rect 23615 34388 23627 34391
rect 24946 34388 24952 34400
rect 23615 34360 24952 34388
rect 23615 34357 23627 34360
rect 23569 34351 23627 34357
rect 24946 34348 24952 34360
rect 25004 34348 25010 34400
rect 25958 34348 25964 34400
rect 26016 34388 26022 34400
rect 30098 34388 30104 34400
rect 26016 34360 30104 34388
rect 26016 34348 26022 34360
rect 30098 34348 30104 34360
rect 30156 34348 30162 34400
rect 30374 34348 30380 34400
rect 30432 34388 30438 34400
rect 31021 34391 31079 34397
rect 31021 34388 31033 34391
rect 30432 34360 31033 34388
rect 30432 34348 30438 34360
rect 31021 34357 31033 34360
rect 31067 34357 31079 34391
rect 31021 34351 31079 34357
rect 47854 34348 47860 34400
rect 47912 34388 47918 34400
rect 47949 34391 48007 34397
rect 47949 34388 47961 34391
rect 47912 34360 47961 34388
rect 47912 34348 47918 34360
rect 47949 34357 47961 34360
rect 47995 34357 48007 34391
rect 47949 34351 48007 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 22646 34184 22652 34196
rect 22607 34156 22652 34184
rect 22646 34144 22652 34156
rect 22704 34144 22710 34196
rect 23198 34184 23204 34196
rect 23159 34156 23204 34184
rect 23198 34144 23204 34156
rect 23256 34144 23262 34196
rect 26510 34144 26516 34196
rect 26568 34184 26574 34196
rect 26605 34187 26663 34193
rect 26605 34184 26617 34187
rect 26568 34156 26617 34184
rect 26568 34144 26574 34156
rect 26605 34153 26617 34156
rect 26651 34153 26663 34187
rect 26605 34147 26663 34153
rect 29733 34187 29791 34193
rect 29733 34153 29745 34187
rect 29779 34184 29791 34187
rect 29822 34184 29828 34196
rect 29779 34156 29828 34184
rect 29779 34153 29791 34156
rect 29733 34147 29791 34153
rect 29822 34144 29828 34156
rect 29880 34144 29886 34196
rect 48041 34187 48099 34193
rect 48041 34184 48053 34187
rect 29932 34156 48053 34184
rect 20806 34076 20812 34128
rect 20864 34116 20870 34128
rect 22002 34116 22008 34128
rect 20864 34088 22008 34116
rect 20864 34076 20870 34088
rect 22002 34076 22008 34088
rect 22060 34116 22066 34128
rect 22060 34088 23152 34116
rect 22060 34076 22066 34088
rect 16942 34008 16948 34060
rect 17000 34048 17006 34060
rect 22281 34051 22339 34057
rect 22281 34048 22293 34051
rect 17000 34020 22293 34048
rect 17000 34008 17006 34020
rect 22281 34017 22293 34020
rect 22327 34017 22339 34051
rect 22281 34011 22339 34017
rect 20806 33980 20812 33992
rect 20767 33952 20812 33980
rect 20806 33940 20812 33952
rect 20864 33940 20870 33992
rect 21910 33980 21916 33992
rect 21871 33952 21916 33980
rect 21910 33940 21916 33952
rect 21968 33940 21974 33992
rect 22192 33983 22250 33989
rect 22085 33977 22143 33983
rect 22085 33943 22097 33977
rect 22131 33943 22143 33977
rect 22192 33949 22204 33983
rect 22238 33949 22250 33983
rect 22192 33943 22250 33949
rect 22465 33983 22523 33989
rect 22465 33949 22477 33983
rect 22511 33980 22523 33983
rect 22738 33980 22744 33992
rect 22511 33952 22744 33980
rect 22511 33949 22523 33952
rect 22465 33943 22523 33949
rect 22085 33937 22143 33943
rect 20898 33844 20904 33856
rect 20859 33816 20904 33844
rect 20898 33804 20904 33816
rect 20956 33804 20962 33856
rect 22099 33844 22127 33937
rect 22204 33912 22232 33943
rect 22738 33940 22744 33952
rect 22796 33940 22802 33992
rect 23124 33989 23152 34088
rect 29546 34076 29552 34128
rect 29604 34116 29610 34128
rect 29932 34116 29960 34156
rect 48041 34153 48053 34156
rect 48087 34153 48099 34187
rect 48041 34147 48099 34153
rect 29604 34088 29960 34116
rect 29604 34076 29610 34088
rect 24210 34008 24216 34060
rect 24268 34048 24274 34060
rect 24397 34051 24455 34057
rect 24397 34048 24409 34051
rect 24268 34020 24409 34048
rect 24268 34008 24274 34020
rect 24397 34017 24409 34020
rect 24443 34048 24455 34051
rect 24670 34048 24676 34060
rect 24443 34020 24676 34048
rect 24443 34017 24455 34020
rect 24397 34011 24455 34017
rect 24670 34008 24676 34020
rect 24728 34008 24734 34060
rect 26510 34008 26516 34060
rect 26568 34048 26574 34060
rect 26789 34051 26847 34057
rect 26568 34020 26740 34048
rect 26568 34008 26574 34020
rect 23109 33983 23167 33989
rect 23109 33949 23121 33983
rect 23155 33949 23167 33983
rect 23109 33943 23167 33949
rect 26142 33940 26148 33992
rect 26200 33980 26206 33992
rect 26605 33983 26663 33989
rect 26605 33980 26617 33983
rect 26200 33952 26617 33980
rect 26200 33940 26206 33952
rect 26605 33949 26617 33952
rect 26651 33949 26663 33983
rect 26712 33980 26740 34020
rect 26789 34017 26801 34051
rect 26835 34048 26847 34051
rect 27246 34048 27252 34060
rect 26835 34020 27252 34048
rect 26835 34017 26847 34020
rect 26789 34011 26847 34017
rect 27246 34008 27252 34020
rect 27304 34008 27310 34060
rect 28721 34051 28779 34057
rect 28721 34017 28733 34051
rect 28767 34048 28779 34051
rect 28994 34048 29000 34060
rect 28767 34020 29000 34048
rect 28767 34017 28779 34020
rect 28721 34011 28779 34017
rect 28994 34008 29000 34020
rect 29052 34008 29058 34060
rect 30285 34051 30343 34057
rect 30285 34017 30297 34051
rect 30331 34048 30343 34051
rect 30374 34048 30380 34060
rect 30331 34020 30380 34048
rect 30331 34017 30343 34020
rect 30285 34011 30343 34017
rect 30374 34008 30380 34020
rect 30432 34008 30438 34060
rect 31110 34048 31116 34060
rect 31071 34020 31116 34048
rect 31110 34008 31116 34020
rect 31168 34008 31174 34060
rect 26881 33983 26939 33989
rect 26881 33980 26893 33983
rect 26712 33952 26893 33980
rect 26605 33943 26663 33949
rect 26881 33949 26893 33952
rect 26927 33949 26939 33983
rect 28442 33980 28448 33992
rect 28403 33952 28448 33980
rect 26881 33943 26939 33949
rect 28442 33940 28448 33952
rect 28500 33940 28506 33992
rect 28537 33983 28595 33989
rect 28537 33949 28549 33983
rect 28583 33980 28595 33983
rect 29638 33980 29644 33992
rect 28583 33952 29644 33980
rect 28583 33949 28595 33952
rect 28537 33943 28595 33949
rect 29638 33940 29644 33952
rect 29696 33940 29702 33992
rect 29917 33983 29975 33989
rect 29917 33980 29929 33983
rect 29748 33952 29929 33980
rect 22830 33912 22836 33924
rect 22204 33884 22836 33912
rect 22830 33872 22836 33884
rect 22888 33872 22894 33924
rect 24670 33912 24676 33924
rect 24631 33884 24676 33912
rect 24670 33872 24676 33884
rect 24728 33872 24734 33924
rect 25130 33872 25136 33924
rect 25188 33872 25194 33924
rect 29362 33912 29368 33924
rect 25976 33884 29368 33912
rect 22278 33844 22284 33856
rect 22099 33816 22284 33844
rect 22278 33804 22284 33816
rect 22336 33844 22342 33856
rect 25976 33844 26004 33884
rect 29362 33872 29368 33884
rect 29420 33872 29426 33924
rect 26142 33844 26148 33856
rect 22336 33816 26004 33844
rect 26103 33816 26148 33844
rect 22336 33804 22342 33816
rect 26142 33804 26148 33816
rect 26200 33804 26206 33856
rect 27062 33844 27068 33856
rect 27023 33816 27068 33844
rect 27062 33804 27068 33816
rect 27120 33804 27126 33856
rect 27154 33804 27160 33856
rect 27212 33844 27218 33856
rect 28721 33847 28779 33853
rect 28721 33844 28733 33847
rect 27212 33816 28733 33844
rect 27212 33804 27218 33816
rect 28721 33813 28733 33816
rect 28767 33813 28779 33847
rect 29748 33844 29776 33952
rect 29917 33949 29929 33952
rect 29963 33949 29975 33983
rect 29917 33943 29975 33949
rect 30009 33983 30067 33989
rect 30009 33949 30021 33983
rect 30055 33949 30067 33983
rect 33318 33980 33324 33992
rect 33279 33952 33324 33980
rect 30009 33943 30067 33949
rect 29822 33872 29828 33924
rect 29880 33912 29886 33924
rect 30024 33912 30052 33943
rect 33318 33940 33324 33952
rect 33376 33940 33382 33992
rect 33502 33980 33508 33992
rect 33463 33952 33508 33980
rect 33502 33940 33508 33952
rect 33560 33940 33566 33992
rect 47857 33983 47915 33989
rect 47857 33949 47869 33983
rect 47903 33980 47915 33983
rect 47946 33980 47952 33992
rect 47903 33952 47952 33980
rect 47903 33949 47915 33952
rect 47857 33943 47915 33949
rect 47946 33940 47952 33952
rect 48004 33940 48010 33992
rect 29880 33884 30052 33912
rect 29880 33872 29886 33884
rect 30098 33872 30104 33924
rect 30156 33912 30162 33924
rect 30377 33915 30435 33921
rect 30377 33912 30389 33915
rect 30156 33884 30389 33912
rect 30156 33872 30162 33884
rect 30377 33881 30389 33884
rect 30423 33881 30435 33915
rect 31386 33912 31392 33924
rect 31347 33884 31392 33912
rect 30377 33875 30435 33881
rect 31386 33872 31392 33884
rect 31444 33872 31450 33924
rect 31846 33872 31852 33924
rect 31904 33872 31910 33924
rect 30282 33844 30288 33856
rect 29748 33816 30288 33844
rect 28721 33807 28779 33813
rect 30282 33804 30288 33816
rect 30340 33804 30346 33856
rect 31294 33804 31300 33856
rect 31352 33844 31358 33856
rect 32398 33844 32404 33856
rect 31352 33816 32404 33844
rect 31352 33804 31358 33816
rect 32398 33804 32404 33816
rect 32456 33844 32462 33856
rect 32861 33847 32919 33853
rect 32861 33844 32873 33847
rect 32456 33816 32873 33844
rect 32456 33804 32462 33816
rect 32861 33813 32873 33816
rect 32907 33813 32919 33847
rect 33502 33844 33508 33856
rect 33463 33816 33508 33844
rect 32861 33807 32919 33813
rect 33502 33804 33508 33816
rect 33560 33804 33566 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 23474 33640 23480 33652
rect 19536 33612 23480 33640
rect 16022 33572 16028 33584
rect 15983 33544 16028 33572
rect 16022 33532 16028 33544
rect 16080 33532 16086 33584
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33504 1731 33507
rect 2682 33504 2688 33516
rect 1719 33476 2688 33504
rect 1719 33473 1731 33476
rect 1673 33467 1731 33473
rect 2682 33464 2688 33476
rect 2740 33464 2746 33516
rect 19536 33513 19564 33612
rect 23474 33600 23480 33612
rect 23532 33600 23538 33652
rect 24670 33600 24676 33652
rect 24728 33640 24734 33652
rect 25041 33643 25099 33649
rect 25041 33640 25053 33643
rect 24728 33612 25053 33640
rect 24728 33600 24734 33612
rect 25041 33609 25053 33612
rect 25087 33609 25099 33643
rect 27154 33640 27160 33652
rect 25041 33603 25099 33609
rect 25700 33612 27160 33640
rect 19521 33507 19579 33513
rect 19521 33473 19533 33507
rect 19567 33473 19579 33507
rect 19521 33467 19579 33473
rect 20898 33464 20904 33516
rect 20956 33464 20962 33516
rect 24857 33507 24915 33513
rect 24857 33473 24869 33507
rect 24903 33504 24915 33507
rect 25700 33504 25728 33612
rect 27154 33600 27160 33612
rect 27212 33600 27218 33652
rect 27338 33640 27344 33652
rect 27299 33612 27344 33640
rect 27338 33600 27344 33612
rect 27396 33600 27402 33652
rect 27798 33600 27804 33652
rect 27856 33640 27862 33652
rect 28537 33643 28595 33649
rect 28537 33640 28549 33643
rect 27856 33612 28549 33640
rect 27856 33600 27862 33612
rect 28537 33609 28549 33612
rect 28583 33609 28595 33643
rect 28537 33603 28595 33609
rect 28994 33600 29000 33652
rect 29052 33640 29058 33652
rect 29822 33640 29828 33652
rect 29052 33612 29828 33640
rect 29052 33600 29058 33612
rect 29822 33600 29828 33612
rect 29880 33600 29886 33652
rect 31386 33600 31392 33652
rect 31444 33640 31450 33652
rect 31573 33643 31631 33649
rect 31573 33640 31585 33643
rect 31444 33612 31585 33640
rect 31444 33600 31450 33612
rect 31573 33609 31585 33612
rect 31619 33609 31631 33643
rect 33134 33640 33140 33652
rect 31573 33603 31631 33609
rect 31772 33612 33140 33640
rect 25777 33575 25835 33581
rect 25777 33541 25789 33575
rect 25823 33572 25835 33575
rect 27062 33572 27068 33584
rect 25823 33544 27068 33572
rect 25823 33541 25835 33544
rect 25777 33535 25835 33541
rect 27062 33532 27068 33544
rect 27120 33532 27126 33584
rect 29365 33575 29423 33581
rect 29365 33572 29377 33575
rect 27816 33544 29377 33572
rect 24903 33476 25728 33504
rect 24903 33473 24915 33476
rect 24857 33467 24915 33473
rect 25866 33464 25872 33516
rect 25924 33504 25930 33516
rect 25961 33507 26019 33513
rect 25961 33504 25973 33507
rect 25924 33476 25973 33504
rect 25924 33464 25930 33476
rect 25961 33473 25973 33476
rect 26007 33473 26019 33507
rect 25961 33467 26019 33473
rect 26878 33464 26884 33516
rect 26936 33504 26942 33516
rect 26973 33507 27031 33513
rect 26973 33504 26985 33507
rect 26936 33476 26985 33504
rect 26936 33464 26942 33476
rect 26973 33473 26985 33476
rect 27019 33473 27031 33507
rect 26973 33467 27031 33473
rect 27157 33507 27215 33513
rect 27157 33473 27169 33507
rect 27203 33504 27215 33507
rect 27246 33504 27252 33516
rect 27203 33476 27252 33504
rect 27203 33473 27215 33476
rect 27157 33467 27215 33473
rect 27246 33464 27252 33476
rect 27304 33464 27310 33516
rect 27816 33513 27844 33544
rect 29365 33541 29377 33544
rect 29411 33541 29423 33575
rect 29365 33535 29423 33541
rect 29454 33532 29460 33584
rect 29512 33572 29518 33584
rect 29512 33544 31064 33572
rect 29512 33532 29518 33544
rect 27801 33507 27859 33513
rect 27801 33473 27813 33507
rect 27847 33473 27859 33507
rect 27985 33507 28043 33513
rect 27985 33504 27997 33507
rect 27801 33467 27859 33473
rect 27908 33476 27997 33504
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 13630 33396 13636 33448
rect 13688 33436 13694 33448
rect 14185 33439 14243 33445
rect 14185 33436 14197 33439
rect 13688 33408 14197 33436
rect 13688 33396 13694 33408
rect 14185 33405 14197 33408
rect 14231 33405 14243 33439
rect 14366 33436 14372 33448
rect 14327 33408 14372 33436
rect 14185 33399 14243 33405
rect 14366 33396 14372 33408
rect 14424 33396 14430 33448
rect 19797 33439 19855 33445
rect 19797 33405 19809 33439
rect 19843 33436 19855 33439
rect 22002 33436 22008 33448
rect 19843 33408 22008 33436
rect 19843 33405 19855 33408
rect 19797 33399 19855 33405
rect 22002 33396 22008 33408
rect 22060 33396 22066 33448
rect 24302 33396 24308 33448
rect 24360 33436 24366 33448
rect 24397 33439 24455 33445
rect 24397 33436 24409 33439
rect 24360 33408 24409 33436
rect 24360 33396 24366 33408
rect 24397 33405 24409 33408
rect 24443 33405 24455 33439
rect 24397 33399 24455 33405
rect 24765 33439 24823 33445
rect 24765 33405 24777 33439
rect 24811 33436 24823 33439
rect 26142 33436 26148 33448
rect 24811 33408 26148 33436
rect 24811 33405 24823 33408
rect 24765 33399 24823 33405
rect 26142 33396 26148 33408
rect 26200 33396 26206 33448
rect 22370 33328 22376 33380
rect 22428 33368 22434 33380
rect 27908 33368 27936 33476
rect 27985 33473 27997 33476
rect 28031 33504 28043 33507
rect 28353 33507 28411 33513
rect 28031 33476 28304 33504
rect 28031 33473 28043 33476
rect 27985 33467 28043 33473
rect 28074 33436 28080 33448
rect 28035 33408 28080 33436
rect 28074 33396 28080 33408
rect 28132 33396 28138 33448
rect 28169 33439 28227 33445
rect 28169 33405 28181 33439
rect 28215 33405 28227 33439
rect 28276 33436 28304 33476
rect 28353 33473 28365 33507
rect 28399 33504 28411 33507
rect 28442 33504 28448 33516
rect 28399 33476 28448 33504
rect 28399 33473 28411 33476
rect 28353 33467 28411 33473
rect 28442 33464 28448 33476
rect 28500 33464 28506 33516
rect 28994 33464 29000 33516
rect 29052 33504 29058 33516
rect 29178 33504 29184 33516
rect 29052 33476 29097 33504
rect 29139 33476 29184 33504
rect 29052 33464 29058 33476
rect 29178 33464 29184 33476
rect 29236 33464 29242 33516
rect 30009 33507 30067 33513
rect 30009 33473 30021 33507
rect 30055 33504 30067 33507
rect 30190 33504 30196 33516
rect 30055 33476 30196 33504
rect 30055 33473 30067 33476
rect 30009 33467 30067 33473
rect 30190 33464 30196 33476
rect 30248 33464 30254 33516
rect 30834 33504 30840 33516
rect 30795 33476 30840 33504
rect 30834 33464 30840 33476
rect 30892 33464 30898 33516
rect 31036 33513 31064 33544
rect 31021 33507 31079 33513
rect 31021 33473 31033 33507
rect 31067 33473 31079 33507
rect 31021 33467 31079 33473
rect 31113 33507 31171 33513
rect 31113 33473 31125 33507
rect 31159 33504 31171 33507
rect 31294 33504 31300 33516
rect 31159 33476 31300 33504
rect 31159 33473 31171 33476
rect 31113 33467 31171 33473
rect 31294 33464 31300 33476
rect 31352 33464 31358 33516
rect 31389 33507 31447 33513
rect 31389 33473 31401 33507
rect 31435 33504 31447 33507
rect 31772 33504 31800 33612
rect 33134 33600 33140 33612
rect 33192 33600 33198 33652
rect 35897 33643 35955 33649
rect 35897 33640 35909 33643
rect 33244 33612 35909 33640
rect 32950 33532 32956 33584
rect 33008 33572 33014 33584
rect 33244 33572 33272 33612
rect 35897 33609 35909 33612
rect 35943 33609 35955 33643
rect 35897 33603 35955 33609
rect 33008 33544 33272 33572
rect 33008 33532 33014 33544
rect 31435 33476 31800 33504
rect 31435 33473 31447 33476
rect 31389 33467 31447 33473
rect 28534 33436 28540 33448
rect 28276 33408 28540 33436
rect 28169 33399 28227 33405
rect 22428 33340 27936 33368
rect 22428 33328 22434 33340
rect 28184 33312 28212 33399
rect 28534 33396 28540 33408
rect 28592 33396 28598 33448
rect 31205 33439 31263 33445
rect 31205 33405 31217 33439
rect 31251 33436 31263 33439
rect 31662 33436 31668 33448
rect 31251 33408 31668 33436
rect 31251 33405 31263 33408
rect 31205 33399 31263 33405
rect 31662 33396 31668 33408
rect 31720 33396 31726 33448
rect 31772 33368 31800 33476
rect 32125 33507 32183 33513
rect 32125 33473 32137 33507
rect 32171 33504 32183 33507
rect 32398 33504 32404 33516
rect 32171 33476 32260 33504
rect 32359 33476 32404 33504
rect 32171 33473 32183 33476
rect 32125 33467 32183 33473
rect 29288 33340 31800 33368
rect 32232 33368 32260 33476
rect 32398 33464 32404 33476
rect 32456 33464 32462 33516
rect 32766 33464 32772 33516
rect 32824 33504 32830 33516
rect 33244 33513 33272 33544
rect 35434 33532 35440 33584
rect 35492 33532 35498 33584
rect 46106 33532 46112 33584
rect 46164 33572 46170 33584
rect 46164 33544 47624 33572
rect 46164 33532 46170 33544
rect 47596 33513 47624 33544
rect 33045 33507 33103 33513
rect 33045 33504 33057 33507
rect 32824 33476 33057 33504
rect 32824 33464 32830 33476
rect 33045 33473 33057 33476
rect 33091 33473 33103 33507
rect 33045 33467 33103 33473
rect 33229 33507 33287 33513
rect 33229 33473 33241 33507
rect 33275 33473 33287 33507
rect 33229 33467 33287 33473
rect 47029 33507 47087 33513
rect 47029 33473 47041 33507
rect 47075 33473 47087 33507
rect 47029 33467 47087 33473
rect 47581 33507 47639 33513
rect 47581 33473 47593 33507
rect 47627 33473 47639 33507
rect 47581 33467 47639 33473
rect 32309 33439 32367 33445
rect 32309 33405 32321 33439
rect 32355 33436 32367 33439
rect 32950 33436 32956 33448
rect 32355 33408 32956 33436
rect 32355 33405 32367 33408
rect 32309 33399 32367 33405
rect 32950 33396 32956 33408
rect 33008 33396 33014 33448
rect 33686 33396 33692 33448
rect 33744 33436 33750 33448
rect 34149 33439 34207 33445
rect 34149 33436 34161 33439
rect 33744 33408 34161 33436
rect 33744 33396 33750 33408
rect 34149 33405 34161 33408
rect 34195 33405 34207 33439
rect 34422 33436 34428 33448
rect 34383 33408 34428 33436
rect 34149 33399 34207 33405
rect 34422 33396 34428 33408
rect 34480 33396 34486 33448
rect 47044 33436 47072 33467
rect 48041 33439 48099 33445
rect 48041 33436 48053 33439
rect 47044 33408 48053 33436
rect 48041 33405 48053 33408
rect 48087 33405 48099 33439
rect 48041 33399 48099 33405
rect 33410 33368 33416 33380
rect 32232 33340 32720 33368
rect 33371 33340 33416 33368
rect 2774 33300 2780 33312
rect 2735 33272 2780 33300
rect 2774 33260 2780 33272
rect 2832 33260 2838 33312
rect 3145 33303 3203 33309
rect 3145 33269 3157 33303
rect 3191 33300 3203 33303
rect 3970 33300 3976 33312
rect 3191 33272 3976 33300
rect 3191 33269 3203 33272
rect 3145 33263 3203 33269
rect 3970 33260 3976 33272
rect 4028 33260 4034 33312
rect 21269 33303 21327 33309
rect 21269 33269 21281 33303
rect 21315 33300 21327 33303
rect 21726 33300 21732 33312
rect 21315 33272 21732 33300
rect 21315 33269 21327 33272
rect 21269 33263 21327 33269
rect 21726 33260 21732 33272
rect 21784 33260 21790 33312
rect 21910 33260 21916 33312
rect 21968 33300 21974 33312
rect 23382 33300 23388 33312
rect 21968 33272 23388 33300
rect 21968 33260 21974 33272
rect 23382 33260 23388 33272
rect 23440 33260 23446 33312
rect 25130 33260 25136 33312
rect 25188 33300 25194 33312
rect 26145 33303 26203 33309
rect 26145 33300 26157 33303
rect 25188 33272 26157 33300
rect 25188 33260 25194 33272
rect 26145 33269 26157 33272
rect 26191 33269 26203 33303
rect 26970 33300 26976 33312
rect 26931 33272 26976 33300
rect 26145 33263 26203 33269
rect 26970 33260 26976 33272
rect 27028 33260 27034 33312
rect 28166 33260 28172 33312
rect 28224 33260 28230 33312
rect 28442 33260 28448 33312
rect 28500 33300 28506 33312
rect 29288 33300 29316 33340
rect 32692 33312 32720 33340
rect 33410 33328 33416 33340
rect 33468 33328 33474 33380
rect 28500 33272 29316 33300
rect 28500 33260 28506 33272
rect 30282 33260 30288 33312
rect 30340 33300 30346 33312
rect 32125 33303 32183 33309
rect 32125 33300 32137 33303
rect 30340 33272 32137 33300
rect 30340 33260 30346 33272
rect 32125 33269 32137 33272
rect 32171 33269 32183 33303
rect 32582 33300 32588 33312
rect 32543 33272 32588 33300
rect 32125 33263 32183 33269
rect 32582 33260 32588 33272
rect 32640 33260 32646 33312
rect 32674 33260 32680 33312
rect 32732 33300 32738 33312
rect 33045 33303 33103 33309
rect 33045 33300 33057 33303
rect 32732 33272 33057 33300
rect 32732 33260 32738 33272
rect 33045 33269 33057 33272
rect 33091 33269 33103 33303
rect 33045 33263 33103 33269
rect 46845 33303 46903 33309
rect 46845 33269 46857 33303
rect 46891 33300 46903 33303
rect 47302 33300 47308 33312
rect 46891 33272 47308 33300
rect 46891 33269 46903 33272
rect 46845 33263 46903 33269
rect 47302 33260 47308 33272
rect 47360 33260 47366 33312
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 11698 33056 11704 33108
rect 11756 33056 11762 33108
rect 22002 33056 22008 33108
rect 22060 33096 22066 33108
rect 22925 33099 22983 33105
rect 22925 33096 22937 33099
rect 22060 33068 22937 33096
rect 22060 33056 22066 33068
rect 22925 33065 22937 33068
rect 22971 33065 22983 33099
rect 25130 33096 25136 33108
rect 25091 33068 25136 33096
rect 22925 33059 22983 33065
rect 25130 33056 25136 33068
rect 25188 33056 25194 33108
rect 26050 33096 26056 33108
rect 26011 33068 26056 33096
rect 26050 33056 26056 33068
rect 26108 33056 26114 33108
rect 27985 33099 28043 33105
rect 27985 33065 27997 33099
rect 28031 33096 28043 33099
rect 29086 33096 29092 33108
rect 28031 33068 29092 33096
rect 28031 33065 28043 33068
rect 27985 33059 28043 33065
rect 29086 33056 29092 33068
rect 29144 33056 29150 33108
rect 30561 33099 30619 33105
rect 30561 33065 30573 33099
rect 30607 33096 30619 33099
rect 30834 33096 30840 33108
rect 30607 33068 30840 33096
rect 30607 33065 30619 33068
rect 30561 33059 30619 33065
rect 30834 33056 30840 33068
rect 30892 33056 30898 33108
rect 32398 33056 32404 33108
rect 32456 33096 32462 33108
rect 32766 33096 32772 33108
rect 32456 33068 32772 33096
rect 32456 33056 32462 33068
rect 32766 33056 32772 33068
rect 32824 33056 32830 33108
rect 32861 33099 32919 33105
rect 32861 33065 32873 33099
rect 32907 33096 32919 33099
rect 33318 33096 33324 33108
rect 32907 33068 33324 33096
rect 32907 33065 32919 33068
rect 32861 33059 32919 33065
rect 33318 33056 33324 33068
rect 33376 33056 33382 33108
rect 34149 33099 34207 33105
rect 34149 33065 34161 33099
rect 34195 33096 34207 33099
rect 34422 33096 34428 33108
rect 34195 33068 34428 33096
rect 34195 33065 34207 33068
rect 34149 33059 34207 33065
rect 34422 33056 34428 33068
rect 34480 33056 34486 33108
rect 35345 33099 35403 33105
rect 35345 33065 35357 33099
rect 35391 33096 35403 33099
rect 35434 33096 35440 33108
rect 35391 33068 35440 33096
rect 35391 33065 35403 33068
rect 35345 33059 35403 33065
rect 35434 33056 35440 33068
rect 35492 33056 35498 33108
rect 1486 33028 1492 33040
rect 1412 33000 1492 33028
rect 1412 32969 1440 33000
rect 1486 32988 1492 33000
rect 1544 32988 1550 33040
rect 11716 33028 11744 33056
rect 23566 33028 23572 33040
rect 11716 33000 23572 33028
rect 23566 32988 23572 33000
rect 23624 32988 23630 33040
rect 27341 33031 27399 33037
rect 27341 32997 27353 33031
rect 27387 33028 27399 33031
rect 28074 33028 28080 33040
rect 27387 33000 28080 33028
rect 27387 32997 27399 33000
rect 27341 32991 27399 32997
rect 28074 32988 28080 33000
rect 28132 32988 28138 33040
rect 28534 32988 28540 33040
rect 28592 33028 28598 33040
rect 29822 33028 29828 33040
rect 28592 33000 29828 33028
rect 28592 32988 28598 33000
rect 29822 32988 29828 33000
rect 29880 32988 29886 33040
rect 33134 32988 33140 33040
rect 33192 33028 33198 33040
rect 33192 33000 34008 33028
rect 33192 32988 33198 33000
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32929 1455 32963
rect 11698 32960 11704 32972
rect 11659 32932 11704 32960
rect 1397 32923 1455 32929
rect 11698 32920 11704 32932
rect 11756 32920 11762 32972
rect 14185 32963 14243 32969
rect 14185 32960 14197 32963
rect 13280 32932 14197 32960
rect 13280 32904 13308 32932
rect 14185 32929 14197 32932
rect 14231 32929 14243 32963
rect 14185 32923 14243 32929
rect 16025 32963 16083 32969
rect 16025 32929 16037 32963
rect 16071 32960 16083 32963
rect 16114 32960 16120 32972
rect 16071 32932 16120 32960
rect 16071 32929 16083 32932
rect 16025 32923 16083 32929
rect 16114 32920 16120 32932
rect 16172 32920 16178 32972
rect 25866 32960 25872 32972
rect 25827 32932 25872 32960
rect 25866 32920 25872 32932
rect 25924 32920 25930 32972
rect 26234 32920 26240 32972
rect 26292 32960 26298 32972
rect 26878 32960 26884 32972
rect 26292 32932 26884 32960
rect 26292 32920 26298 32932
rect 26878 32920 26884 32932
rect 26936 32920 26942 32972
rect 27798 32920 27804 32972
rect 27856 32960 27862 32972
rect 30098 32960 30104 32972
rect 27856 32932 30104 32960
rect 27856 32920 27862 32932
rect 30098 32920 30104 32932
rect 30156 32920 30162 32972
rect 31294 32960 31300 32972
rect 30852 32932 31300 32960
rect 3970 32892 3976 32904
rect 3931 32864 3976 32892
rect 3970 32852 3976 32864
rect 4028 32852 4034 32904
rect 11609 32895 11667 32901
rect 11609 32861 11621 32895
rect 11655 32892 11667 32895
rect 13262 32892 13268 32904
rect 11655 32864 13268 32892
rect 11655 32861 11667 32864
rect 11609 32855 11667 32861
rect 13262 32852 13268 32864
rect 13320 32852 13326 32904
rect 13357 32895 13415 32901
rect 13357 32861 13369 32895
rect 13403 32892 13415 32895
rect 13538 32892 13544 32904
rect 13403 32864 13544 32892
rect 13403 32861 13415 32864
rect 13357 32855 13415 32861
rect 1581 32827 1639 32833
rect 1581 32793 1593 32827
rect 1627 32793 1639 32827
rect 3234 32824 3240 32836
rect 3195 32796 3240 32824
rect 1581 32787 1639 32793
rect 1596 32756 1624 32787
rect 3234 32784 3240 32796
rect 3292 32784 3298 32836
rect 9674 32784 9680 32836
rect 9732 32824 9738 32836
rect 13372 32824 13400 32855
rect 13538 32852 13544 32864
rect 13596 32852 13602 32904
rect 20346 32852 20352 32904
rect 20404 32892 20410 32904
rect 21361 32895 21419 32901
rect 21361 32892 21373 32895
rect 20404 32864 21373 32892
rect 20404 32852 20410 32864
rect 21361 32861 21373 32864
rect 21407 32861 21419 32895
rect 21361 32855 21419 32861
rect 21729 32895 21787 32901
rect 21729 32861 21741 32895
rect 21775 32892 21787 32895
rect 22189 32895 22247 32901
rect 22189 32892 22201 32895
rect 21775 32864 22201 32892
rect 21775 32861 21787 32864
rect 21729 32855 21787 32861
rect 22189 32861 22201 32864
rect 22235 32861 22247 32895
rect 22370 32892 22376 32904
rect 22331 32864 22376 32892
rect 22189 32855 22247 32861
rect 22370 32852 22376 32864
rect 22428 32852 22434 32904
rect 22462 32852 22468 32904
rect 22520 32892 22526 32904
rect 22646 32901 22652 32904
rect 22603 32895 22652 32901
rect 22520 32864 22565 32892
rect 22520 32852 22526 32864
rect 22603 32861 22615 32895
rect 22649 32861 22652 32895
rect 22603 32855 22652 32861
rect 22646 32852 22652 32855
rect 22704 32852 22710 32904
rect 22741 32895 22799 32901
rect 22741 32861 22753 32895
rect 22787 32861 22799 32895
rect 24946 32892 24952 32904
rect 24907 32864 24952 32892
rect 22741 32855 22799 32861
rect 9732 32796 13400 32824
rect 13449 32827 13507 32833
rect 9732 32784 9738 32796
rect 13449 32793 13461 32827
rect 13495 32824 13507 32827
rect 14369 32827 14427 32833
rect 14369 32824 14381 32827
rect 13495 32796 14381 32824
rect 13495 32793 13507 32796
rect 13449 32787 13507 32793
rect 14369 32793 14381 32796
rect 14415 32793 14427 32827
rect 14369 32787 14427 32793
rect 21545 32827 21603 32833
rect 21545 32793 21557 32827
rect 21591 32793 21603 32827
rect 21545 32787 21603 32793
rect 3789 32759 3847 32765
rect 3789 32756 3801 32759
rect 1596 32728 3801 32756
rect 3789 32725 3801 32728
rect 3835 32725 3847 32759
rect 3789 32719 3847 32725
rect 11790 32716 11796 32768
rect 11848 32756 11854 32768
rect 11977 32759 12035 32765
rect 11977 32756 11989 32759
rect 11848 32728 11989 32756
rect 11848 32716 11854 32728
rect 11977 32725 11989 32728
rect 12023 32725 12035 32759
rect 21560 32756 21588 32787
rect 22002 32784 22008 32836
rect 22060 32824 22066 32836
rect 22756 32824 22784 32855
rect 24946 32852 24952 32864
rect 25004 32852 25010 32904
rect 25222 32892 25228 32904
rect 25183 32864 25228 32892
rect 25222 32852 25228 32864
rect 25280 32852 25286 32904
rect 26053 32895 26111 32901
rect 26053 32861 26065 32895
rect 26099 32892 26111 32895
rect 26142 32892 26148 32904
rect 26099 32864 26148 32892
rect 26099 32861 26111 32864
rect 26053 32855 26111 32861
rect 26142 32852 26148 32864
rect 26200 32852 26206 32904
rect 26973 32895 27031 32901
rect 26973 32861 26985 32895
rect 27019 32892 27031 32895
rect 27246 32892 27252 32904
rect 27019 32864 27252 32892
rect 27019 32861 27031 32864
rect 26973 32855 27031 32861
rect 27246 32852 27252 32864
rect 27304 32852 27310 32904
rect 28721 32895 28779 32901
rect 27816 32864 28120 32892
rect 25774 32824 25780 32836
rect 22060 32796 22784 32824
rect 25735 32796 25780 32824
rect 22060 32784 22066 32796
rect 25774 32784 25780 32796
rect 25832 32784 25838 32836
rect 27816 32833 27844 32864
rect 27801 32827 27859 32833
rect 27801 32793 27813 32827
rect 27847 32793 27859 32827
rect 27801 32787 27859 32793
rect 27982 32784 27988 32836
rect 28040 32833 28046 32836
rect 28040 32827 28059 32833
rect 28047 32793 28059 32827
rect 28092 32824 28120 32864
rect 28721 32861 28733 32895
rect 28767 32892 28779 32895
rect 28994 32892 29000 32904
rect 28767 32864 29000 32892
rect 28767 32861 28779 32864
rect 28721 32855 28779 32861
rect 28994 32852 29000 32864
rect 29052 32892 29058 32904
rect 29549 32895 29607 32901
rect 29549 32892 29561 32895
rect 29052 32864 29561 32892
rect 29052 32852 29058 32864
rect 29549 32861 29561 32864
rect 29595 32861 29607 32895
rect 29549 32855 29607 32861
rect 30374 32852 30380 32904
rect 30432 32892 30438 32904
rect 30852 32901 30880 32932
rect 31294 32920 31300 32932
rect 31352 32920 31358 32972
rect 32950 32960 32956 32972
rect 32911 32932 32956 32960
rect 32950 32920 32956 32932
rect 33008 32920 33014 32972
rect 33502 32920 33508 32972
rect 33560 32960 33566 32972
rect 33689 32963 33747 32969
rect 33689 32960 33701 32963
rect 33560 32932 33701 32960
rect 33560 32920 33566 32932
rect 33689 32929 33701 32932
rect 33735 32929 33747 32963
rect 33689 32923 33747 32929
rect 30745 32895 30803 32901
rect 30745 32892 30757 32895
rect 30432 32864 30757 32892
rect 30432 32852 30438 32864
rect 30745 32861 30757 32864
rect 30791 32861 30803 32895
rect 30745 32855 30803 32861
rect 30837 32895 30895 32901
rect 30837 32861 30849 32895
rect 30883 32861 30895 32895
rect 30837 32855 30895 32861
rect 31021 32895 31079 32901
rect 31021 32861 31033 32895
rect 31067 32861 31079 32895
rect 31021 32855 31079 32861
rect 31113 32895 31171 32901
rect 31113 32861 31125 32895
rect 31159 32892 31171 32895
rect 31202 32892 31208 32904
rect 31159 32864 31208 32892
rect 31159 32861 31171 32864
rect 31113 32855 31171 32861
rect 29178 32824 29184 32836
rect 28092 32796 29184 32824
rect 28040 32787 28059 32793
rect 28040 32784 28046 32787
rect 29178 32784 29184 32796
rect 29236 32784 29242 32836
rect 29638 32784 29644 32836
rect 29696 32824 29702 32836
rect 31036 32824 31064 32855
rect 31202 32852 31208 32864
rect 31260 32852 31266 32904
rect 32674 32892 32680 32904
rect 32635 32864 32680 32892
rect 32674 32852 32680 32864
rect 32732 32852 32738 32904
rect 33410 32892 33416 32904
rect 33371 32864 33416 32892
rect 33410 32852 33416 32864
rect 33468 32852 33474 32904
rect 33594 32892 33600 32904
rect 33555 32864 33600 32892
rect 33594 32852 33600 32864
rect 33652 32852 33658 32904
rect 33781 32895 33839 32901
rect 33781 32861 33793 32895
rect 33827 32861 33839 32895
rect 33781 32855 33839 32861
rect 29696 32796 31064 32824
rect 33796 32824 33824 32855
rect 33870 32852 33876 32904
rect 33928 32892 33934 32904
rect 33980 32901 34008 33000
rect 47118 32960 47124 32972
rect 47079 32932 47124 32960
rect 47118 32920 47124 32932
rect 47176 32920 47182 32972
rect 47394 32960 47400 32972
rect 47355 32932 47400 32960
rect 47394 32920 47400 32932
rect 47452 32920 47458 32972
rect 33965 32895 34023 32901
rect 33965 32892 33977 32895
rect 33928 32864 33977 32892
rect 33928 32852 33934 32864
rect 33965 32861 33977 32864
rect 34011 32861 34023 32895
rect 33965 32855 34023 32861
rect 34698 32852 34704 32904
rect 34756 32892 34762 32904
rect 35253 32895 35311 32901
rect 35253 32892 35265 32895
rect 34756 32864 35265 32892
rect 34756 32852 34762 32864
rect 35253 32861 35265 32864
rect 35299 32861 35311 32895
rect 35253 32855 35311 32861
rect 46290 32852 46296 32904
rect 46348 32892 46354 32904
rect 46569 32895 46627 32901
rect 46569 32892 46581 32895
rect 46348 32864 46581 32892
rect 46348 32852 46354 32864
rect 46569 32861 46581 32864
rect 46615 32861 46627 32895
rect 46569 32855 46627 32861
rect 46474 32824 46480 32836
rect 33796 32796 46480 32824
rect 29696 32784 29702 32796
rect 46474 32784 46480 32796
rect 46532 32784 46538 32836
rect 47213 32827 47271 32833
rect 47213 32793 47225 32827
rect 47259 32824 47271 32827
rect 47302 32824 47308 32836
rect 47259 32796 47308 32824
rect 47259 32793 47271 32796
rect 47213 32787 47271 32793
rect 47302 32784 47308 32796
rect 47360 32784 47366 32836
rect 22186 32756 22192 32768
rect 21560 32728 22192 32756
rect 11977 32719 12035 32725
rect 22186 32716 22192 32728
rect 22244 32716 22250 32768
rect 23198 32716 23204 32768
rect 23256 32756 23262 32768
rect 24765 32759 24823 32765
rect 24765 32756 24777 32759
rect 23256 32728 24777 32756
rect 23256 32716 23262 32728
rect 24765 32725 24777 32728
rect 24811 32725 24823 32759
rect 26234 32756 26240 32768
rect 26195 32728 26240 32756
rect 24765 32719 24823 32725
rect 26234 32716 26240 32728
rect 26292 32716 26298 32768
rect 27430 32716 27436 32768
rect 27488 32756 27494 32768
rect 28169 32759 28227 32765
rect 28169 32756 28181 32759
rect 27488 32728 28181 32756
rect 27488 32716 27494 32728
rect 28169 32725 28181 32728
rect 28215 32725 28227 32759
rect 28169 32719 28227 32725
rect 28534 32716 28540 32768
rect 28592 32756 28598 32768
rect 28905 32759 28963 32765
rect 28905 32756 28917 32759
rect 28592 32728 28917 32756
rect 28592 32716 28598 32728
rect 28905 32725 28917 32728
rect 28951 32725 28963 32759
rect 28905 32719 28963 32725
rect 29362 32716 29368 32768
rect 29420 32756 29426 32768
rect 29733 32759 29791 32765
rect 29733 32756 29745 32759
rect 29420 32728 29745 32756
rect 29420 32716 29426 32728
rect 29733 32725 29745 32728
rect 29779 32725 29791 32759
rect 29733 32719 29791 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 14277 32555 14335 32561
rect 14277 32521 14289 32555
rect 14323 32552 14335 32555
rect 14366 32552 14372 32564
rect 14323 32524 14372 32552
rect 14323 32521 14335 32524
rect 14277 32515 14335 32521
rect 14366 32512 14372 32524
rect 14424 32512 14430 32564
rect 22373 32555 22431 32561
rect 22373 32521 22385 32555
rect 22419 32552 22431 32555
rect 22462 32552 22468 32564
rect 22419 32524 22468 32552
rect 22419 32521 22431 32524
rect 22373 32515 22431 32521
rect 22462 32512 22468 32524
rect 22520 32512 22526 32564
rect 23382 32552 23388 32564
rect 23343 32524 23388 32552
rect 23382 32512 23388 32524
rect 23440 32512 23446 32564
rect 28534 32552 28540 32564
rect 24596 32524 28540 32552
rect 24596 32496 24624 32524
rect 28534 32512 28540 32524
rect 28592 32512 28598 32564
rect 29270 32552 29276 32564
rect 28644 32524 29276 32552
rect 2682 32484 2688 32496
rect 2643 32456 2688 32484
rect 2682 32444 2688 32456
rect 2740 32444 2746 32496
rect 11790 32484 11796 32496
rect 11751 32456 11796 32484
rect 11790 32444 11796 32456
rect 11848 32444 11854 32496
rect 12802 32444 12808 32496
rect 12860 32444 12866 32496
rect 22646 32444 22652 32496
rect 22704 32484 22710 32496
rect 24578 32484 24584 32496
rect 22704 32456 24584 32484
rect 22704 32444 22710 32456
rect 24578 32444 24584 32456
rect 24636 32444 24642 32496
rect 25130 32444 25136 32496
rect 25188 32484 25194 32496
rect 25317 32487 25375 32493
rect 25317 32484 25329 32487
rect 25188 32456 25329 32484
rect 25188 32444 25194 32456
rect 25317 32453 25329 32456
rect 25363 32453 25375 32487
rect 25317 32447 25375 32453
rect 26050 32444 26056 32496
rect 26108 32484 26114 32496
rect 27982 32484 27988 32496
rect 26108 32456 27988 32484
rect 26108 32444 26114 32456
rect 27982 32444 27988 32456
rect 28040 32444 28046 32496
rect 28644 32493 28672 32524
rect 29270 32512 29276 32524
rect 29328 32552 29334 32564
rect 29546 32552 29552 32564
rect 29328 32524 29552 32552
rect 29328 32512 29334 32524
rect 29546 32512 29552 32524
rect 29604 32512 29610 32564
rect 29638 32512 29644 32564
rect 29696 32552 29702 32564
rect 30193 32555 30251 32561
rect 30193 32552 30205 32555
rect 29696 32524 30205 32552
rect 29696 32512 29702 32524
rect 30193 32521 30205 32524
rect 30239 32521 30251 32555
rect 30193 32515 30251 32521
rect 33410 32512 33416 32564
rect 33468 32552 33474 32564
rect 33597 32555 33655 32561
rect 33597 32552 33609 32555
rect 33468 32524 33609 32552
rect 33468 32512 33474 32524
rect 33597 32521 33609 32524
rect 33643 32521 33655 32555
rect 37642 32552 37648 32564
rect 37603 32524 37648 32552
rect 33597 32515 33655 32521
rect 37642 32512 37648 32524
rect 37700 32512 37706 32564
rect 28629 32487 28687 32493
rect 28629 32453 28641 32487
rect 28675 32453 28687 32487
rect 28629 32447 28687 32453
rect 28810 32444 28816 32496
rect 28868 32484 28874 32496
rect 28994 32484 29000 32496
rect 28868 32456 29000 32484
rect 28868 32444 28874 32456
rect 28994 32444 29000 32456
rect 29052 32444 29058 32496
rect 29273 32453 29331 32459
rect 29273 32450 29285 32453
rect 29196 32440 29285 32450
rect 13538 32376 13544 32428
rect 13596 32416 13602 32428
rect 14185 32419 14243 32425
rect 14185 32416 14197 32419
rect 13596 32388 14197 32416
rect 13596 32376 13602 32388
rect 14185 32385 14197 32388
rect 14231 32385 14243 32419
rect 14185 32379 14243 32385
rect 21726 32376 21732 32428
rect 21784 32416 21790 32428
rect 22002 32416 22008 32428
rect 21784 32388 22008 32416
rect 21784 32376 21790 32388
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22370 32376 22376 32428
rect 22428 32416 22434 32428
rect 22833 32419 22891 32425
rect 22833 32416 22845 32419
rect 22428 32388 22845 32416
rect 22428 32376 22434 32388
rect 22833 32385 22845 32388
rect 22879 32385 22891 32419
rect 22833 32379 22891 32385
rect 24946 32376 24952 32428
rect 25004 32416 25010 32428
rect 25593 32419 25651 32425
rect 25593 32416 25605 32419
rect 25004 32388 25605 32416
rect 25004 32376 25010 32388
rect 25593 32385 25605 32388
rect 25639 32385 25651 32419
rect 28902 32416 28908 32428
rect 25593 32379 25651 32385
rect 27265 32388 28908 32416
rect 2501 32351 2559 32357
rect 2501 32317 2513 32351
rect 2547 32317 2559 32351
rect 3234 32348 3240 32360
rect 3195 32320 3240 32348
rect 2501 32311 2559 32317
rect 2516 32280 2544 32311
rect 3234 32308 3240 32320
rect 3292 32308 3298 32360
rect 11514 32348 11520 32360
rect 11475 32320 11520 32348
rect 11514 32308 11520 32320
rect 11572 32308 11578 32360
rect 14090 32348 14096 32360
rect 11624 32320 14096 32348
rect 2516 32252 6914 32280
rect 1946 32172 1952 32224
rect 2004 32212 2010 32224
rect 2041 32215 2099 32221
rect 2041 32212 2053 32215
rect 2004 32184 2053 32212
rect 2004 32172 2010 32184
rect 2041 32181 2053 32184
rect 2087 32181 2099 32215
rect 6886 32212 6914 32252
rect 9398 32240 9404 32292
rect 9456 32280 9462 32292
rect 11624 32280 11652 32320
rect 14090 32308 14096 32320
rect 14148 32308 14154 32360
rect 22097 32351 22155 32357
rect 22097 32317 22109 32351
rect 22143 32348 22155 32351
rect 22462 32348 22468 32360
rect 22143 32320 22468 32348
rect 22143 32317 22155 32320
rect 22097 32311 22155 32317
rect 22462 32308 22468 32320
rect 22520 32308 22526 32360
rect 23106 32308 23112 32360
rect 23164 32348 23170 32360
rect 25501 32351 25559 32357
rect 23164 32320 23209 32348
rect 23164 32308 23170 32320
rect 25501 32317 25513 32351
rect 25547 32348 25559 32351
rect 25866 32348 25872 32360
rect 25547 32320 25872 32348
rect 25547 32317 25559 32320
rect 25501 32311 25559 32317
rect 25866 32308 25872 32320
rect 25924 32348 25930 32360
rect 27265 32348 27293 32388
rect 28902 32376 28908 32388
rect 28960 32416 28966 32428
rect 29104 32422 29285 32440
rect 29104 32416 29224 32422
rect 28960 32412 29224 32416
rect 29273 32419 29285 32422
rect 29319 32419 29331 32453
rect 29454 32444 29460 32496
rect 29512 32493 29518 32496
rect 29512 32484 29523 32493
rect 32582 32484 32588 32496
rect 29512 32456 29557 32484
rect 30208 32456 32588 32484
rect 29512 32447 29523 32456
rect 29512 32444 29518 32447
rect 29273 32413 29331 32419
rect 28960 32388 29132 32412
rect 28960 32376 28966 32388
rect 30098 32376 30104 32428
rect 30156 32425 30162 32428
rect 30156 32416 30165 32425
rect 30208 32416 30236 32456
rect 32582 32444 32588 32456
rect 32640 32444 32646 32496
rect 32950 32444 32956 32496
rect 33008 32484 33014 32496
rect 33008 32456 33456 32484
rect 33008 32444 33014 32456
rect 30285 32419 30343 32425
rect 30156 32388 30249 32416
rect 30156 32379 30165 32388
rect 30285 32385 30297 32419
rect 30331 32385 30343 32419
rect 31202 32416 31208 32428
rect 31163 32388 31208 32416
rect 30285 32379 30343 32385
rect 30156 32376 30162 32379
rect 25924 32320 27293 32348
rect 28813 32351 28871 32357
rect 25924 32308 25930 32320
rect 28813 32317 28825 32351
rect 28859 32348 28871 32351
rect 29178 32348 29184 32360
rect 28859 32320 29184 32348
rect 28859 32317 28871 32320
rect 28813 32311 28871 32317
rect 29178 32308 29184 32320
rect 29236 32308 29242 32360
rect 29638 32348 29644 32360
rect 29551 32320 29644 32348
rect 29638 32308 29644 32320
rect 29696 32348 29702 32360
rect 30300 32348 30328 32379
rect 31202 32376 31208 32388
rect 31260 32376 31266 32428
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32416 32367 32419
rect 33226 32416 33232 32428
rect 32355 32388 32628 32416
rect 33187 32388 33232 32416
rect 32355 32385 32367 32388
rect 32309 32379 32367 32385
rect 32600 32360 32628 32388
rect 33226 32376 33232 32388
rect 33284 32376 33290 32428
rect 33428 32425 33456 32456
rect 45922 32444 45928 32496
rect 45980 32484 45986 32496
rect 45980 32456 47532 32484
rect 45980 32444 45986 32456
rect 47504 32428 47532 32456
rect 33413 32419 33471 32425
rect 33413 32385 33425 32419
rect 33459 32385 33471 32419
rect 33413 32379 33471 32385
rect 36633 32419 36691 32425
rect 36633 32385 36645 32419
rect 36679 32416 36691 32419
rect 46474 32416 46480 32428
rect 36679 32388 37320 32416
rect 46435 32388 46480 32416
rect 36679 32385 36691 32388
rect 36633 32379 36691 32385
rect 32398 32348 32404 32360
rect 29696 32320 32404 32348
rect 29696 32308 29702 32320
rect 32398 32308 32404 32320
rect 32456 32308 32462 32360
rect 32582 32308 32588 32360
rect 32640 32308 32646 32360
rect 22002 32280 22008 32292
rect 9456 32252 11652 32280
rect 12820 32252 22008 32280
rect 9456 32240 9462 32252
rect 12820 32212 12848 32252
rect 22002 32240 22008 32252
rect 22060 32240 22066 32292
rect 22646 32240 22652 32292
rect 22704 32280 22710 32292
rect 25777 32283 25835 32289
rect 25777 32280 25789 32283
rect 22704 32252 25789 32280
rect 22704 32240 22710 32252
rect 25777 32249 25789 32252
rect 25823 32249 25835 32283
rect 25777 32243 25835 32249
rect 26786 32240 26792 32292
rect 26844 32280 26850 32292
rect 27522 32280 27528 32292
rect 26844 32252 27528 32280
rect 26844 32240 26850 32252
rect 27522 32240 27528 32252
rect 27580 32240 27586 32292
rect 27982 32240 27988 32292
rect 28040 32280 28046 32292
rect 29454 32280 29460 32292
rect 28040 32252 29460 32280
rect 28040 32240 28046 32252
rect 29454 32240 29460 32252
rect 29512 32240 29518 32292
rect 29822 32240 29828 32292
rect 29880 32280 29886 32292
rect 31389 32283 31447 32289
rect 31389 32280 31401 32283
rect 29880 32252 31401 32280
rect 29880 32240 29886 32252
rect 31389 32249 31401 32252
rect 31435 32280 31447 32283
rect 33594 32280 33600 32292
rect 31435 32252 33600 32280
rect 31435 32249 31447 32252
rect 31389 32243 31447 32249
rect 33594 32240 33600 32252
rect 33652 32240 33658 32292
rect 34514 32240 34520 32292
rect 34572 32280 34578 32292
rect 37292 32289 37320 32388
rect 46474 32376 46480 32388
rect 46532 32376 46538 32428
rect 47486 32376 47492 32428
rect 47544 32416 47550 32428
rect 47581 32419 47639 32425
rect 47581 32416 47593 32419
rect 47544 32388 47593 32416
rect 47544 32376 47550 32388
rect 47581 32385 47593 32388
rect 47627 32385 47639 32419
rect 47581 32379 47639 32385
rect 37734 32348 37740 32360
rect 37695 32320 37740 32348
rect 37734 32308 37740 32320
rect 37792 32308 37798 32360
rect 37829 32351 37887 32357
rect 37829 32317 37841 32351
rect 37875 32317 37887 32351
rect 46198 32348 46204 32360
rect 46159 32320 46204 32348
rect 37829 32311 37887 32317
rect 37277 32283 37335 32289
rect 34572 32252 36860 32280
rect 34572 32240 34578 32252
rect 13262 32212 13268 32224
rect 6886 32184 12848 32212
rect 13175 32184 13268 32212
rect 2041 32175 2099 32181
rect 13262 32172 13268 32184
rect 13320 32212 13326 32224
rect 13722 32212 13728 32224
rect 13320 32184 13728 32212
rect 13320 32172 13326 32184
rect 13722 32172 13728 32184
rect 13780 32172 13786 32224
rect 23198 32212 23204 32224
rect 23159 32184 23204 32212
rect 23198 32172 23204 32184
rect 23256 32172 23262 32224
rect 25593 32215 25651 32221
rect 25593 32181 25605 32215
rect 25639 32212 25651 32215
rect 27798 32212 27804 32224
rect 25639 32184 27804 32212
rect 25639 32181 25651 32184
rect 25593 32175 25651 32181
rect 27798 32172 27804 32184
rect 27856 32172 27862 32224
rect 28534 32172 28540 32224
rect 28592 32212 28598 32224
rect 31018 32212 31024 32224
rect 28592 32184 31024 32212
rect 28592 32172 28598 32184
rect 31018 32172 31024 32184
rect 31076 32172 31082 32224
rect 31754 32172 31760 32224
rect 31812 32212 31818 32224
rect 32677 32215 32735 32221
rect 32677 32212 32689 32215
rect 31812 32184 32689 32212
rect 31812 32172 31818 32184
rect 32677 32181 32689 32184
rect 32723 32181 32735 32215
rect 32677 32175 32735 32181
rect 36170 32172 36176 32224
rect 36228 32212 36234 32224
rect 36449 32215 36507 32221
rect 36449 32212 36461 32215
rect 36228 32184 36461 32212
rect 36228 32172 36234 32184
rect 36449 32181 36461 32184
rect 36495 32181 36507 32215
rect 36832 32212 36860 32252
rect 37277 32249 37289 32283
rect 37323 32249 37335 32283
rect 37277 32243 37335 32249
rect 37844 32212 37872 32311
rect 46198 32308 46204 32320
rect 46256 32308 46262 32360
rect 36832 32184 37872 32212
rect 36449 32175 36507 32181
rect 46474 32172 46480 32224
rect 46532 32212 46538 32224
rect 47673 32215 47731 32221
rect 47673 32212 47685 32215
rect 46532 32184 47685 32212
rect 46532 32172 46538 32184
rect 47673 32181 47685 32184
rect 47719 32181 47731 32215
rect 47673 32175 47731 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1397 32011 1455 32017
rect 1397 31977 1409 32011
rect 1443 32008 1455 32011
rect 2774 32008 2780 32020
rect 1443 31980 2780 32008
rect 1443 31977 1455 31980
rect 1397 31971 1455 31977
rect 2774 31968 2780 31980
rect 2832 31968 2838 32020
rect 8294 31968 8300 32020
rect 8352 32008 8358 32020
rect 9858 32008 9864 32020
rect 8352 31980 9864 32008
rect 8352 31968 8358 31980
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 11698 31968 11704 32020
rect 11756 32008 11762 32020
rect 12069 32011 12127 32017
rect 12069 32008 12081 32011
rect 11756 31980 12081 32008
rect 11756 31968 11762 31980
rect 12069 31977 12081 31980
rect 12115 31977 12127 32011
rect 12069 31971 12127 31977
rect 12713 32011 12771 32017
rect 12713 31977 12725 32011
rect 12759 32008 12771 32011
rect 12802 32008 12808 32020
rect 12759 31980 12808 32008
rect 12759 31977 12771 31980
rect 12713 31971 12771 31977
rect 12802 31968 12808 31980
rect 12860 31968 12866 32020
rect 25498 32008 25504 32020
rect 16546 31980 25504 32008
rect 3050 31900 3056 31952
rect 3108 31940 3114 31952
rect 16546 31940 16574 31980
rect 25498 31968 25504 31980
rect 25556 31968 25562 32020
rect 25700 31980 29224 32008
rect 3108 31912 16574 31940
rect 3108 31900 3114 31912
rect 23566 31900 23572 31952
rect 23624 31940 23630 31952
rect 23624 31912 25268 31940
rect 23624 31900 23630 31912
rect 9398 31872 9404 31884
rect 9359 31844 9404 31872
rect 9398 31832 9404 31844
rect 9456 31832 9462 31884
rect 9585 31875 9643 31881
rect 9585 31841 9597 31875
rect 9631 31872 9643 31875
rect 9766 31872 9772 31884
rect 9631 31844 9772 31872
rect 9631 31841 9643 31844
rect 9585 31835 9643 31841
rect 9766 31832 9772 31844
rect 9824 31832 9830 31884
rect 9858 31832 9864 31884
rect 9916 31872 9922 31884
rect 12894 31872 12900 31884
rect 9916 31844 9961 31872
rect 11992 31844 12900 31872
rect 9916 31832 9922 31844
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 2777 31807 2835 31813
rect 2777 31773 2789 31807
rect 2823 31804 2835 31807
rect 3050 31804 3056 31816
rect 2823 31776 3056 31804
rect 2823 31773 2835 31776
rect 2777 31767 2835 31773
rect 3050 31764 3056 31776
rect 3108 31764 3114 31816
rect 11992 31813 12020 31844
rect 12894 31832 12900 31844
rect 12952 31832 12958 31884
rect 15105 31875 15163 31881
rect 15105 31841 15117 31875
rect 15151 31872 15163 31875
rect 15194 31872 15200 31884
rect 15151 31844 15200 31872
rect 15151 31841 15163 31844
rect 15105 31835 15163 31841
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 20806 31872 20812 31884
rect 20272 31844 20812 31872
rect 11977 31807 12035 31813
rect 11977 31773 11989 31807
rect 12023 31773 12035 31807
rect 11977 31767 12035 31773
rect 12161 31807 12219 31813
rect 12161 31773 12173 31807
rect 12207 31804 12219 31807
rect 12618 31804 12624 31816
rect 12207 31776 12480 31804
rect 12579 31776 12624 31804
rect 12207 31773 12219 31776
rect 12161 31767 12219 31773
rect 12452 31736 12480 31776
rect 12618 31764 12624 31776
rect 12676 31764 12682 31816
rect 15013 31807 15071 31813
rect 15013 31773 15025 31807
rect 15059 31804 15071 31807
rect 16574 31804 16580 31816
rect 15059 31776 16580 31804
rect 15059 31773 15071 31776
rect 15013 31767 15071 31773
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 20272 31813 20300 31844
rect 20806 31832 20812 31844
rect 20864 31872 20870 31884
rect 24762 31872 24768 31884
rect 20864 31844 20944 31872
rect 20864 31832 20870 31844
rect 20257 31807 20315 31813
rect 20257 31773 20269 31807
rect 20303 31773 20315 31807
rect 20257 31767 20315 31773
rect 20349 31807 20407 31813
rect 20349 31773 20361 31807
rect 20395 31804 20407 31807
rect 20438 31804 20444 31816
rect 20395 31776 20444 31804
rect 20395 31773 20407 31776
rect 20349 31767 20407 31773
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 20916 31813 20944 31844
rect 22020 31844 24768 31872
rect 22020 31813 22048 31844
rect 24762 31832 24768 31844
rect 24820 31832 24826 31884
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31773 20959 31807
rect 20901 31767 20959 31773
rect 22005 31807 22063 31813
rect 22005 31773 22017 31807
rect 22051 31773 22063 31807
rect 22005 31767 22063 31773
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31804 22339 31807
rect 22370 31804 22376 31816
rect 22327 31776 22376 31804
rect 22327 31773 22339 31776
rect 22281 31767 22339 31773
rect 22370 31764 22376 31776
rect 22428 31764 22434 31816
rect 22646 31764 22652 31816
rect 22704 31764 22710 31816
rect 23658 31764 23664 31816
rect 23716 31804 23722 31816
rect 24670 31804 24676 31816
rect 23716 31776 24676 31804
rect 23716 31764 23722 31776
rect 24670 31764 24676 31776
rect 24728 31764 24734 31816
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31773 24915 31807
rect 24857 31767 24915 31773
rect 25133 31807 25191 31813
rect 25133 31773 25145 31807
rect 25179 31804 25191 31807
rect 25240 31804 25268 31912
rect 25700 31872 25728 31980
rect 27982 31940 27988 31952
rect 27943 31912 27988 31940
rect 27982 31900 27988 31912
rect 28040 31900 28046 31952
rect 28074 31900 28080 31952
rect 28132 31940 28138 31952
rect 28626 31940 28632 31952
rect 28132 31912 28632 31940
rect 28132 31900 28138 31912
rect 28626 31900 28632 31912
rect 28684 31940 28690 31952
rect 28721 31943 28779 31949
rect 28721 31940 28733 31943
rect 28684 31912 28733 31940
rect 28684 31900 28690 31912
rect 28721 31909 28733 31912
rect 28767 31909 28779 31943
rect 28721 31903 28779 31909
rect 25958 31872 25964 31884
rect 25179 31776 25268 31804
rect 25516 31844 25728 31872
rect 25884 31844 25964 31872
rect 25179 31773 25191 31776
rect 25133 31767 25191 31773
rect 12526 31736 12532 31748
rect 12452 31708 12532 31736
rect 12526 31696 12532 31708
rect 12584 31696 12590 31748
rect 22664 31736 22692 31764
rect 22020 31708 22692 31736
rect 22020 31680 22048 31708
rect 2866 31668 2872 31680
rect 2827 31640 2872 31668
rect 2866 31628 2872 31640
rect 2924 31628 2930 31680
rect 15378 31668 15384 31680
rect 15339 31640 15384 31668
rect 15378 31628 15384 31640
rect 15436 31628 15442 31680
rect 20806 31628 20812 31680
rect 20864 31668 20870 31680
rect 20993 31671 21051 31677
rect 20993 31668 21005 31671
rect 20864 31640 21005 31668
rect 20864 31628 20870 31640
rect 20993 31637 21005 31640
rect 21039 31637 21051 31671
rect 20993 31631 21051 31637
rect 21821 31671 21879 31677
rect 21821 31637 21833 31671
rect 21867 31668 21879 31671
rect 21910 31668 21916 31680
rect 21867 31640 21916 31668
rect 21867 31637 21879 31640
rect 21821 31631 21879 31637
rect 21910 31628 21916 31640
rect 21968 31628 21974 31680
rect 22002 31628 22008 31680
rect 22060 31628 22066 31680
rect 22186 31628 22192 31680
rect 22244 31668 22250 31680
rect 24394 31668 24400 31680
rect 22244 31640 24400 31668
rect 22244 31628 22250 31640
rect 24394 31628 24400 31640
rect 24452 31628 24458 31680
rect 24486 31628 24492 31680
rect 24544 31668 24550 31680
rect 24673 31671 24731 31677
rect 24673 31668 24685 31671
rect 24544 31640 24685 31668
rect 24544 31628 24550 31640
rect 24673 31637 24685 31640
rect 24719 31637 24731 31671
rect 24872 31668 24900 31767
rect 25041 31739 25099 31745
rect 25041 31705 25053 31739
rect 25087 31736 25099 31739
rect 25516 31736 25544 31844
rect 25682 31804 25688 31816
rect 25643 31776 25688 31804
rect 25682 31764 25688 31776
rect 25740 31764 25746 31816
rect 25884 31813 25912 31844
rect 25958 31832 25964 31844
rect 26016 31832 26022 31884
rect 29086 31872 29092 31884
rect 28552 31844 29092 31872
rect 25869 31807 25927 31813
rect 25869 31773 25881 31807
rect 25915 31773 25927 31807
rect 25869 31767 25927 31773
rect 26099 31807 26157 31813
rect 26099 31773 26111 31807
rect 26145 31804 26157 31807
rect 26786 31804 26792 31816
rect 26145 31776 26792 31804
rect 26145 31773 26157 31776
rect 26099 31767 26157 31773
rect 26786 31764 26792 31776
rect 26844 31804 26850 31816
rect 26970 31804 26976 31816
rect 26844 31776 26976 31804
rect 26844 31764 26850 31776
rect 26970 31764 26976 31776
rect 27028 31764 27034 31816
rect 27798 31804 27804 31816
rect 27759 31776 27804 31804
rect 27798 31764 27804 31776
rect 27856 31764 27862 31816
rect 28552 31813 28580 31844
rect 29086 31832 29092 31844
rect 29144 31832 29150 31884
rect 29196 31872 29224 31980
rect 33045 31943 33103 31949
rect 31772 31912 32996 31940
rect 31772 31872 31800 31912
rect 29196 31844 31800 31872
rect 31849 31875 31907 31881
rect 31849 31841 31861 31875
rect 31895 31872 31907 31875
rect 31895 31844 32444 31872
rect 31895 31841 31907 31844
rect 31849 31835 31907 31841
rect 28537 31807 28595 31813
rect 28537 31773 28549 31807
rect 28583 31773 28595 31807
rect 28537 31767 28595 31773
rect 29196 31776 30420 31804
rect 25087 31708 25544 31736
rect 25087 31705 25099 31708
rect 25041 31699 25099 31705
rect 25774 31696 25780 31748
rect 25832 31736 25838 31748
rect 25961 31739 26019 31745
rect 25961 31736 25973 31739
rect 25832 31708 25973 31736
rect 25832 31696 25838 31708
rect 25961 31705 25973 31708
rect 26007 31705 26019 31739
rect 25961 31699 26019 31705
rect 27062 31696 27068 31748
rect 27120 31736 27126 31748
rect 29196 31736 29224 31776
rect 27120 31708 29224 31736
rect 27120 31696 27126 31708
rect 26237 31671 26295 31677
rect 26237 31668 26249 31671
rect 24872 31640 26249 31668
rect 24673 31631 24731 31637
rect 26237 31637 26249 31640
rect 26283 31637 26295 31671
rect 30392 31668 30420 31776
rect 30466 31764 30472 31816
rect 30524 31804 30530 31816
rect 31202 31804 31208 31816
rect 30524 31776 31208 31804
rect 30524 31764 30530 31776
rect 31202 31764 31208 31776
rect 31260 31804 31266 31816
rect 31754 31804 31760 31816
rect 31260 31776 31616 31804
rect 31715 31776 31760 31804
rect 31260 31764 31266 31776
rect 31588 31736 31616 31776
rect 31754 31764 31760 31776
rect 31812 31764 31818 31816
rect 32416 31813 32444 31844
rect 32674 31832 32680 31884
rect 32732 31832 32738 31884
rect 32582 31813 32588 31816
rect 31941 31807 31999 31813
rect 31941 31804 31953 31807
rect 31864 31776 31953 31804
rect 31864 31736 31892 31776
rect 31941 31773 31953 31776
rect 31987 31773 31999 31807
rect 31941 31767 31999 31773
rect 32401 31807 32459 31813
rect 32401 31773 32413 31807
rect 32447 31773 32459 31807
rect 32401 31767 32459 31773
rect 32549 31807 32588 31813
rect 32549 31773 32561 31807
rect 32549 31767 32588 31773
rect 32582 31764 32588 31767
rect 32640 31764 32646 31816
rect 32692 31804 32720 31832
rect 32866 31807 32924 31813
rect 32866 31804 32878 31807
rect 32692 31776 32878 31804
rect 32866 31773 32878 31776
rect 32912 31773 32924 31807
rect 32866 31767 32924 31773
rect 31588 31708 31892 31736
rect 32214 31696 32220 31748
rect 32272 31736 32278 31748
rect 32677 31739 32735 31745
rect 32677 31736 32689 31739
rect 32272 31708 32689 31736
rect 32272 31696 32278 31708
rect 32677 31705 32689 31708
rect 32723 31705 32735 31739
rect 32677 31699 32735 31705
rect 32766 31696 32772 31748
rect 32824 31736 32830 31748
rect 32968 31736 32996 31912
rect 33045 31909 33057 31943
rect 33091 31940 33103 31943
rect 33410 31940 33416 31952
rect 33091 31912 33416 31940
rect 33091 31909 33103 31912
rect 33045 31903 33103 31909
rect 33410 31900 33416 31912
rect 33468 31900 33474 31952
rect 33686 31832 33692 31884
rect 33744 31872 33750 31884
rect 35897 31875 35955 31881
rect 35897 31872 35909 31875
rect 33744 31844 35909 31872
rect 33744 31832 33750 31844
rect 35897 31841 35909 31844
rect 35943 31841 35955 31875
rect 36170 31872 36176 31884
rect 36131 31844 36176 31872
rect 35897 31835 35955 31841
rect 36170 31832 36176 31844
rect 36228 31832 36234 31884
rect 36630 31832 36636 31884
rect 36688 31872 36694 31884
rect 37645 31875 37703 31881
rect 37645 31872 37657 31875
rect 36688 31844 37657 31872
rect 36688 31832 36694 31844
rect 37645 31841 37657 31844
rect 37691 31841 37703 31875
rect 46290 31872 46296 31884
rect 46251 31844 46296 31872
rect 37645 31835 37703 31841
rect 46290 31832 46296 31844
rect 46348 31832 46354 31884
rect 46474 31872 46480 31884
rect 46435 31844 46480 31872
rect 46474 31832 46480 31844
rect 46532 31832 46538 31884
rect 48130 31872 48136 31884
rect 48091 31844 48136 31872
rect 48130 31832 48136 31844
rect 48188 31832 48194 31884
rect 34698 31804 34704 31816
rect 34659 31776 34704 31804
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 34790 31764 34796 31816
rect 34848 31804 34854 31816
rect 34848 31776 34893 31804
rect 34848 31764 34854 31776
rect 37458 31736 37464 31748
rect 32824 31708 32996 31736
rect 37398 31708 37464 31736
rect 32824 31696 32830 31708
rect 37458 31696 37464 31708
rect 37516 31696 37522 31748
rect 32950 31668 32956 31680
rect 30392 31640 32956 31668
rect 26237 31631 26295 31637
rect 32950 31628 32956 31640
rect 33008 31668 33014 31680
rect 37550 31668 37556 31680
rect 33008 31640 37556 31668
rect 33008 31628 33014 31640
rect 37550 31628 37556 31640
rect 37608 31628 37614 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 9766 31464 9772 31476
rect 9727 31436 9772 31464
rect 9766 31424 9772 31436
rect 9824 31424 9830 31476
rect 11514 31424 11520 31476
rect 11572 31464 11578 31476
rect 11609 31467 11667 31473
rect 11609 31464 11621 31467
rect 11572 31436 11621 31464
rect 11572 31424 11578 31436
rect 11609 31433 11621 31436
rect 11655 31433 11667 31467
rect 11609 31427 11667 31433
rect 14090 31424 14096 31476
rect 14148 31464 14154 31476
rect 15381 31467 15439 31473
rect 15381 31464 15393 31467
rect 14148 31436 15393 31464
rect 14148 31424 14154 31436
rect 15381 31433 15393 31436
rect 15427 31433 15439 31467
rect 15381 31427 15439 31433
rect 25498 31424 25504 31476
rect 25556 31464 25562 31476
rect 26418 31464 26424 31476
rect 25556 31436 26424 31464
rect 25556 31424 25562 31436
rect 26418 31424 26424 31436
rect 26476 31424 26482 31476
rect 32582 31424 32588 31476
rect 32640 31464 32646 31476
rect 34885 31467 34943 31473
rect 34885 31464 34897 31467
rect 32640 31436 34897 31464
rect 32640 31424 32646 31436
rect 34885 31433 34897 31436
rect 34931 31433 34943 31467
rect 34885 31427 34943 31433
rect 37369 31467 37427 31473
rect 37369 31433 37381 31467
rect 37415 31464 37427 31467
rect 37458 31464 37464 31476
rect 37415 31436 37464 31464
rect 37415 31433 37427 31436
rect 37369 31427 37427 31433
rect 37458 31424 37464 31436
rect 37516 31424 37522 31476
rect 2133 31399 2191 31405
rect 2133 31365 2145 31399
rect 2179 31396 2191 31399
rect 2866 31396 2872 31408
rect 2179 31368 2872 31396
rect 2179 31365 2191 31368
rect 2133 31359 2191 31365
rect 2866 31356 2872 31368
rect 2924 31356 2930 31408
rect 15933 31399 15991 31405
rect 15933 31396 15945 31399
rect 15134 31368 15945 31396
rect 15933 31365 15945 31368
rect 15979 31365 15991 31399
rect 15933 31359 15991 31365
rect 20438 31356 20444 31408
rect 20496 31356 20502 31408
rect 21818 31356 21824 31408
rect 21876 31396 21882 31408
rect 23477 31399 23535 31405
rect 23477 31396 23489 31399
rect 21876 31368 23489 31396
rect 21876 31356 21882 31368
rect 23477 31365 23489 31368
rect 23523 31365 23535 31399
rect 24486 31396 24492 31408
rect 24447 31368 24492 31396
rect 23477 31359 23535 31365
rect 24486 31356 24492 31368
rect 24544 31356 24550 31408
rect 25958 31356 25964 31408
rect 26016 31396 26022 31408
rect 26602 31396 26608 31408
rect 26016 31368 26608 31396
rect 26016 31356 26022 31368
rect 26602 31356 26608 31368
rect 26660 31356 26666 31408
rect 27893 31399 27951 31405
rect 27893 31365 27905 31399
rect 27939 31396 27951 31399
rect 28442 31396 28448 31408
rect 27939 31368 28448 31396
rect 27939 31365 27951 31368
rect 27893 31359 27951 31365
rect 28442 31356 28448 31368
rect 28500 31356 28506 31408
rect 29178 31356 29184 31408
rect 29236 31396 29242 31408
rect 29362 31396 29368 31408
rect 29236 31368 29368 31396
rect 29236 31356 29242 31368
rect 29362 31356 29368 31368
rect 29420 31396 29426 31408
rect 30101 31399 30159 31405
rect 30101 31396 30113 31399
rect 29420 31368 30113 31396
rect 29420 31356 29426 31368
rect 30101 31365 30113 31368
rect 30147 31365 30159 31399
rect 30101 31359 30159 31365
rect 30317 31399 30375 31405
rect 30317 31365 30329 31399
rect 30363 31396 30375 31399
rect 30558 31396 30564 31408
rect 30363 31368 30564 31396
rect 30363 31365 30375 31368
rect 30317 31359 30375 31365
rect 30558 31356 30564 31368
rect 30616 31356 30622 31408
rect 33686 31396 33692 31408
rect 33152 31368 33692 31396
rect 1946 31328 1952 31340
rect 1907 31300 1952 31328
rect 1946 31288 1952 31300
rect 2004 31288 2010 31340
rect 9674 31328 9680 31340
rect 9635 31300 9680 31328
rect 9674 31288 9680 31300
rect 9732 31288 9738 31340
rect 10962 31288 10968 31340
rect 11020 31328 11026 31340
rect 11517 31331 11575 31337
rect 11517 31328 11529 31331
rect 11020 31300 11529 31328
rect 11020 31288 11026 31300
rect 11517 31297 11529 31300
rect 11563 31297 11575 31331
rect 11517 31291 11575 31297
rect 15562 31288 15568 31340
rect 15620 31328 15626 31340
rect 15841 31331 15899 31337
rect 15841 31328 15853 31331
rect 15620 31300 15853 31328
rect 15620 31288 15626 31300
rect 15841 31297 15853 31300
rect 15887 31328 15899 31331
rect 16761 31331 16819 31337
rect 16761 31328 16773 31331
rect 15887 31300 16773 31328
rect 15887 31297 15899 31300
rect 15841 31291 15899 31297
rect 16761 31297 16773 31300
rect 16807 31297 16819 31331
rect 16761 31291 16819 31297
rect 23293 31331 23351 31337
rect 23293 31297 23305 31331
rect 23339 31297 23351 31331
rect 26418 31328 26424 31340
rect 25622 31300 26424 31328
rect 23293 31291 23351 31297
rect 2958 31260 2964 31272
rect 2919 31232 2964 31260
rect 2958 31220 2964 31232
rect 3016 31220 3022 31272
rect 13633 31263 13691 31269
rect 13633 31229 13645 31263
rect 13679 31229 13691 31263
rect 13906 31260 13912 31272
rect 13867 31232 13912 31260
rect 13633 31223 13691 31229
rect 13648 31124 13676 31223
rect 13906 31220 13912 31232
rect 13964 31220 13970 31272
rect 19150 31260 19156 31272
rect 19111 31232 19156 31260
rect 19150 31220 19156 31232
rect 19208 31220 19214 31272
rect 19429 31263 19487 31269
rect 19429 31229 19441 31263
rect 19475 31260 19487 31263
rect 20714 31260 20720 31272
rect 19475 31232 20720 31260
rect 19475 31229 19487 31232
rect 19429 31223 19487 31229
rect 20714 31220 20720 31232
rect 20772 31220 20778 31272
rect 22002 31260 22008 31272
rect 21963 31232 22008 31260
rect 22002 31220 22008 31232
rect 22060 31220 22066 31272
rect 22281 31263 22339 31269
rect 22281 31229 22293 31263
rect 22327 31260 22339 31263
rect 22370 31260 22376 31272
rect 22327 31232 22376 31260
rect 22327 31229 22339 31232
rect 22281 31223 22339 31229
rect 22370 31220 22376 31232
rect 22428 31260 22434 31272
rect 22554 31260 22560 31272
rect 22428 31232 22560 31260
rect 22428 31220 22434 31232
rect 22554 31220 22560 31232
rect 22612 31260 22618 31272
rect 23308 31260 23336 31291
rect 26418 31288 26424 31300
rect 26476 31288 26482 31340
rect 27709 31331 27767 31337
rect 27709 31297 27721 31331
rect 27755 31297 27767 31331
rect 27709 31291 27767 31297
rect 24210 31260 24216 31272
rect 22612 31232 23336 31260
rect 24171 31232 24216 31260
rect 22612 31220 22618 31232
rect 24210 31220 24216 31232
rect 24268 31220 24274 31272
rect 24486 31220 24492 31272
rect 24544 31260 24550 31272
rect 27724 31260 27752 31291
rect 31110 31288 31116 31340
rect 31168 31328 31174 31340
rect 31386 31328 31392 31340
rect 31168 31300 31392 31328
rect 31168 31288 31174 31300
rect 31386 31288 31392 31300
rect 31444 31328 31450 31340
rect 33152 31328 33180 31368
rect 33686 31356 33692 31368
rect 33744 31356 33750 31408
rect 34790 31396 34796 31408
rect 34638 31368 34796 31396
rect 34790 31356 34796 31368
rect 34848 31356 34854 31408
rect 34900 31368 37320 31396
rect 31444 31300 33180 31328
rect 31444 31288 31450 31300
rect 33152 31272 33180 31300
rect 34698 31288 34704 31340
rect 34756 31328 34762 31340
rect 34900 31328 34928 31368
rect 34756 31300 34928 31328
rect 34756 31288 34762 31300
rect 36170 31288 36176 31340
rect 36228 31328 36234 31340
rect 36357 31331 36415 31337
rect 36357 31328 36369 31331
rect 36228 31300 36369 31328
rect 36228 31288 36234 31300
rect 36357 31297 36369 31300
rect 36403 31328 36415 31331
rect 36630 31328 36636 31340
rect 36403 31300 36636 31328
rect 36403 31297 36415 31300
rect 36357 31291 36415 31297
rect 36630 31288 36636 31300
rect 36688 31288 36694 31340
rect 37292 31337 37320 31368
rect 37550 31356 37556 31408
rect 37608 31396 37614 31408
rect 46017 31399 46075 31405
rect 46017 31396 46029 31399
rect 37608 31368 46029 31396
rect 37608 31356 37614 31368
rect 46017 31365 46029 31368
rect 46063 31365 46075 31399
rect 46017 31359 46075 31365
rect 46106 31356 46112 31408
rect 46164 31396 46170 31408
rect 47029 31399 47087 31405
rect 46164 31368 46209 31396
rect 46164 31356 46170 31368
rect 47029 31365 47041 31399
rect 47075 31396 47087 31399
rect 47394 31396 47400 31408
rect 47075 31368 47400 31396
rect 47075 31365 47087 31368
rect 47029 31359 47087 31365
rect 37277 31331 37335 31337
rect 37277 31297 37289 31331
rect 37323 31297 37335 31331
rect 37277 31291 37335 31297
rect 27890 31260 27896 31272
rect 24544 31232 27896 31260
rect 24544 31220 24550 31232
rect 27890 31220 27896 31232
rect 27948 31220 27954 31272
rect 33134 31260 33140 31272
rect 33095 31232 33140 31260
rect 33134 31220 33140 31232
rect 33192 31220 33198 31272
rect 33410 31260 33416 31272
rect 33371 31232 33416 31260
rect 33410 31220 33416 31232
rect 33468 31220 33474 31272
rect 36265 31263 36323 31269
rect 36265 31260 36277 31263
rect 34440 31232 36277 31260
rect 14642 31124 14648 31136
rect 13648 31096 14648 31124
rect 14642 31084 14648 31096
rect 14700 31084 14706 31136
rect 16758 31084 16764 31136
rect 16816 31124 16822 31136
rect 16853 31127 16911 31133
rect 16853 31124 16865 31127
rect 16816 31096 16865 31124
rect 16816 31084 16822 31096
rect 16853 31093 16865 31096
rect 16899 31093 16911 31127
rect 20898 31124 20904 31136
rect 20811 31096 20904 31124
rect 16853 31087 16911 31093
rect 20898 31084 20904 31096
rect 20956 31124 20962 31136
rect 21818 31124 21824 31136
rect 20956 31096 21824 31124
rect 20956 31084 20962 31096
rect 21818 31084 21824 31096
rect 21876 31084 21882 31136
rect 22462 31084 22468 31136
rect 22520 31124 22526 31136
rect 23661 31127 23719 31133
rect 23661 31124 23673 31127
rect 22520 31096 23673 31124
rect 22520 31084 22526 31096
rect 23661 31093 23673 31096
rect 23707 31093 23719 31127
rect 23661 31087 23719 31093
rect 25774 31084 25780 31136
rect 25832 31124 25838 31136
rect 25961 31127 26019 31133
rect 25961 31124 25973 31127
rect 25832 31096 25973 31124
rect 25832 31084 25838 31096
rect 25961 31093 25973 31096
rect 26007 31093 26019 31127
rect 25961 31087 26019 31093
rect 29086 31084 29092 31136
rect 29144 31124 29150 31136
rect 30285 31127 30343 31133
rect 30285 31124 30297 31127
rect 29144 31096 30297 31124
rect 29144 31084 29150 31096
rect 30285 31093 30297 31096
rect 30331 31093 30343 31127
rect 30285 31087 30343 31093
rect 30469 31127 30527 31133
rect 30469 31093 30481 31127
rect 30515 31124 30527 31127
rect 34440 31124 34468 31232
rect 36265 31229 36277 31232
rect 36311 31229 36323 31263
rect 36265 31223 36323 31229
rect 36725 31263 36783 31269
rect 36725 31229 36737 31263
rect 36771 31260 36783 31263
rect 37734 31260 37740 31272
rect 36771 31232 37740 31260
rect 36771 31229 36783 31232
rect 36725 31223 36783 31229
rect 37734 31220 37740 31232
rect 37792 31220 37798 31272
rect 44174 31220 44180 31272
rect 44232 31260 44238 31272
rect 47044 31260 47072 31359
rect 47394 31356 47400 31368
rect 47452 31356 47458 31408
rect 44232 31232 47072 31260
rect 44232 31220 44238 31232
rect 30515 31096 34468 31124
rect 30515 31093 30527 31096
rect 30469 31087 30527 31093
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 15194 30920 15200 30932
rect 15155 30892 15200 30920
rect 15194 30880 15200 30892
rect 15252 30880 15258 30932
rect 20714 30880 20720 30932
rect 20772 30920 20778 30932
rect 22097 30923 22155 30929
rect 22097 30920 22109 30923
rect 20772 30892 22109 30920
rect 20772 30880 20778 30892
rect 22097 30889 22109 30892
rect 22143 30889 22155 30923
rect 22097 30883 22155 30889
rect 22462 30880 22468 30932
rect 22520 30920 22526 30932
rect 22925 30923 22983 30929
rect 22925 30920 22937 30923
rect 22520 30892 22937 30920
rect 22520 30880 22526 30892
rect 22925 30889 22937 30892
rect 22971 30889 22983 30923
rect 22925 30883 22983 30889
rect 25682 30880 25688 30932
rect 25740 30920 25746 30932
rect 25777 30923 25835 30929
rect 25777 30920 25789 30923
rect 25740 30892 25789 30920
rect 25740 30880 25746 30892
rect 25777 30889 25789 30892
rect 25823 30889 25835 30923
rect 26418 30920 26424 30932
rect 26379 30892 26424 30920
rect 25777 30883 25835 30889
rect 26418 30880 26424 30892
rect 26476 30880 26482 30932
rect 12894 30812 12900 30864
rect 12952 30852 12958 30864
rect 14090 30852 14096 30864
rect 12952 30824 13952 30852
rect 14051 30824 14096 30852
rect 12952 30812 12958 30824
rect 12529 30787 12587 30793
rect 12529 30753 12541 30787
rect 12575 30784 12587 30787
rect 13262 30784 13268 30796
rect 12575 30756 13268 30784
rect 12575 30753 12587 30756
rect 12529 30747 12587 30753
rect 13262 30744 13268 30756
rect 13320 30744 13326 30796
rect 13924 30784 13952 30824
rect 14090 30812 14096 30824
rect 14148 30812 14154 30864
rect 13924 30756 15148 30784
rect 10962 30716 10968 30728
rect 10923 30688 10968 30716
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 11698 30716 11704 30728
rect 11659 30688 11704 30716
rect 11698 30676 11704 30688
rect 11756 30676 11762 30728
rect 11885 30719 11943 30725
rect 11885 30685 11897 30719
rect 11931 30716 11943 30719
rect 13078 30716 13084 30728
rect 11931 30688 13084 30716
rect 11931 30685 11943 30688
rect 11885 30679 11943 30685
rect 13078 30676 13084 30688
rect 13136 30676 13142 30728
rect 13722 30716 13728 30728
rect 13188 30688 13728 30716
rect 11054 30648 11060 30660
rect 11015 30620 11060 30648
rect 11054 30608 11060 30620
rect 11112 30608 11118 30660
rect 12710 30648 12716 30660
rect 12623 30620 12716 30648
rect 12710 30608 12716 30620
rect 12768 30648 12774 30660
rect 13188 30648 13216 30688
rect 13722 30676 13728 30688
rect 13780 30716 13786 30728
rect 15120 30725 15148 30756
rect 15378 30744 15384 30796
rect 15436 30784 15442 30796
rect 16025 30787 16083 30793
rect 16025 30784 16037 30787
rect 15436 30756 16037 30784
rect 15436 30744 15442 30756
rect 16025 30753 16037 30756
rect 16071 30753 16083 30787
rect 16025 30747 16083 30753
rect 19150 30744 19156 30796
rect 19208 30784 19214 30796
rect 19245 30787 19303 30793
rect 19245 30784 19257 30787
rect 19208 30756 19257 30784
rect 19208 30744 19214 30756
rect 19245 30753 19257 30756
rect 19291 30784 19303 30787
rect 24210 30784 24216 30796
rect 19291 30756 24216 30784
rect 19291 30753 19303 30756
rect 19245 30747 19303 30753
rect 24210 30744 24216 30756
rect 24268 30744 24274 30796
rect 25593 30787 25651 30793
rect 25593 30753 25605 30787
rect 25639 30784 25651 30787
rect 25682 30784 25688 30796
rect 25639 30756 25688 30784
rect 25639 30753 25651 30756
rect 25593 30747 25651 30753
rect 25682 30744 25688 30756
rect 25740 30784 25746 30796
rect 26050 30784 26056 30796
rect 25740 30756 26056 30784
rect 25740 30744 25746 30756
rect 26050 30744 26056 30756
rect 26108 30744 26114 30796
rect 14369 30719 14427 30725
rect 14369 30716 14381 30719
rect 13780 30688 14381 30716
rect 13780 30676 13786 30688
rect 14369 30685 14381 30688
rect 14415 30685 14427 30719
rect 14369 30679 14427 30685
rect 15105 30719 15163 30725
rect 15105 30685 15117 30719
rect 15151 30685 15163 30719
rect 15105 30679 15163 30685
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30685 15347 30719
rect 15746 30716 15752 30728
rect 15707 30688 15752 30716
rect 15289 30679 15347 30685
rect 12768 30620 13216 30648
rect 12768 30608 12774 30620
rect 13538 30608 13544 30660
rect 13596 30648 13602 30660
rect 14461 30651 14519 30657
rect 14461 30648 14473 30651
rect 13596 30620 14473 30648
rect 13596 30608 13602 30620
rect 14461 30617 14473 30620
rect 14507 30617 14519 30651
rect 15304 30648 15332 30679
rect 15746 30676 15752 30688
rect 15804 30676 15810 30728
rect 21818 30716 21824 30728
rect 21779 30688 21824 30716
rect 21818 30676 21824 30688
rect 21876 30676 21882 30728
rect 21910 30676 21916 30728
rect 21968 30716 21974 30728
rect 21968 30688 22013 30716
rect 21968 30676 21974 30688
rect 22370 30676 22376 30728
rect 22428 30716 22434 30728
rect 22741 30719 22799 30725
rect 22741 30716 22753 30719
rect 22428 30688 22753 30716
rect 22428 30676 22434 30688
rect 22741 30685 22753 30688
rect 22787 30685 22799 30719
rect 22741 30679 22799 30685
rect 23017 30719 23075 30725
rect 23017 30685 23029 30719
rect 23063 30685 23075 30719
rect 23017 30679 23075 30685
rect 25501 30719 25559 30725
rect 25501 30685 25513 30719
rect 25547 30716 25559 30719
rect 25774 30716 25780 30728
rect 25547 30688 25780 30716
rect 25547 30685 25559 30688
rect 25501 30679 25559 30685
rect 14461 30611 14519 30617
rect 14752 30620 15332 30648
rect 14752 30592 14780 30620
rect 16758 30608 16764 30660
rect 16816 30608 16822 30660
rect 19521 30651 19579 30657
rect 19521 30617 19533 30651
rect 19567 30617 19579 30651
rect 20806 30648 20812 30660
rect 20746 30620 20812 30648
rect 19521 30611 19579 30617
rect 11790 30580 11796 30592
rect 11751 30552 11796 30580
rect 11790 30540 11796 30552
rect 11848 30540 11854 30592
rect 12526 30540 12532 30592
rect 12584 30580 12590 30592
rect 12805 30583 12863 30589
rect 12805 30580 12817 30583
rect 12584 30552 12817 30580
rect 12584 30540 12590 30552
rect 12805 30549 12817 30552
rect 12851 30549 12863 30583
rect 12805 30543 12863 30549
rect 12894 30540 12900 30592
rect 12952 30580 12958 30592
rect 12952 30552 12997 30580
rect 12952 30540 12958 30552
rect 13078 30540 13084 30592
rect 13136 30580 13142 30592
rect 13136 30552 13181 30580
rect 13136 30540 13142 30552
rect 13262 30540 13268 30592
rect 13320 30580 13326 30592
rect 14277 30583 14335 30589
rect 14277 30580 14289 30583
rect 13320 30552 14289 30580
rect 13320 30540 13326 30552
rect 14277 30549 14289 30552
rect 14323 30549 14335 30583
rect 14277 30543 14335 30549
rect 14645 30583 14703 30589
rect 14645 30549 14657 30583
rect 14691 30580 14703 30583
rect 14734 30580 14740 30592
rect 14691 30552 14740 30580
rect 14691 30549 14703 30552
rect 14645 30543 14703 30549
rect 14734 30540 14740 30552
rect 14792 30540 14798 30592
rect 16666 30540 16672 30592
rect 16724 30580 16730 30592
rect 17494 30580 17500 30592
rect 16724 30552 17500 30580
rect 16724 30540 16730 30552
rect 17494 30540 17500 30552
rect 17552 30540 17558 30592
rect 19536 30580 19564 30611
rect 20806 30608 20812 30620
rect 20864 30608 20870 30660
rect 21082 30648 21088 30660
rect 20916 30620 21088 30648
rect 20916 30580 20944 30620
rect 21082 30608 21088 30620
rect 21140 30608 21146 30660
rect 21726 30608 21732 30660
rect 21784 30648 21790 30660
rect 23032 30648 23060 30679
rect 25774 30676 25780 30688
rect 25832 30676 25838 30728
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30716 26387 30719
rect 28261 30719 28319 30725
rect 28261 30716 28273 30719
rect 26375 30688 28273 30716
rect 26375 30685 26387 30688
rect 26329 30679 26387 30685
rect 28261 30685 28273 30688
rect 28307 30716 28319 30719
rect 28626 30716 28632 30728
rect 28307 30688 28632 30716
rect 28307 30685 28319 30688
rect 28261 30679 28319 30685
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 30190 30676 30196 30728
rect 30248 30716 30254 30728
rect 33226 30716 33232 30728
rect 30248 30688 33232 30716
rect 30248 30676 30254 30688
rect 33226 30676 33232 30688
rect 33284 30716 33290 30728
rect 33413 30719 33471 30725
rect 33413 30716 33425 30719
rect 33284 30688 33425 30716
rect 33284 30676 33290 30688
rect 33413 30685 33425 30688
rect 33459 30685 33471 30719
rect 33413 30679 33471 30685
rect 21784 30620 23060 30648
rect 24673 30651 24731 30657
rect 21784 30608 21790 30620
rect 24673 30617 24685 30651
rect 24719 30648 24731 30651
rect 24854 30648 24860 30660
rect 24719 30620 24860 30648
rect 24719 30617 24731 30620
rect 24673 30611 24731 30617
rect 24854 30608 24860 30620
rect 24912 30608 24918 30660
rect 31294 30648 31300 30660
rect 31255 30620 31300 30648
rect 31294 30608 31300 30620
rect 31352 30608 31358 30660
rect 33597 30651 33655 30657
rect 33597 30617 33609 30651
rect 33643 30648 33655 30651
rect 33686 30648 33692 30660
rect 33643 30620 33692 30648
rect 33643 30617 33655 30620
rect 33597 30611 33655 30617
rect 33686 30608 33692 30620
rect 33744 30608 33750 30660
rect 19536 30552 20944 30580
rect 20990 30540 20996 30592
rect 21048 30580 21054 30592
rect 21450 30580 21456 30592
rect 21048 30552 21093 30580
rect 21411 30552 21456 30580
rect 21048 30540 21054 30552
rect 21450 30540 21456 30552
rect 21508 30540 21514 30592
rect 22557 30583 22615 30589
rect 22557 30549 22569 30583
rect 22603 30580 22615 30583
rect 22646 30580 22652 30592
rect 22603 30552 22652 30580
rect 22603 30549 22615 30552
rect 22557 30543 22615 30549
rect 22646 30540 22652 30552
rect 22704 30540 22710 30592
rect 24210 30540 24216 30592
rect 24268 30580 24274 30592
rect 24765 30583 24823 30589
rect 24765 30580 24777 30583
rect 24268 30552 24777 30580
rect 24268 30540 24274 30552
rect 24765 30549 24777 30552
rect 24811 30580 24823 30583
rect 25038 30580 25044 30592
rect 24811 30552 25044 30580
rect 24811 30549 24823 30552
rect 24765 30543 24823 30549
rect 25038 30540 25044 30552
rect 25096 30540 25102 30592
rect 28350 30580 28356 30592
rect 28311 30552 28356 30580
rect 28350 30540 28356 30552
rect 28408 30540 28414 30592
rect 30374 30540 30380 30592
rect 30432 30580 30438 30592
rect 31386 30580 31392 30592
rect 30432 30552 31392 30580
rect 30432 30540 30438 30552
rect 31386 30540 31392 30552
rect 31444 30540 31450 30592
rect 33318 30540 33324 30592
rect 33376 30580 33382 30592
rect 33781 30583 33839 30589
rect 33781 30580 33793 30583
rect 33376 30552 33793 30580
rect 33376 30540 33382 30552
rect 33781 30549 33793 30552
rect 33827 30549 33839 30583
rect 33781 30543 33839 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 13262 30376 13268 30388
rect 13223 30348 13268 30376
rect 13262 30336 13268 30348
rect 13320 30336 13326 30388
rect 13817 30379 13875 30385
rect 13817 30345 13829 30379
rect 13863 30376 13875 30379
rect 13906 30376 13912 30388
rect 13863 30348 13912 30376
rect 13863 30345 13875 30348
rect 13817 30339 13875 30345
rect 13906 30336 13912 30348
rect 13964 30336 13970 30388
rect 15746 30336 15752 30388
rect 15804 30376 15810 30388
rect 15841 30379 15899 30385
rect 15841 30376 15853 30379
rect 15804 30348 15853 30376
rect 15804 30336 15810 30348
rect 15841 30345 15853 30348
rect 15887 30345 15899 30379
rect 24486 30376 24492 30388
rect 24447 30348 24492 30376
rect 15841 30339 15899 30345
rect 24486 30336 24492 30348
rect 24544 30336 24550 30388
rect 25314 30336 25320 30388
rect 25372 30376 25378 30388
rect 46842 30376 46848 30388
rect 25372 30348 46848 30376
rect 25372 30336 25378 30348
rect 46842 30336 46848 30348
rect 46900 30336 46906 30388
rect 11790 30308 11796 30320
rect 11751 30280 11796 30308
rect 11790 30268 11796 30280
rect 11848 30268 11854 30320
rect 12434 30268 12440 30320
rect 12492 30268 12498 30320
rect 14642 30268 14648 30320
rect 14700 30308 14706 30320
rect 14829 30311 14887 30317
rect 14829 30308 14841 30311
rect 14700 30280 14841 30308
rect 14700 30268 14706 30280
rect 14829 30277 14841 30280
rect 14875 30277 14887 30311
rect 14829 30271 14887 30277
rect 21082 30268 21088 30320
rect 21140 30308 21146 30320
rect 22833 30311 22891 30317
rect 22833 30308 22845 30311
rect 21140 30280 22845 30308
rect 21140 30268 21146 30280
rect 22833 30277 22845 30280
rect 22879 30277 22891 30311
rect 26418 30308 26424 30320
rect 22833 30271 22891 30277
rect 24504 30280 26424 30308
rect 11054 30200 11060 30252
rect 11112 30240 11118 30252
rect 11517 30243 11575 30249
rect 11517 30240 11529 30243
rect 11112 30212 11529 30240
rect 11112 30200 11118 30212
rect 11517 30209 11529 30212
rect 11563 30209 11575 30243
rect 11517 30203 11575 30209
rect 14001 30243 14059 30249
rect 14001 30209 14013 30243
rect 14047 30240 14059 30243
rect 14737 30243 14795 30249
rect 14047 30212 14688 30240
rect 14047 30209 14059 30212
rect 14001 30203 14059 30209
rect 13078 30132 13084 30184
rect 13136 30172 13142 30184
rect 14185 30175 14243 30181
rect 14185 30172 14197 30175
rect 13136 30144 14197 30172
rect 13136 30132 13142 30144
rect 14185 30141 14197 30144
rect 14231 30141 14243 30175
rect 14185 30135 14243 30141
rect 14277 30175 14335 30181
rect 14277 30141 14289 30175
rect 14323 30141 14335 30175
rect 14660 30172 14688 30212
rect 14737 30209 14749 30243
rect 14783 30240 14795 30243
rect 15841 30243 15899 30249
rect 15841 30240 15853 30243
rect 14783 30212 15853 30240
rect 14783 30209 14795 30212
rect 14737 30203 14795 30209
rect 15841 30209 15853 30212
rect 15887 30240 15899 30243
rect 16114 30240 16120 30252
rect 15887 30212 16120 30240
rect 15887 30209 15899 30212
rect 15841 30203 15899 30209
rect 16114 30200 16120 30212
rect 16172 30200 16178 30252
rect 20898 30240 20904 30252
rect 20859 30212 20904 30240
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 22152 30212 22197 30240
rect 22152 30200 22158 30212
rect 22278 30200 22284 30252
rect 22336 30240 22342 30252
rect 22649 30243 22707 30249
rect 22336 30212 22381 30240
rect 22336 30200 22342 30212
rect 22649 30209 22661 30243
rect 22695 30240 22707 30243
rect 22738 30240 22744 30252
rect 22695 30212 22744 30240
rect 22695 30209 22707 30212
rect 22649 30203 22707 30209
rect 22738 30200 22744 30212
rect 22796 30200 22802 30252
rect 23014 30200 23020 30252
rect 23072 30240 23078 30252
rect 24504 30249 24532 30280
rect 26418 30268 26424 30280
rect 26476 30268 26482 30320
rect 28350 30268 28356 30320
rect 28408 30268 28414 30320
rect 30374 30308 30380 30320
rect 29840 30280 30380 30308
rect 24486 30243 24544 30249
rect 24486 30240 24498 30243
rect 23072 30212 24498 30240
rect 23072 30200 23078 30212
rect 24486 30209 24498 30212
rect 24532 30209 24544 30243
rect 24486 30203 24544 30209
rect 25038 30200 25044 30252
rect 25096 30240 25102 30252
rect 29840 30249 29868 30280
rect 30374 30268 30380 30280
rect 30432 30268 30438 30320
rect 33134 30268 33140 30320
rect 33192 30308 33198 30320
rect 33192 30280 34560 30308
rect 33192 30268 33198 30280
rect 27341 30243 27399 30249
rect 27341 30240 27353 30243
rect 25096 30212 27353 30240
rect 25096 30200 25102 30212
rect 27341 30209 27353 30212
rect 27387 30209 27399 30243
rect 27341 30203 27399 30209
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 32490 30240 32496 30252
rect 31234 30212 32496 30240
rect 29825 30203 29883 30209
rect 32490 30200 32496 30212
rect 32548 30200 32554 30252
rect 33318 30240 33324 30252
rect 33279 30212 33324 30240
rect 33318 30200 33324 30212
rect 33376 30200 33382 30252
rect 33502 30240 33508 30252
rect 33463 30212 33508 30240
rect 33502 30200 33508 30212
rect 33560 30200 33566 30252
rect 33870 30240 33876 30252
rect 33831 30212 33876 30240
rect 33870 30200 33876 30212
rect 33928 30200 33934 30252
rect 34532 30249 34560 30280
rect 35342 30268 35348 30320
rect 35400 30268 35406 30320
rect 34517 30243 34575 30249
rect 34517 30209 34529 30243
rect 34563 30209 34575 30243
rect 34517 30203 34575 30209
rect 15194 30172 15200 30184
rect 14660 30144 15200 30172
rect 14277 30135 14335 30141
rect 14090 30064 14096 30116
rect 14148 30104 14154 30116
rect 14292 30104 14320 30135
rect 15194 30132 15200 30144
rect 15252 30132 15258 30184
rect 20990 30172 20996 30184
rect 20903 30144 20996 30172
rect 20990 30132 20996 30144
rect 21048 30172 21054 30184
rect 22370 30172 22376 30184
rect 21048 30144 22376 30172
rect 21048 30132 21054 30144
rect 22370 30132 22376 30144
rect 22428 30132 22434 30184
rect 22465 30175 22523 30181
rect 22465 30141 22477 30175
rect 22511 30172 22523 30175
rect 23382 30172 23388 30184
rect 22511 30144 23388 30172
rect 22511 30141 22523 30144
rect 22465 30135 22523 30141
rect 23382 30132 23388 30144
rect 23440 30132 23446 30184
rect 24946 30172 24952 30184
rect 24907 30144 24952 30172
rect 24946 30132 24952 30144
rect 25004 30132 25010 30184
rect 27614 30172 27620 30184
rect 27575 30144 27620 30172
rect 27614 30132 27620 30144
rect 27672 30132 27678 30184
rect 30101 30175 30159 30181
rect 30101 30141 30113 30175
rect 30147 30172 30159 30175
rect 30650 30172 30656 30184
rect 30147 30144 30656 30172
rect 30147 30141 30159 30144
rect 30101 30135 30159 30141
rect 30650 30132 30656 30144
rect 30708 30132 30714 30184
rect 31110 30132 31116 30184
rect 31168 30172 31174 30184
rect 33226 30172 33232 30184
rect 31168 30144 33232 30172
rect 31168 30132 31174 30144
rect 33226 30132 33232 30144
rect 33284 30132 33290 30184
rect 33594 30172 33600 30184
rect 33555 30144 33600 30172
rect 33594 30132 33600 30144
rect 33652 30132 33658 30184
rect 33689 30175 33747 30181
rect 33689 30141 33701 30175
rect 33735 30141 33747 30175
rect 33689 30135 33747 30141
rect 34057 30175 34115 30181
rect 34057 30141 34069 30175
rect 34103 30172 34115 30175
rect 34793 30175 34851 30181
rect 34793 30172 34805 30175
rect 34103 30144 34805 30172
rect 34103 30141 34115 30144
rect 34057 30135 34115 30141
rect 34793 30141 34805 30144
rect 34839 30141 34851 30175
rect 34793 30135 34851 30141
rect 21726 30104 21732 30116
rect 14148 30076 14320 30104
rect 21100 30076 21732 30104
rect 14148 30064 14154 30076
rect 21100 30045 21128 30076
rect 21726 30064 21732 30076
rect 21784 30064 21790 30116
rect 24302 30104 24308 30116
rect 24263 30076 24308 30104
rect 24302 30064 24308 30076
rect 24360 30064 24366 30116
rect 24857 30107 24915 30113
rect 24857 30073 24869 30107
rect 24903 30104 24915 30107
rect 26234 30104 26240 30116
rect 24903 30076 26240 30104
rect 24903 30073 24915 30076
rect 24857 30067 24915 30073
rect 26234 30064 26240 30076
rect 26292 30064 26298 30116
rect 28626 30064 28632 30116
rect 28684 30104 28690 30116
rect 32398 30104 32404 30116
rect 28684 30076 29960 30104
rect 28684 30064 28690 30076
rect 21085 30039 21143 30045
rect 21085 30005 21097 30039
rect 21131 30005 21143 30039
rect 21266 30036 21272 30048
rect 21227 30008 21272 30036
rect 21085 29999 21143 30005
rect 21266 29996 21272 30008
rect 21324 29996 21330 30048
rect 24762 29996 24768 30048
rect 24820 30036 24826 30048
rect 27062 30036 27068 30048
rect 24820 30008 27068 30036
rect 24820 29996 24826 30008
rect 27062 29996 27068 30008
rect 27120 29996 27126 30048
rect 27338 29996 27344 30048
rect 27396 30036 27402 30048
rect 28644 30036 28672 30064
rect 29086 30036 29092 30048
rect 27396 30008 28672 30036
rect 29047 30008 29092 30036
rect 27396 29996 27402 30008
rect 29086 29996 29092 30008
rect 29144 29996 29150 30048
rect 29932 30036 29960 30076
rect 31404 30076 32404 30104
rect 31404 30036 31432 30076
rect 32398 30064 32404 30076
rect 32456 30064 32462 30116
rect 31570 30036 31576 30048
rect 29932 30008 31432 30036
rect 31531 30008 31576 30036
rect 31570 29996 31576 30008
rect 31628 29996 31634 30048
rect 33704 30036 33732 30135
rect 44450 30104 44456 30116
rect 36188 30076 44456 30104
rect 36188 30036 36216 30076
rect 44450 30064 44456 30076
rect 44508 30064 44514 30116
rect 33704 30008 36216 30036
rect 36262 29996 36268 30048
rect 36320 30036 36326 30048
rect 36320 30008 36365 30036
rect 36320 29996 36326 30008
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 11698 29792 11704 29844
rect 11756 29832 11762 29844
rect 11793 29835 11851 29841
rect 11793 29832 11805 29835
rect 11756 29804 11805 29832
rect 11756 29792 11762 29804
rect 11793 29801 11805 29804
rect 11839 29801 11851 29835
rect 11793 29795 11851 29801
rect 12434 29792 12440 29844
rect 12492 29832 12498 29844
rect 21450 29832 21456 29844
rect 12492 29804 12537 29832
rect 21411 29804 21456 29832
rect 12492 29792 12498 29804
rect 21450 29792 21456 29804
rect 21508 29792 21514 29844
rect 22005 29835 22063 29841
rect 22005 29801 22017 29835
rect 22051 29832 22063 29835
rect 22462 29832 22468 29844
rect 22051 29804 22468 29832
rect 22051 29801 22063 29804
rect 22005 29795 22063 29801
rect 22462 29792 22468 29804
rect 22520 29792 22526 29844
rect 22646 29832 22652 29844
rect 22607 29804 22652 29832
rect 22646 29792 22652 29804
rect 22704 29792 22710 29844
rect 24946 29792 24952 29844
rect 25004 29832 25010 29844
rect 26234 29832 26240 29844
rect 25004 29804 26240 29832
rect 25004 29792 25010 29804
rect 26234 29792 26240 29804
rect 26292 29792 26298 29844
rect 27614 29792 27620 29844
rect 27672 29832 27678 29844
rect 27801 29835 27859 29841
rect 27801 29832 27813 29835
rect 27672 29804 27813 29832
rect 27672 29792 27678 29804
rect 27801 29801 27813 29804
rect 27847 29801 27859 29835
rect 27801 29795 27859 29801
rect 28813 29835 28871 29841
rect 28813 29801 28825 29835
rect 28859 29801 28871 29835
rect 28813 29795 28871 29801
rect 22094 29724 22100 29776
rect 22152 29764 22158 29776
rect 23109 29767 23167 29773
rect 23109 29764 23121 29767
rect 22152 29736 23121 29764
rect 22152 29724 22158 29736
rect 23109 29733 23121 29736
rect 23155 29733 23167 29767
rect 23109 29727 23167 29733
rect 24302 29724 24308 29776
rect 24360 29764 24366 29776
rect 28828 29764 28856 29795
rect 28994 29792 29000 29844
rect 29052 29832 29058 29844
rect 30834 29832 30840 29844
rect 29052 29804 29097 29832
rect 30795 29804 30840 29832
rect 29052 29792 29058 29804
rect 30834 29792 30840 29804
rect 30892 29792 30898 29844
rect 31110 29792 31116 29844
rect 31168 29832 31174 29844
rect 31757 29835 31815 29841
rect 31757 29832 31769 29835
rect 31168 29804 31769 29832
rect 31168 29792 31174 29804
rect 31757 29801 31769 29804
rect 31803 29801 31815 29835
rect 32490 29832 32496 29844
rect 32451 29804 32496 29832
rect 31757 29795 31815 29801
rect 32490 29792 32496 29804
rect 32548 29792 32554 29844
rect 33594 29792 33600 29844
rect 33652 29832 33658 29844
rect 33781 29835 33839 29841
rect 33781 29832 33793 29835
rect 33652 29804 33793 29832
rect 33652 29792 33658 29804
rect 33781 29801 33793 29804
rect 33827 29801 33839 29835
rect 33781 29795 33839 29801
rect 35161 29835 35219 29841
rect 35161 29801 35173 29835
rect 35207 29832 35219 29835
rect 35342 29832 35348 29844
rect 35207 29804 35348 29832
rect 35207 29801 35219 29804
rect 35161 29795 35219 29801
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 36173 29835 36231 29841
rect 36173 29801 36185 29835
rect 36219 29832 36231 29835
rect 36446 29832 36452 29844
rect 36219 29804 36452 29832
rect 36219 29801 36231 29804
rect 36173 29795 36231 29801
rect 36446 29792 36452 29804
rect 36504 29792 36510 29844
rect 29086 29764 29092 29776
rect 24360 29736 28764 29764
rect 28828 29736 29092 29764
rect 24360 29724 24366 29736
rect 11609 29699 11667 29705
rect 11609 29665 11621 29699
rect 11655 29696 11667 29699
rect 12710 29696 12716 29708
rect 11655 29668 12716 29696
rect 11655 29665 11667 29668
rect 11609 29659 11667 29665
rect 12710 29656 12716 29668
rect 12768 29656 12774 29708
rect 16114 29696 16120 29708
rect 15672 29668 16120 29696
rect 11238 29588 11244 29640
rect 11296 29628 11302 29640
rect 11425 29631 11483 29637
rect 11425 29628 11437 29631
rect 11296 29600 11437 29628
rect 11296 29588 11302 29600
rect 11425 29597 11437 29600
rect 11471 29597 11483 29631
rect 11425 29591 11483 29597
rect 11793 29631 11851 29637
rect 11793 29597 11805 29631
rect 11839 29597 11851 29631
rect 11793 29591 11851 29597
rect 12345 29631 12403 29637
rect 12345 29597 12357 29631
rect 12391 29628 12403 29631
rect 12618 29628 12624 29640
rect 12391 29600 12624 29628
rect 12391 29597 12403 29600
rect 12345 29591 12403 29597
rect 9122 29520 9128 29572
rect 9180 29560 9186 29572
rect 11808 29560 11836 29591
rect 12618 29588 12624 29600
rect 12676 29628 12682 29640
rect 15562 29628 15568 29640
rect 12676 29600 15568 29628
rect 12676 29588 12682 29600
rect 15562 29588 15568 29600
rect 15620 29588 15626 29640
rect 15672 29637 15700 29668
rect 16114 29656 16120 29668
rect 16172 29656 16178 29708
rect 24946 29696 24952 29708
rect 22112 29668 24952 29696
rect 22112 29637 22140 29668
rect 24946 29656 24952 29668
rect 25004 29656 25010 29708
rect 25682 29696 25688 29708
rect 25643 29668 25688 29696
rect 25682 29656 25688 29668
rect 25740 29696 25746 29708
rect 26050 29696 26056 29708
rect 25740 29668 26056 29696
rect 25740 29656 25746 29668
rect 26050 29656 26056 29668
rect 26108 29656 26114 29708
rect 26605 29699 26663 29705
rect 26605 29665 26617 29699
rect 26651 29696 26663 29699
rect 28626 29696 28632 29708
rect 26651 29668 28632 29696
rect 26651 29665 26663 29668
rect 26605 29659 26663 29665
rect 28626 29656 28632 29668
rect 28684 29656 28690 29708
rect 28736 29696 28764 29736
rect 29086 29724 29092 29736
rect 29144 29764 29150 29776
rect 46842 29764 46848 29776
rect 29144 29736 29592 29764
rect 29144 29724 29150 29736
rect 29564 29705 29592 29736
rect 29656 29736 46848 29764
rect 29549 29699 29607 29705
rect 28736 29668 28948 29696
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29597 15715 29631
rect 15657 29591 15715 29597
rect 15749 29631 15807 29637
rect 15749 29597 15761 29631
rect 15795 29628 15807 29631
rect 16209 29631 16267 29637
rect 16209 29628 16221 29631
rect 15795 29600 16221 29628
rect 15795 29597 15807 29600
rect 15749 29591 15807 29597
rect 16209 29597 16221 29600
rect 16255 29597 16267 29631
rect 16209 29591 16267 29597
rect 21634 29631 21692 29637
rect 21634 29597 21646 29631
rect 21680 29597 21692 29631
rect 21634 29591 21692 29597
rect 22097 29631 22155 29637
rect 22097 29597 22109 29631
rect 22143 29597 22155 29631
rect 22097 29591 22155 29597
rect 13262 29560 13268 29572
rect 9180 29532 13268 29560
rect 9180 29520 9186 29532
rect 13262 29520 13268 29532
rect 13320 29520 13326 29572
rect 15930 29520 15936 29572
rect 15988 29560 15994 29572
rect 16485 29563 16543 29569
rect 16485 29560 16497 29563
rect 15988 29532 16497 29560
rect 15988 29520 15994 29532
rect 16485 29529 16497 29532
rect 16531 29529 16543 29563
rect 16485 29523 16543 29529
rect 17034 29520 17040 29572
rect 17092 29520 17098 29572
rect 21649 29560 21677 29591
rect 22186 29588 22192 29640
rect 22244 29628 22250 29640
rect 22557 29631 22615 29637
rect 22557 29628 22569 29631
rect 22244 29600 22569 29628
rect 22244 29588 22250 29600
rect 22557 29597 22569 29600
rect 22603 29597 22615 29631
rect 22557 29591 22615 29597
rect 22925 29631 22983 29637
rect 22925 29597 22937 29631
rect 22971 29628 22983 29631
rect 23106 29628 23112 29640
rect 22971 29600 23112 29628
rect 22971 29597 22983 29600
rect 22925 29591 22983 29597
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 25501 29631 25559 29637
rect 25501 29597 25513 29631
rect 25547 29597 25559 29631
rect 25774 29628 25780 29640
rect 25687 29600 25780 29628
rect 25501 29591 25559 29597
rect 23014 29560 23020 29572
rect 21649 29532 23020 29560
rect 23014 29520 23020 29532
rect 23072 29520 23078 29572
rect 24670 29520 24676 29572
rect 24728 29560 24734 29572
rect 25516 29560 25544 29591
rect 25774 29588 25780 29600
rect 25832 29628 25838 29640
rect 26237 29631 26295 29637
rect 26237 29628 26249 29631
rect 25832 29600 26249 29628
rect 25832 29588 25838 29600
rect 26237 29597 26249 29600
rect 26283 29597 26295 29631
rect 27154 29628 27160 29640
rect 27115 29600 27160 29628
rect 26237 29591 26295 29597
rect 27154 29588 27160 29600
rect 27212 29588 27218 29640
rect 27246 29588 27252 29640
rect 27304 29628 27310 29640
rect 27663 29631 27721 29637
rect 27304 29600 27349 29628
rect 27304 29588 27310 29600
rect 27663 29597 27675 29631
rect 27709 29628 27721 29631
rect 28258 29628 28264 29640
rect 27709 29600 28264 29628
rect 27709 29597 27721 29600
rect 27663 29591 27721 29597
rect 28258 29588 28264 29600
rect 28316 29588 28322 29640
rect 28810 29628 28816 29640
rect 28771 29600 28816 29628
rect 28810 29588 28816 29600
rect 28868 29588 28874 29640
rect 28920 29628 28948 29668
rect 29549 29665 29561 29699
rect 29595 29665 29607 29699
rect 29549 29659 29607 29665
rect 29656 29628 29684 29736
rect 46842 29724 46848 29736
rect 46900 29724 46906 29776
rect 30374 29656 30380 29708
rect 30432 29696 30438 29708
rect 30929 29699 30987 29705
rect 30929 29696 30941 29699
rect 30432 29668 30941 29696
rect 30432 29656 30438 29668
rect 30929 29665 30941 29668
rect 30975 29696 30987 29699
rect 31386 29696 31392 29708
rect 30975 29668 31392 29696
rect 30975 29665 30987 29668
rect 30929 29659 30987 29665
rect 31386 29656 31392 29668
rect 31444 29696 31450 29708
rect 31570 29696 31576 29708
rect 31444 29668 31576 29696
rect 31444 29656 31450 29668
rect 31570 29656 31576 29668
rect 31628 29696 31634 29708
rect 31941 29699 31999 29705
rect 31941 29696 31953 29699
rect 31628 29668 31953 29696
rect 31628 29656 31634 29668
rect 31941 29665 31953 29668
rect 31987 29665 31999 29699
rect 33505 29699 33563 29705
rect 33505 29696 33517 29699
rect 31941 29659 31999 29665
rect 33428 29668 33517 29696
rect 33428 29640 33456 29668
rect 33505 29665 33517 29668
rect 33551 29665 33563 29699
rect 34422 29696 34428 29708
rect 33505 29659 33563 29665
rect 33888 29668 34428 29696
rect 28920 29600 29684 29628
rect 30282 29588 30288 29640
rect 30340 29628 30346 29640
rect 30837 29631 30895 29637
rect 30837 29628 30849 29631
rect 30340 29600 30849 29628
rect 30340 29588 30346 29600
rect 30837 29597 30849 29600
rect 30883 29597 30895 29631
rect 30837 29591 30895 29597
rect 31018 29588 31024 29640
rect 31076 29628 31082 29640
rect 31665 29631 31723 29637
rect 31665 29628 31677 29631
rect 31076 29600 31677 29628
rect 31076 29588 31082 29600
rect 31665 29597 31677 29600
rect 31711 29597 31723 29631
rect 32398 29628 32404 29640
rect 32359 29600 32404 29628
rect 31665 29591 31723 29597
rect 32398 29588 32404 29600
rect 32456 29588 32462 29640
rect 33410 29588 33416 29640
rect 33468 29588 33474 29640
rect 33583 29631 33641 29637
rect 33583 29597 33595 29631
rect 33629 29622 33641 29631
rect 33686 29622 33692 29640
rect 33629 29597 33692 29622
rect 33583 29594 33692 29597
rect 33583 29591 33641 29594
rect 33686 29588 33692 29594
rect 33744 29628 33750 29640
rect 33888 29628 33916 29668
rect 34422 29656 34428 29668
rect 34480 29656 34486 29708
rect 36078 29696 36084 29708
rect 36039 29668 36084 29696
rect 36078 29656 36084 29668
rect 36136 29656 36142 29708
rect 33744 29600 33916 29628
rect 33744 29588 33750 29600
rect 33962 29588 33968 29640
rect 34020 29628 34026 29640
rect 35069 29631 35127 29637
rect 35069 29628 35081 29631
rect 34020 29600 35081 29628
rect 34020 29588 34026 29600
rect 35069 29597 35081 29600
rect 35115 29597 35127 29631
rect 36170 29628 36176 29640
rect 36131 29600 36176 29628
rect 35069 29591 35127 29597
rect 36170 29588 36176 29600
rect 36228 29588 36234 29640
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 47581 29631 47639 29637
rect 47581 29597 47593 29631
rect 47627 29628 47639 29631
rect 47762 29628 47768 29640
rect 47627 29600 47768 29628
rect 47627 29597 47639 29600
rect 47581 29591 47639 29597
rect 47762 29588 47768 29600
rect 47820 29588 47826 29640
rect 26142 29560 26148 29572
rect 24728 29532 26148 29560
rect 24728 29520 24734 29532
rect 26142 29520 26148 29532
rect 26200 29560 26206 29572
rect 26421 29563 26479 29569
rect 26421 29560 26433 29563
rect 26200 29532 26433 29560
rect 26200 29520 26206 29532
rect 26421 29529 26433 29532
rect 26467 29529 26479 29563
rect 26421 29523 26479 29529
rect 27062 29520 27068 29572
rect 27120 29560 27126 29572
rect 27433 29563 27491 29569
rect 27433 29560 27445 29563
rect 27120 29532 27445 29560
rect 27120 29520 27126 29532
rect 27433 29529 27445 29532
rect 27479 29529 27491 29563
rect 27433 29523 27491 29529
rect 27525 29563 27583 29569
rect 27525 29529 27537 29563
rect 27571 29560 27583 29563
rect 28074 29560 28080 29572
rect 27571 29532 28080 29560
rect 27571 29529 27583 29532
rect 27525 29523 27583 29529
rect 28074 29520 28080 29532
rect 28132 29560 28138 29572
rect 28350 29560 28356 29572
rect 28132 29532 28356 29560
rect 28132 29520 28138 29532
rect 28350 29520 28356 29532
rect 28408 29520 28414 29572
rect 28537 29563 28595 29569
rect 28537 29529 28549 29563
rect 28583 29560 28595 29563
rect 28583 29532 34100 29560
rect 28583 29529 28595 29532
rect 28537 29523 28595 29529
rect 11517 29495 11575 29501
rect 11517 29461 11529 29495
rect 11563 29492 11575 29495
rect 12434 29492 12440 29504
rect 11563 29464 12440 29492
rect 11563 29461 11575 29464
rect 11517 29455 11575 29461
rect 12434 29452 12440 29464
rect 12492 29452 12498 29504
rect 17957 29495 18015 29501
rect 17957 29461 17969 29495
rect 18003 29492 18015 29495
rect 18046 29492 18052 29504
rect 18003 29464 18052 29492
rect 18003 29461 18015 29464
rect 17957 29455 18015 29461
rect 18046 29452 18052 29464
rect 18104 29452 18110 29504
rect 21542 29452 21548 29504
rect 21600 29492 21606 29504
rect 21637 29495 21695 29501
rect 21637 29492 21649 29495
rect 21600 29464 21649 29492
rect 21600 29452 21606 29464
rect 21637 29461 21649 29464
rect 21683 29461 21695 29495
rect 21637 29455 21695 29461
rect 25317 29495 25375 29501
rect 25317 29461 25329 29495
rect 25363 29492 25375 29495
rect 25866 29492 25872 29504
rect 25363 29464 25872 29492
rect 25363 29461 25375 29464
rect 25317 29455 25375 29461
rect 25866 29452 25872 29464
rect 25924 29452 25930 29504
rect 27246 29452 27252 29504
rect 27304 29492 27310 29504
rect 29779 29495 29837 29501
rect 29779 29492 29791 29495
rect 27304 29464 29791 29492
rect 27304 29452 27310 29464
rect 29779 29461 29791 29464
rect 29825 29492 29837 29495
rect 30834 29492 30840 29504
rect 29825 29464 30840 29492
rect 29825 29461 29837 29464
rect 29779 29455 29837 29461
rect 30834 29452 30840 29464
rect 30892 29452 30898 29504
rect 30926 29452 30932 29504
rect 30984 29492 30990 29504
rect 31205 29495 31263 29501
rect 31205 29492 31217 29495
rect 30984 29464 31217 29492
rect 30984 29452 30990 29464
rect 31205 29461 31217 29464
rect 31251 29461 31263 29495
rect 31205 29455 31263 29461
rect 31478 29452 31484 29504
rect 31536 29492 31542 29504
rect 31941 29495 31999 29501
rect 31941 29492 31953 29495
rect 31536 29464 31953 29492
rect 31536 29452 31542 29464
rect 31941 29461 31953 29464
rect 31987 29461 31999 29495
rect 31941 29455 31999 29461
rect 32398 29452 32404 29504
rect 32456 29492 32462 29504
rect 33962 29492 33968 29504
rect 32456 29464 33968 29492
rect 32456 29452 32462 29464
rect 33962 29452 33968 29464
rect 34020 29452 34026 29504
rect 34072 29492 34100 29532
rect 34422 29520 34428 29572
rect 34480 29560 34486 29572
rect 35897 29563 35955 29569
rect 35897 29560 35909 29563
rect 34480 29532 35909 29560
rect 34480 29520 34486 29532
rect 35897 29529 35909 29532
rect 35943 29560 35955 29563
rect 36262 29560 36268 29572
rect 35943 29532 36268 29560
rect 35943 29529 35955 29532
rect 35897 29523 35955 29529
rect 36262 29520 36268 29532
rect 36320 29520 36326 29572
rect 36357 29495 36415 29501
rect 36357 29492 36369 29495
rect 34072 29464 36369 29492
rect 36357 29461 36369 29464
rect 36403 29461 36415 29495
rect 36357 29455 36415 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 17034 29288 17040 29300
rect 16995 29260 17040 29288
rect 17034 29248 17040 29260
rect 17092 29248 17098 29300
rect 26145 29291 26203 29297
rect 26145 29288 26157 29291
rect 24412 29260 26157 29288
rect 1762 29180 1768 29232
rect 1820 29220 1826 29232
rect 1820 29192 6914 29220
rect 1820 29180 1826 29192
rect 6886 29016 6914 29192
rect 9030 29180 9036 29232
rect 9088 29220 9094 29232
rect 9088 29192 10548 29220
rect 9088 29180 9094 29192
rect 9122 29152 9128 29164
rect 9083 29124 9128 29152
rect 9122 29112 9128 29124
rect 9180 29112 9186 29164
rect 9309 29087 9367 29093
rect 9309 29053 9321 29087
rect 9355 29084 9367 29087
rect 9766 29084 9772 29096
rect 9355 29056 9772 29084
rect 9355 29053 9367 29056
rect 9309 29047 9367 29053
rect 9766 29044 9772 29056
rect 9824 29044 9830 29096
rect 10520 29093 10548 29192
rect 12894 29180 12900 29232
rect 12952 29220 12958 29232
rect 13541 29223 13599 29229
rect 13541 29220 13553 29223
rect 12952 29192 13553 29220
rect 12952 29180 12958 29192
rect 13541 29189 13553 29192
rect 13587 29220 13599 29223
rect 14645 29223 14703 29229
rect 14645 29220 14657 29223
rect 13587 29192 14657 29220
rect 13587 29189 13599 29192
rect 13541 29183 13599 29189
rect 14645 29189 14657 29192
rect 14691 29189 14703 29223
rect 18046 29220 18052 29232
rect 14645 29183 14703 29189
rect 15580 29192 18052 29220
rect 12713 29155 12771 29161
rect 12713 29121 12725 29155
rect 12759 29152 12771 29155
rect 13446 29152 13452 29164
rect 12759 29124 13452 29152
rect 12759 29121 12771 29124
rect 12713 29115 12771 29121
rect 13446 29112 13452 29124
rect 13504 29112 13510 29164
rect 14458 29152 14464 29164
rect 14419 29124 14464 29152
rect 14458 29112 14464 29124
rect 14516 29112 14522 29164
rect 15470 29112 15476 29164
rect 15528 29152 15534 29164
rect 15580 29161 15608 29192
rect 18046 29180 18052 29192
rect 18104 29180 18110 29232
rect 19981 29223 20039 29229
rect 19981 29189 19993 29223
rect 20027 29220 20039 29223
rect 24302 29220 24308 29232
rect 20027 29192 24308 29220
rect 20027 29189 20039 29192
rect 19981 29183 20039 29189
rect 24302 29180 24308 29192
rect 24360 29180 24366 29232
rect 15565 29155 15623 29161
rect 15565 29152 15577 29155
rect 15528 29124 15577 29152
rect 15528 29112 15534 29124
rect 15565 29121 15577 29124
rect 15611 29121 15623 29155
rect 15565 29115 15623 29121
rect 15746 29112 15752 29164
rect 15804 29152 15810 29164
rect 16945 29155 17003 29161
rect 16945 29152 16957 29155
rect 15804 29124 16957 29152
rect 15804 29112 15810 29124
rect 16945 29121 16957 29124
rect 16991 29121 17003 29155
rect 16945 29115 17003 29121
rect 21266 29112 21272 29164
rect 21324 29152 21330 29164
rect 21634 29152 21640 29164
rect 21324 29124 21640 29152
rect 21324 29112 21330 29124
rect 21634 29112 21640 29124
rect 21692 29152 21698 29164
rect 21821 29155 21879 29161
rect 21821 29152 21833 29155
rect 21692 29124 21833 29152
rect 21692 29112 21698 29124
rect 21821 29121 21833 29124
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29152 22063 29155
rect 22554 29152 22560 29164
rect 22051 29124 22560 29152
rect 22051 29121 22063 29124
rect 22005 29115 22063 29121
rect 22554 29112 22560 29124
rect 22612 29112 22618 29164
rect 24412 29161 24440 29260
rect 26145 29257 26157 29260
rect 26191 29257 26203 29291
rect 26145 29251 26203 29257
rect 27157 29291 27215 29297
rect 27157 29257 27169 29291
rect 27203 29288 27215 29291
rect 27338 29288 27344 29300
rect 27203 29260 27344 29288
rect 27203 29257 27215 29260
rect 27157 29251 27215 29257
rect 27338 29248 27344 29260
rect 27396 29248 27402 29300
rect 28810 29248 28816 29300
rect 28868 29288 28874 29300
rect 30374 29288 30380 29300
rect 28868 29260 30380 29288
rect 28868 29248 28874 29260
rect 30374 29248 30380 29260
rect 30432 29248 30438 29300
rect 30650 29288 30656 29300
rect 30611 29260 30656 29288
rect 30650 29248 30656 29260
rect 30708 29248 30714 29300
rect 33962 29288 33968 29300
rect 31726 29260 33968 29288
rect 29822 29180 29828 29232
rect 29880 29220 29886 29232
rect 31726 29220 31754 29260
rect 33962 29248 33968 29260
rect 34020 29248 34026 29300
rect 34793 29223 34851 29229
rect 34793 29220 34805 29223
rect 29880 29192 30144 29220
rect 29880 29180 29886 29192
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29121 24455 29155
rect 24578 29152 24584 29164
rect 24539 29124 24584 29152
rect 24397 29115 24455 29121
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 24670 29112 24676 29164
rect 24728 29152 24734 29164
rect 24949 29155 25007 29161
rect 24949 29152 24961 29155
rect 24728 29124 24773 29152
rect 24872 29124 24961 29152
rect 24728 29112 24734 29124
rect 10505 29087 10563 29093
rect 10505 29053 10517 29087
rect 10551 29053 10563 29087
rect 14274 29084 14280 29096
rect 14235 29056 14280 29084
rect 10505 29047 10563 29053
rect 14274 29044 14280 29056
rect 14332 29044 14338 29096
rect 15194 29044 15200 29096
rect 15252 29084 15258 29096
rect 15654 29084 15660 29096
rect 15252 29056 15660 29084
rect 15252 29044 15258 29056
rect 15654 29044 15660 29056
rect 15712 29044 15718 29096
rect 15930 29084 15936 29096
rect 15891 29056 15936 29084
rect 15930 29044 15936 29056
rect 15988 29044 15994 29096
rect 18138 29084 18144 29096
rect 18099 29056 18144 29084
rect 18138 29044 18144 29056
rect 18196 29044 18202 29096
rect 18322 29084 18328 29096
rect 18283 29056 18328 29084
rect 18322 29044 18328 29056
rect 18380 29044 18386 29096
rect 24765 29087 24823 29093
rect 24765 29053 24777 29087
rect 24811 29053 24823 29087
rect 24765 29047 24823 29053
rect 24780 29016 24808 29047
rect 6886 28988 24808 29016
rect 24872 29016 24900 29124
rect 24949 29121 24961 29124
rect 24995 29121 25007 29155
rect 24949 29115 25007 29121
rect 25593 29155 25651 29161
rect 25593 29121 25605 29155
rect 25639 29121 25651 29155
rect 25866 29152 25872 29164
rect 25827 29124 25872 29152
rect 25593 29115 25651 29121
rect 25608 29084 25636 29115
rect 25866 29112 25872 29124
rect 25924 29112 25930 29164
rect 25958 29112 25964 29164
rect 26016 29152 26022 29164
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26016 29124 26985 29152
rect 26016 29112 26022 29124
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 27706 29152 27712 29164
rect 27667 29124 27712 29152
rect 26973 29115 27031 29121
rect 27706 29112 27712 29124
rect 27764 29112 27770 29164
rect 28994 29112 29000 29164
rect 29052 29152 29058 29164
rect 29730 29152 29736 29164
rect 29052 29124 29736 29152
rect 29052 29112 29058 29124
rect 29730 29112 29736 29124
rect 29788 29112 29794 29164
rect 29914 29152 29920 29164
rect 29875 29124 29920 29152
rect 29914 29112 29920 29124
rect 29972 29112 29978 29164
rect 30116 29161 30144 29192
rect 30484 29192 31754 29220
rect 32692 29192 34805 29220
rect 30101 29155 30159 29161
rect 30101 29121 30113 29155
rect 30147 29121 30159 29155
rect 30101 29115 30159 29121
rect 30193 29155 30251 29161
rect 30193 29121 30205 29155
rect 30239 29152 30251 29155
rect 30374 29152 30380 29164
rect 30239 29124 30380 29152
rect 30239 29121 30251 29124
rect 30193 29115 30251 29121
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 30484 29161 30512 29192
rect 30469 29155 30527 29161
rect 30469 29121 30481 29155
rect 30515 29121 30527 29155
rect 30469 29115 30527 29121
rect 27062 29084 27068 29096
rect 25608 29056 27068 29084
rect 27062 29044 27068 29056
rect 27120 29044 27126 29096
rect 29454 29044 29460 29096
rect 29512 29084 29518 29096
rect 30285 29087 30343 29093
rect 30285 29084 30297 29087
rect 29512 29056 30297 29084
rect 29512 29044 29518 29056
rect 30285 29053 30297 29056
rect 30331 29053 30343 29087
rect 30484 29084 30512 29115
rect 30834 29112 30840 29164
rect 30892 29112 30898 29164
rect 31018 29112 31024 29164
rect 31076 29152 31082 29164
rect 31113 29155 31171 29161
rect 31113 29152 31125 29155
rect 31076 29124 31125 29152
rect 31076 29112 31082 29124
rect 31113 29121 31125 29124
rect 31159 29121 31171 29155
rect 31386 29152 31392 29164
rect 31347 29124 31392 29152
rect 31113 29115 31171 29121
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 31570 29112 31576 29164
rect 31628 29152 31634 29164
rect 32217 29155 32275 29161
rect 32217 29152 32229 29155
rect 31628 29124 32229 29152
rect 31628 29112 31634 29124
rect 32217 29121 32229 29124
rect 32263 29121 32275 29155
rect 32582 29152 32588 29164
rect 32543 29124 32588 29152
rect 32217 29115 32275 29121
rect 32582 29112 32588 29124
rect 32640 29112 32646 29164
rect 30285 29047 30343 29053
rect 30392 29056 30512 29084
rect 30852 29084 30880 29112
rect 31297 29087 31355 29093
rect 30852 29056 31156 29084
rect 30392 29016 30420 29056
rect 24872 28988 30420 29016
rect 12618 28908 12624 28960
rect 12676 28948 12682 28960
rect 12897 28951 12955 28957
rect 12897 28948 12909 28951
rect 12676 28920 12909 28948
rect 12676 28908 12682 28920
rect 12897 28917 12909 28920
rect 12943 28917 12955 28951
rect 12897 28911 12955 28917
rect 13633 28951 13691 28957
rect 13633 28917 13645 28951
rect 13679 28948 13691 28951
rect 14642 28948 14648 28960
rect 13679 28920 14648 28948
rect 13679 28917 13691 28920
rect 13633 28911 13691 28917
rect 14642 28908 14648 28920
rect 14700 28908 14706 28960
rect 22094 28908 22100 28960
rect 22152 28948 22158 28960
rect 22189 28951 22247 28957
rect 22189 28948 22201 28951
rect 22152 28920 22201 28948
rect 22152 28908 22158 28920
rect 22189 28917 22201 28920
rect 22235 28917 22247 28951
rect 22189 28911 22247 28917
rect 24762 28908 24768 28960
rect 24820 28948 24826 28960
rect 24872 28948 24900 28988
rect 25130 28948 25136 28960
rect 24820 28920 24900 28948
rect 25091 28920 25136 28948
rect 24820 28908 24826 28920
rect 25130 28908 25136 28920
rect 25188 28908 25194 28960
rect 25682 28948 25688 28960
rect 25643 28920 25688 28948
rect 25682 28908 25688 28920
rect 25740 28908 25746 28960
rect 28902 28908 28908 28960
rect 28960 28948 28966 28960
rect 31128 28957 31156 29056
rect 31297 29053 31309 29087
rect 31343 29053 31355 29087
rect 31297 29047 31355 29053
rect 31312 29016 31340 29047
rect 32692 29016 32720 29192
rect 34793 29189 34805 29192
rect 34839 29189 34851 29223
rect 34793 29183 34851 29189
rect 33229 29155 33287 29161
rect 33229 29152 33241 29155
rect 32784 29124 33241 29152
rect 32784 29025 32812 29124
rect 33229 29121 33241 29124
rect 33275 29121 33287 29155
rect 33229 29115 33287 29121
rect 33413 29155 33471 29161
rect 33413 29121 33425 29155
rect 33459 29121 33471 29155
rect 33413 29115 33471 29121
rect 33505 29155 33563 29161
rect 33505 29121 33517 29155
rect 33551 29152 33563 29155
rect 33781 29155 33839 29161
rect 33551 29124 33732 29152
rect 33551 29121 33563 29124
rect 33505 29115 33563 29121
rect 31312 28988 32720 29016
rect 32769 29019 32827 29025
rect 32769 28985 32781 29019
rect 32815 28985 32827 29019
rect 32769 28979 32827 28985
rect 33226 28976 33232 29028
rect 33284 29016 33290 29028
rect 33428 29016 33456 29115
rect 33704 29096 33732 29124
rect 33781 29121 33793 29155
rect 33827 29152 33839 29155
rect 33870 29152 33876 29164
rect 33827 29124 33876 29152
rect 33827 29121 33839 29124
rect 33781 29115 33839 29121
rect 33870 29112 33876 29124
rect 33928 29112 33934 29164
rect 34422 29152 34428 29164
rect 34383 29124 34428 29152
rect 34422 29112 34428 29124
rect 34480 29112 34486 29164
rect 34609 29155 34667 29161
rect 34609 29121 34621 29155
rect 34655 29152 34667 29155
rect 36078 29152 36084 29164
rect 34655 29124 36084 29152
rect 34655 29121 34667 29124
rect 34609 29115 34667 29121
rect 33597 29087 33655 29093
rect 33597 29053 33609 29087
rect 33643 29053 33655 29087
rect 33597 29047 33655 29053
rect 33502 29016 33508 29028
rect 33284 28988 33508 29016
rect 33284 28976 33290 28988
rect 33502 28976 33508 28988
rect 33560 28976 33566 29028
rect 33612 28960 33640 29047
rect 33686 29044 33692 29096
rect 33744 29084 33750 29096
rect 34624 29084 34652 29115
rect 36078 29112 36084 29124
rect 36136 29112 36142 29164
rect 33744 29056 34652 29084
rect 33744 29044 33750 29056
rect 33965 29019 34023 29025
rect 33965 28985 33977 29019
rect 34011 29016 34023 29019
rect 34606 29016 34612 29028
rect 34011 28988 34612 29016
rect 34011 28985 34023 28988
rect 33965 28979 34023 28985
rect 34606 28976 34612 28988
rect 34664 28976 34670 29028
rect 28997 28951 29055 28957
rect 28997 28948 29009 28951
rect 28960 28920 29009 28948
rect 28960 28908 28966 28920
rect 28997 28917 29009 28920
rect 29043 28917 29055 28951
rect 28997 28911 29055 28917
rect 31113 28951 31171 28957
rect 31113 28917 31125 28951
rect 31159 28917 31171 28951
rect 31113 28911 31171 28917
rect 31202 28908 31208 28960
rect 31260 28948 31266 28960
rect 31570 28948 31576 28960
rect 31260 28920 31576 28948
rect 31260 28908 31266 28920
rect 31570 28908 31576 28920
rect 31628 28908 31634 28960
rect 32306 28948 32312 28960
rect 32267 28920 32312 28948
rect 32306 28908 32312 28920
rect 32364 28908 32370 28960
rect 33594 28908 33600 28960
rect 33652 28908 33658 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 9766 28744 9772 28756
rect 9727 28716 9772 28744
rect 9766 28704 9772 28716
rect 9824 28704 9830 28756
rect 13354 28704 13360 28756
rect 13412 28744 13418 28756
rect 23474 28744 23480 28756
rect 13412 28716 23480 28744
rect 13412 28704 13418 28716
rect 23474 28704 23480 28716
rect 23532 28704 23538 28756
rect 25682 28744 25688 28756
rect 24504 28716 25688 28744
rect 11238 28676 11244 28688
rect 10888 28648 11244 28676
rect 10888 28617 10916 28648
rect 11238 28636 11244 28648
rect 11296 28676 11302 28688
rect 14642 28676 14648 28688
rect 11296 28648 14648 28676
rect 11296 28636 11302 28648
rect 14642 28636 14648 28648
rect 14700 28636 14706 28688
rect 14752 28648 19334 28676
rect 10873 28611 10931 28617
rect 10873 28577 10885 28611
rect 10919 28577 10931 28611
rect 10873 28571 10931 28577
rect 11333 28611 11391 28617
rect 11333 28577 11345 28611
rect 11379 28608 11391 28611
rect 11790 28608 11796 28620
rect 11379 28580 11796 28608
rect 11379 28577 11391 28580
rect 11333 28571 11391 28577
rect 11790 28568 11796 28580
rect 11848 28568 11854 28620
rect 14550 28568 14556 28620
rect 14608 28608 14614 28620
rect 14752 28608 14780 28648
rect 14608 28580 14780 28608
rect 19306 28608 19334 28648
rect 23014 28636 23020 28688
rect 23072 28676 23078 28688
rect 24504 28676 24532 28716
rect 25682 28704 25688 28716
rect 25740 28704 25746 28756
rect 26142 28744 26148 28756
rect 26103 28716 26148 28744
rect 26142 28704 26148 28716
rect 26200 28704 26206 28756
rect 27798 28704 27804 28756
rect 27856 28744 27862 28756
rect 28445 28747 28503 28753
rect 28445 28744 28457 28747
rect 27856 28716 28457 28744
rect 27856 28704 27862 28716
rect 28445 28713 28457 28716
rect 28491 28713 28503 28747
rect 29730 28744 29736 28756
rect 29691 28716 29736 28744
rect 28445 28707 28503 28713
rect 29730 28704 29736 28716
rect 29788 28704 29794 28756
rect 29822 28704 29828 28756
rect 29880 28744 29886 28756
rect 30837 28747 30895 28753
rect 30837 28744 30849 28747
rect 29880 28716 30849 28744
rect 29880 28704 29886 28716
rect 30837 28713 30849 28716
rect 30883 28713 30895 28747
rect 30837 28707 30895 28713
rect 32582 28704 32588 28756
rect 32640 28744 32646 28756
rect 33045 28747 33103 28753
rect 33045 28744 33057 28747
rect 32640 28716 33057 28744
rect 32640 28704 32646 28716
rect 33045 28713 33057 28716
rect 33091 28713 33103 28747
rect 33045 28707 33103 28713
rect 36078 28704 36084 28756
rect 36136 28744 36142 28756
rect 36541 28747 36599 28753
rect 36541 28744 36553 28747
rect 36136 28716 36553 28744
rect 36136 28704 36142 28716
rect 36541 28713 36553 28716
rect 36587 28713 36599 28747
rect 36541 28707 36599 28713
rect 23072 28648 24532 28676
rect 25700 28676 25728 28704
rect 26510 28676 26516 28688
rect 25700 28648 26516 28676
rect 23072 28636 23078 28648
rect 26510 28636 26516 28648
rect 26568 28636 26574 28688
rect 29917 28679 29975 28685
rect 29917 28676 29929 28679
rect 27172 28648 29929 28676
rect 19306 28580 21956 28608
rect 14608 28568 14614 28580
rect 9674 28540 9680 28552
rect 9635 28512 9680 28540
rect 9674 28500 9680 28512
rect 9732 28500 9738 28552
rect 10965 28543 11023 28549
rect 10965 28509 10977 28543
rect 11011 28540 11023 28543
rect 12434 28540 12440 28552
rect 11011 28512 12440 28540
rect 11011 28509 11023 28512
rect 10965 28503 11023 28509
rect 12434 28500 12440 28512
rect 12492 28540 12498 28552
rect 13538 28540 13544 28552
rect 12492 28512 13544 28540
rect 12492 28500 12498 28512
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 15194 28540 15200 28552
rect 14691 28512 15200 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 15378 28540 15384 28552
rect 15339 28512 15384 28540
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 16114 28540 16120 28552
rect 16075 28512 16120 28540
rect 16114 28500 16120 28512
rect 16172 28500 16178 28552
rect 19334 28540 19340 28552
rect 19295 28512 19340 28540
rect 19334 28500 19340 28512
rect 19392 28500 19398 28552
rect 21082 28500 21088 28552
rect 21140 28540 21146 28552
rect 21928 28549 21956 28580
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 24673 28611 24731 28617
rect 22152 28580 23060 28608
rect 22152 28568 22158 28580
rect 23032 28549 23060 28580
rect 24673 28577 24685 28611
rect 24719 28608 24731 28611
rect 25130 28608 25136 28620
rect 24719 28580 25136 28608
rect 24719 28577 24731 28580
rect 24673 28571 24731 28577
rect 25130 28568 25136 28580
rect 25188 28568 25194 28620
rect 27062 28568 27068 28620
rect 27120 28608 27126 28620
rect 27172 28617 27200 28648
rect 29917 28645 29929 28648
rect 29963 28676 29975 28679
rect 30282 28676 30288 28688
rect 29963 28648 30288 28676
rect 29963 28645 29975 28648
rect 29917 28639 29975 28645
rect 30282 28636 30288 28648
rect 30340 28676 30346 28688
rect 31018 28676 31024 28688
rect 30340 28648 31024 28676
rect 30340 28636 30346 28648
rect 31018 28636 31024 28648
rect 31076 28636 31082 28688
rect 32306 28676 32312 28688
rect 31128 28648 32312 28676
rect 27157 28611 27215 28617
rect 27157 28608 27169 28611
rect 27120 28580 27169 28608
rect 27120 28568 27126 28580
rect 27157 28577 27169 28580
rect 27203 28577 27215 28611
rect 27157 28571 27215 28577
rect 27617 28611 27675 28617
rect 27617 28577 27629 28611
rect 27663 28577 27675 28611
rect 31128 28608 31156 28648
rect 32306 28636 32312 28648
rect 32364 28636 32370 28688
rect 27617 28571 27675 28577
rect 28000 28580 31156 28608
rect 21545 28543 21603 28549
rect 21545 28540 21557 28543
rect 21140 28512 21557 28540
rect 21140 28500 21146 28512
rect 21545 28509 21557 28512
rect 21591 28509 21603 28543
rect 21545 28503 21603 28509
rect 21913 28543 21971 28549
rect 21913 28509 21925 28543
rect 21959 28509 21971 28543
rect 21913 28503 21971 28509
rect 22741 28543 22799 28549
rect 22741 28509 22753 28543
rect 22787 28509 22799 28543
rect 22741 28503 22799 28509
rect 23017 28543 23075 28549
rect 23017 28509 23029 28543
rect 23063 28509 23075 28543
rect 24394 28540 24400 28552
rect 24355 28512 24400 28540
rect 23017 28503 23075 28509
rect 13354 28472 13360 28484
rect 13315 28444 13360 28472
rect 13354 28432 13360 28444
rect 13412 28432 13418 28484
rect 13906 28432 13912 28484
rect 13964 28472 13970 28484
rect 14093 28475 14151 28481
rect 14093 28472 14105 28475
rect 13964 28444 14105 28472
rect 13964 28432 13970 28444
rect 14093 28441 14105 28444
rect 14139 28441 14151 28475
rect 14093 28435 14151 28441
rect 14369 28475 14427 28481
rect 14369 28441 14381 28475
rect 14415 28472 14427 28475
rect 14734 28472 14740 28484
rect 14415 28444 14740 28472
rect 14415 28441 14427 28444
rect 14369 28435 14427 28441
rect 14734 28432 14740 28444
rect 14792 28472 14798 28484
rect 14792 28444 14964 28472
rect 14792 28432 14798 28444
rect 13446 28404 13452 28416
rect 13407 28376 13452 28404
rect 13446 28364 13452 28376
rect 13504 28364 13510 28416
rect 14274 28404 14280 28416
rect 14235 28376 14280 28404
rect 14274 28364 14280 28376
rect 14332 28364 14338 28416
rect 14458 28364 14464 28416
rect 14516 28404 14522 28416
rect 14936 28404 14964 28444
rect 15010 28432 15016 28484
rect 15068 28472 15074 28484
rect 15105 28475 15163 28481
rect 15105 28472 15117 28475
rect 15068 28444 15117 28472
rect 15068 28432 15074 28444
rect 15105 28441 15117 28444
rect 15151 28441 15163 28475
rect 15473 28475 15531 28481
rect 15473 28472 15485 28475
rect 15105 28435 15163 28441
rect 15212 28444 15485 28472
rect 15212 28404 15240 28444
rect 15473 28441 15485 28444
rect 15519 28441 15531 28475
rect 15473 28435 15531 28441
rect 19613 28475 19671 28481
rect 19613 28441 19625 28475
rect 19659 28441 19671 28475
rect 19613 28435 19671 28441
rect 14516 28376 14561 28404
rect 14936 28376 15240 28404
rect 14516 28364 14522 28376
rect 15286 28364 15292 28416
rect 15344 28404 15350 28416
rect 15344 28376 15389 28404
rect 15344 28364 15350 28376
rect 15562 28364 15568 28416
rect 15620 28404 15626 28416
rect 15657 28407 15715 28413
rect 15657 28404 15669 28407
rect 15620 28376 15669 28404
rect 15620 28364 15626 28376
rect 15657 28373 15669 28376
rect 15703 28373 15715 28407
rect 15657 28367 15715 28373
rect 16301 28407 16359 28413
rect 16301 28373 16313 28407
rect 16347 28404 16359 28407
rect 16666 28404 16672 28416
rect 16347 28376 16672 28404
rect 16347 28373 16359 28376
rect 16301 28367 16359 28373
rect 16666 28364 16672 28376
rect 16724 28364 16730 28416
rect 19628 28404 19656 28435
rect 20622 28432 20628 28484
rect 20680 28432 20686 28484
rect 21174 28432 21180 28484
rect 21232 28472 21238 28484
rect 21729 28475 21787 28481
rect 21729 28472 21741 28475
rect 21232 28444 21741 28472
rect 21232 28432 21238 28444
rect 21729 28441 21741 28444
rect 21775 28441 21787 28475
rect 21729 28435 21787 28441
rect 21818 28432 21824 28484
rect 21876 28472 21882 28484
rect 21876 28444 21921 28472
rect 21876 28432 21882 28444
rect 20990 28404 20996 28416
rect 19628 28376 20996 28404
rect 20990 28364 20996 28376
rect 21048 28364 21054 28416
rect 21085 28407 21143 28413
rect 21085 28373 21097 28407
rect 21131 28404 21143 28407
rect 21266 28404 21272 28416
rect 21131 28376 21272 28404
rect 21131 28373 21143 28376
rect 21085 28367 21143 28373
rect 21266 28364 21272 28376
rect 21324 28364 21330 28416
rect 22002 28364 22008 28416
rect 22060 28404 22066 28416
rect 22097 28407 22155 28413
rect 22097 28404 22109 28407
rect 22060 28376 22109 28404
rect 22060 28364 22066 28376
rect 22097 28373 22109 28376
rect 22143 28373 22155 28407
rect 22097 28367 22155 28373
rect 22278 28364 22284 28416
rect 22336 28404 22342 28416
rect 22557 28407 22615 28413
rect 22557 28404 22569 28407
rect 22336 28376 22569 28404
rect 22336 28364 22342 28376
rect 22557 28373 22569 28376
rect 22603 28373 22615 28407
rect 22756 28404 22784 28503
rect 24394 28500 24400 28512
rect 24452 28500 24458 28552
rect 27246 28540 27252 28552
rect 27207 28512 27252 28540
rect 27246 28500 27252 28512
rect 27304 28500 27310 28552
rect 22925 28475 22983 28481
rect 22925 28441 22937 28475
rect 22971 28472 22983 28475
rect 24762 28472 24768 28484
rect 22971 28444 24768 28472
rect 22971 28441 22983 28444
rect 22925 28435 22983 28441
rect 24762 28432 24768 28444
rect 24820 28432 24826 28484
rect 25958 28472 25964 28484
rect 25898 28444 25964 28472
rect 25958 28432 25964 28444
rect 26016 28432 26022 28484
rect 26234 28432 26240 28484
rect 26292 28472 26298 28484
rect 27632 28472 27660 28571
rect 26292 28444 27660 28472
rect 26292 28432 26298 28444
rect 26970 28404 26976 28416
rect 22756 28376 26976 28404
rect 22557 28367 22615 28373
rect 26970 28364 26976 28376
rect 27028 28364 27034 28416
rect 27246 28364 27252 28416
rect 27304 28404 27310 28416
rect 28000 28404 28028 28580
rect 31202 28568 31208 28620
rect 31260 28608 31266 28620
rect 33505 28611 33563 28617
rect 31260 28580 32076 28608
rect 31260 28568 31266 28580
rect 28626 28500 28632 28552
rect 28684 28540 28690 28552
rect 29549 28543 29607 28549
rect 29549 28540 29561 28543
rect 28684 28512 29561 28540
rect 28684 28500 28690 28512
rect 29549 28509 29561 28512
rect 29595 28509 29607 28543
rect 29549 28503 29607 28509
rect 29641 28543 29699 28549
rect 29641 28509 29653 28543
rect 29687 28509 29699 28543
rect 29641 28503 29699 28509
rect 30653 28543 30711 28549
rect 30653 28509 30665 28543
rect 30699 28540 30711 28543
rect 31386 28540 31392 28552
rect 30699 28512 31392 28540
rect 30699 28509 30711 28512
rect 30653 28503 30711 28509
rect 28077 28475 28135 28481
rect 28077 28441 28089 28475
rect 28123 28441 28135 28475
rect 28077 28435 28135 28441
rect 28261 28475 28319 28481
rect 28261 28441 28273 28475
rect 28307 28472 28319 28475
rect 28442 28472 28448 28484
rect 28307 28444 28448 28472
rect 28307 28441 28319 28444
rect 28261 28435 28319 28441
rect 27304 28376 28028 28404
rect 28092 28404 28120 28435
rect 28442 28432 28448 28444
rect 28500 28472 28506 28484
rect 29656 28472 29684 28503
rect 31386 28500 31392 28512
rect 31444 28500 31450 28552
rect 31754 28500 31760 28552
rect 31812 28540 31818 28552
rect 32048 28549 32076 28580
rect 33505 28577 33517 28611
rect 33551 28608 33563 28611
rect 34422 28608 34428 28620
rect 33551 28580 34428 28608
rect 33551 28577 33563 28580
rect 33505 28571 33563 28577
rect 34422 28568 34428 28580
rect 34480 28568 34486 28620
rect 34606 28568 34612 28620
rect 34664 28608 34670 28620
rect 35069 28611 35127 28617
rect 35069 28608 35081 28611
rect 34664 28580 35081 28608
rect 34664 28568 34670 28580
rect 35069 28577 35081 28580
rect 35115 28577 35127 28611
rect 35069 28571 35127 28577
rect 31849 28543 31907 28549
rect 31849 28540 31861 28543
rect 31812 28512 31861 28540
rect 31812 28500 31818 28512
rect 31849 28509 31861 28512
rect 31895 28509 31907 28543
rect 31849 28503 31907 28509
rect 32033 28543 32091 28549
rect 32033 28509 32045 28543
rect 32079 28509 32091 28543
rect 32033 28503 32091 28509
rect 33229 28543 33287 28549
rect 33229 28509 33241 28543
rect 33275 28509 33287 28543
rect 33229 28503 33287 28509
rect 28500 28444 29684 28472
rect 28500 28432 28506 28444
rect 30282 28432 30288 28484
rect 30340 28472 30346 28484
rect 30469 28475 30527 28481
rect 30469 28472 30481 28475
rect 30340 28444 30481 28472
rect 30340 28432 30346 28444
rect 30469 28441 30481 28444
rect 30515 28441 30527 28475
rect 33244 28472 33272 28503
rect 33410 28500 33416 28552
rect 33468 28540 33474 28552
rect 33468 28512 33513 28540
rect 33468 28500 33474 28512
rect 34698 28500 34704 28552
rect 34756 28540 34762 28552
rect 34793 28543 34851 28549
rect 34793 28540 34805 28543
rect 34756 28512 34805 28540
rect 34756 28500 34762 28512
rect 34793 28509 34805 28512
rect 34839 28509 34851 28543
rect 34793 28503 34851 28509
rect 46934 28500 46940 28552
rect 46992 28540 46998 28552
rect 47673 28543 47731 28549
rect 47673 28540 47685 28543
rect 46992 28512 47685 28540
rect 46992 28500 46998 28512
rect 47673 28509 47685 28512
rect 47719 28509 47731 28543
rect 47673 28503 47731 28509
rect 33686 28472 33692 28484
rect 33244 28444 33692 28472
rect 30469 28435 30527 28441
rect 33686 28432 33692 28444
rect 33744 28432 33750 28484
rect 36078 28432 36084 28484
rect 36136 28432 36142 28484
rect 29730 28404 29736 28416
rect 28092 28376 29736 28404
rect 27304 28364 27310 28376
rect 29730 28364 29736 28376
rect 29788 28364 29794 28416
rect 32217 28407 32275 28413
rect 32217 28373 32229 28407
rect 32263 28404 32275 28407
rect 32490 28404 32496 28416
rect 32263 28376 32496 28404
rect 32263 28373 32275 28376
rect 32217 28367 32275 28373
rect 32490 28364 32496 28376
rect 32548 28364 32554 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 14461 28203 14519 28209
rect 14461 28169 14473 28203
rect 14507 28169 14519 28203
rect 14461 28163 14519 28169
rect 14553 28203 14611 28209
rect 14553 28169 14565 28203
rect 14599 28200 14611 28203
rect 15562 28200 15568 28212
rect 14599 28172 15568 28200
rect 14599 28169 14611 28172
rect 14553 28163 14611 28169
rect 10962 28132 10968 28144
rect 10888 28104 10968 28132
rect 10888 28073 10916 28104
rect 10962 28092 10968 28104
rect 11020 28092 11026 28144
rect 11790 28132 11796 28144
rect 11751 28104 11796 28132
rect 11790 28092 11796 28104
rect 11848 28092 11854 28144
rect 12434 28092 12440 28144
rect 12492 28092 12498 28144
rect 13538 28132 13544 28144
rect 13499 28104 13544 28132
rect 13538 28092 13544 28104
rect 13596 28092 13602 28144
rect 14476 28132 14504 28163
rect 15562 28160 15568 28172
rect 15620 28160 15626 28212
rect 18230 28160 18236 28212
rect 18288 28200 18294 28212
rect 18417 28203 18475 28209
rect 18417 28200 18429 28203
rect 18288 28172 18429 28200
rect 18288 28160 18294 28172
rect 18417 28169 18429 28172
rect 18463 28169 18475 28203
rect 18417 28163 18475 28169
rect 20533 28203 20591 28209
rect 20533 28169 20545 28203
rect 20579 28200 20591 28203
rect 20622 28200 20628 28212
rect 20579 28172 20628 28200
rect 20579 28169 20591 28172
rect 20533 28163 20591 28169
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 21174 28200 21180 28212
rect 21135 28172 21180 28200
rect 21174 28160 21180 28172
rect 21232 28160 21238 28212
rect 21818 28160 21824 28212
rect 21876 28200 21882 28212
rect 24762 28200 24768 28212
rect 21876 28172 24768 28200
rect 21876 28160 21882 28172
rect 24762 28160 24768 28172
rect 24820 28160 24826 28212
rect 24854 28160 24860 28212
rect 24912 28200 24918 28212
rect 25685 28203 25743 28209
rect 25685 28200 25697 28203
rect 24912 28172 25697 28200
rect 24912 28160 24918 28172
rect 25685 28169 25697 28172
rect 25731 28169 25743 28203
rect 25685 28163 25743 28169
rect 26329 28203 26387 28209
rect 26329 28169 26341 28203
rect 26375 28200 26387 28203
rect 27154 28200 27160 28212
rect 26375 28172 27160 28200
rect 26375 28169 26387 28172
rect 26329 28163 26387 28169
rect 27154 28160 27160 28172
rect 27212 28160 27218 28212
rect 27430 28160 27436 28212
rect 27488 28200 27494 28212
rect 28537 28203 28595 28209
rect 28537 28200 28549 28203
rect 27488 28172 28549 28200
rect 27488 28160 27494 28172
rect 28537 28169 28549 28172
rect 28583 28200 28595 28203
rect 33873 28203 33931 28209
rect 28583 28172 33364 28200
rect 28583 28169 28595 28172
rect 28537 28163 28595 28169
rect 16945 28135 17003 28141
rect 16945 28132 16957 28135
rect 14476 28104 16957 28132
rect 16945 28101 16957 28104
rect 16991 28101 17003 28135
rect 16945 28095 17003 28101
rect 17954 28092 17960 28144
rect 18012 28092 18018 28144
rect 22094 28132 22100 28144
rect 21100 28104 22100 28132
rect 10873 28067 10931 28073
rect 10873 28033 10885 28067
rect 10919 28033 10931 28067
rect 10873 28027 10931 28033
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28064 14703 28067
rect 14734 28064 14740 28076
rect 14691 28036 14740 28064
rect 14691 28033 14703 28036
rect 14645 28027 14703 28033
rect 14734 28024 14740 28036
rect 14792 28024 14798 28076
rect 15010 28024 15016 28076
rect 15068 28064 15074 28076
rect 15289 28067 15347 28073
rect 15289 28064 15301 28067
rect 15068 28036 15301 28064
rect 15068 28024 15074 28036
rect 15289 28033 15301 28036
rect 15335 28033 15347 28067
rect 15470 28064 15476 28076
rect 15431 28036 15476 28064
rect 15289 28027 15347 28033
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11517 27999 11575 28005
rect 11517 27996 11529 27999
rect 11011 27968 11529 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11517 27965 11529 27968
rect 11563 27965 11575 27999
rect 11517 27959 11575 27965
rect 14185 27999 14243 28005
rect 14185 27965 14197 27999
rect 14231 27996 14243 27999
rect 15105 27999 15163 28005
rect 15105 27996 15117 27999
rect 14231 27968 15117 27996
rect 14231 27965 14243 27968
rect 14185 27959 14243 27965
rect 15105 27965 15117 27968
rect 15151 27965 15163 27999
rect 15304 27996 15332 28027
rect 15470 28024 15476 28036
rect 15528 28024 15534 28076
rect 15565 28067 15623 28073
rect 15565 28033 15577 28067
rect 15611 28064 15623 28067
rect 15654 28064 15660 28076
rect 15611 28036 15660 28064
rect 15611 28033 15623 28036
rect 15565 28027 15623 28033
rect 15654 28024 15660 28036
rect 15712 28024 15718 28076
rect 16666 28064 16672 28076
rect 16627 28036 16672 28064
rect 16666 28024 16672 28036
rect 16724 28024 16730 28076
rect 21100 28073 21128 28104
rect 22094 28092 22100 28104
rect 22152 28092 22158 28144
rect 24394 28092 24400 28144
rect 24452 28132 24458 28144
rect 24946 28132 24952 28144
rect 24452 28104 24952 28132
rect 24452 28092 24458 28104
rect 24946 28092 24952 28104
rect 25004 28092 25010 28144
rect 25593 28135 25651 28141
rect 25593 28101 25605 28135
rect 25639 28132 25651 28135
rect 28902 28132 28908 28144
rect 25639 28104 28908 28132
rect 25639 28101 25651 28104
rect 25593 28095 25651 28101
rect 28902 28092 28908 28104
rect 28960 28132 28966 28144
rect 30653 28135 30711 28141
rect 30653 28132 30665 28135
rect 28960 28104 30665 28132
rect 28960 28092 28966 28104
rect 30653 28101 30665 28104
rect 30699 28101 30711 28135
rect 30653 28095 30711 28101
rect 30837 28135 30895 28141
rect 30837 28101 30849 28135
rect 30883 28132 30895 28135
rect 31294 28132 31300 28144
rect 30883 28104 31300 28132
rect 30883 28101 30895 28104
rect 30837 28095 30895 28101
rect 31294 28092 31300 28104
rect 31352 28132 31358 28144
rect 31389 28135 31447 28141
rect 31389 28132 31401 28135
rect 31352 28104 31401 28132
rect 31352 28092 31358 28104
rect 31389 28101 31401 28104
rect 31435 28101 31447 28135
rect 31389 28095 31447 28101
rect 20441 28067 20499 28073
rect 20441 28033 20453 28067
rect 20487 28033 20499 28067
rect 20441 28027 20499 28033
rect 21085 28067 21143 28073
rect 21085 28033 21097 28067
rect 21131 28033 21143 28067
rect 21266 28064 21272 28076
rect 21227 28036 21272 28064
rect 21085 28027 21143 28033
rect 18138 27996 18144 28008
rect 15304 27968 18144 27996
rect 15105 27959 15163 27965
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 20456 27860 20484 28027
rect 21266 28024 21272 28036
rect 21324 28024 21330 28076
rect 22002 28064 22008 28076
rect 21963 28036 22008 28064
rect 22002 28024 22008 28036
rect 22060 28024 22066 28076
rect 22189 28067 22247 28073
rect 22189 28033 22201 28067
rect 22235 28033 22247 28067
rect 22189 28027 22247 28033
rect 20990 27956 20996 28008
rect 21048 27996 21054 28008
rect 21821 27999 21879 28005
rect 21821 27996 21833 27999
rect 21048 27968 21833 27996
rect 21048 27956 21054 27968
rect 21821 27965 21833 27968
rect 21867 27965 21879 27999
rect 22204 27996 22232 28027
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22741 28067 22799 28073
rect 22336 28036 22381 28064
rect 22336 28024 22342 28036
rect 22741 28033 22753 28067
rect 22787 28064 22799 28067
rect 23474 28064 23480 28076
rect 22787 28036 23480 28064
rect 22787 28033 22799 28036
rect 22741 28027 22799 28033
rect 23474 28024 23480 28036
rect 23532 28064 23538 28076
rect 24673 28067 24731 28073
rect 24673 28064 24685 28067
rect 23532 28036 24685 28064
rect 23532 28024 23538 28036
rect 24673 28033 24685 28036
rect 24719 28033 24731 28067
rect 26234 28064 26240 28076
rect 26195 28036 26240 28064
rect 24673 28027 24731 28033
rect 26234 28024 26240 28036
rect 26292 28024 26298 28076
rect 26421 28067 26479 28073
rect 26421 28033 26433 28067
rect 26467 28033 26479 28067
rect 27430 28064 27436 28076
rect 27391 28036 27436 28064
rect 26421 28027 26479 28033
rect 21821 27959 21879 27965
rect 21928 27968 22232 27996
rect 21266 27888 21272 27940
rect 21324 27928 21330 27940
rect 21928 27928 21956 27968
rect 21324 27900 21956 27928
rect 21324 27888 21330 27900
rect 20622 27860 20628 27872
rect 20456 27832 20628 27860
rect 20622 27820 20628 27832
rect 20680 27860 20686 27872
rect 22925 27863 22983 27869
rect 22925 27860 22937 27863
rect 20680 27832 22937 27860
rect 20680 27820 20686 27832
rect 22925 27829 22937 27832
rect 22971 27829 22983 27863
rect 22925 27823 22983 27829
rect 24857 27863 24915 27869
rect 24857 27829 24869 27863
rect 24903 27860 24915 27863
rect 25866 27860 25872 27872
rect 24903 27832 25872 27860
rect 24903 27829 24915 27832
rect 24857 27823 24915 27829
rect 25866 27820 25872 27832
rect 25924 27820 25930 27872
rect 26436 27860 26464 28027
rect 27430 28024 27436 28036
rect 27488 28024 27494 28076
rect 28350 28024 28356 28076
rect 28408 28073 28414 28076
rect 28408 28064 28417 28073
rect 29089 28067 29147 28073
rect 28408 28036 28994 28064
rect 28408 28027 28417 28036
rect 28408 28024 28414 28027
rect 27617 27999 27675 28005
rect 27617 27965 27629 27999
rect 27663 27996 27675 27999
rect 27798 27996 27804 28008
rect 27663 27968 27804 27996
rect 27663 27965 27675 27968
rect 27617 27959 27675 27965
rect 27798 27956 27804 27968
rect 27856 27956 27862 28008
rect 28966 27996 28994 28036
rect 29089 28033 29101 28067
rect 29135 28064 29147 28067
rect 29270 28064 29276 28076
rect 29135 28036 29276 28064
rect 29135 28033 29147 28036
rect 29089 28027 29147 28033
rect 29270 28024 29276 28036
rect 29328 28024 29334 28076
rect 29733 28067 29791 28073
rect 29733 28033 29745 28067
rect 29779 28064 29791 28067
rect 29914 28064 29920 28076
rect 29779 28036 29920 28064
rect 29779 28033 29791 28036
rect 29733 28027 29791 28033
rect 29914 28024 29920 28036
rect 29972 28024 29978 28076
rect 32122 28024 32128 28076
rect 32180 28064 32186 28076
rect 32309 28067 32367 28073
rect 32309 28064 32321 28067
rect 32180 28036 32321 28064
rect 32180 28024 32186 28036
rect 32309 28033 32321 28036
rect 32355 28033 32367 28067
rect 32490 28064 32496 28076
rect 32451 28036 32496 28064
rect 32309 28027 32367 28033
rect 32490 28024 32496 28036
rect 32548 28024 32554 28076
rect 33336 28064 33364 28172
rect 33873 28169 33885 28203
rect 33919 28200 33931 28203
rect 33962 28200 33968 28212
rect 33919 28172 33968 28200
rect 33919 28169 33931 28172
rect 33873 28163 33931 28169
rect 33962 28160 33968 28172
rect 34020 28160 34026 28212
rect 34609 28203 34667 28209
rect 34609 28169 34621 28203
rect 34655 28200 34667 28203
rect 34790 28200 34796 28212
rect 34655 28172 34796 28200
rect 34655 28169 34667 28172
rect 34609 28163 34667 28169
rect 34790 28160 34796 28172
rect 34848 28160 34854 28212
rect 35989 28203 36047 28209
rect 35989 28169 36001 28203
rect 36035 28200 36047 28203
rect 36078 28200 36084 28212
rect 36035 28172 36084 28200
rect 36035 28169 36047 28172
rect 35989 28163 36047 28169
rect 36078 28160 36084 28172
rect 36136 28160 36142 28212
rect 34514 28132 34520 28144
rect 33888 28104 34520 28132
rect 33781 28067 33839 28073
rect 33781 28064 33793 28067
rect 33336 28036 33793 28064
rect 33781 28033 33793 28036
rect 33827 28064 33839 28067
rect 33888 28064 33916 28104
rect 34514 28092 34520 28104
rect 34572 28092 34578 28144
rect 34422 28064 34428 28076
rect 33827 28036 33916 28064
rect 34383 28036 34428 28064
rect 33827 28033 33839 28036
rect 33781 28027 33839 28033
rect 34422 28024 34428 28036
rect 34480 28024 34486 28076
rect 34808 28064 34836 28160
rect 35253 28067 35311 28073
rect 35253 28064 35265 28067
rect 34808 28036 35265 28064
rect 35253 28033 35265 28036
rect 35299 28064 35311 28067
rect 35897 28067 35955 28073
rect 35897 28064 35909 28067
rect 35299 28036 35909 28064
rect 35299 28033 35311 28036
rect 35253 28027 35311 28033
rect 35897 28033 35909 28036
rect 35943 28033 35955 28067
rect 35897 28027 35955 28033
rect 45646 28024 45652 28076
rect 45704 28064 45710 28076
rect 45741 28067 45799 28073
rect 45741 28064 45753 28067
rect 45704 28036 45753 28064
rect 45704 28024 45710 28036
rect 45741 28033 45753 28036
rect 45787 28033 45799 28067
rect 47578 28064 47584 28076
rect 47539 28036 47584 28064
rect 45741 28027 45799 28033
rect 47578 28024 47584 28036
rect 47636 28024 47642 28076
rect 29825 27999 29883 28005
rect 29825 27996 29837 27999
rect 28966 27968 29837 27996
rect 29825 27965 29837 27968
rect 29871 27965 29883 27999
rect 29825 27959 29883 27965
rect 30558 27956 30564 28008
rect 30616 27996 30622 28008
rect 32585 27999 32643 28005
rect 32585 27996 32597 27999
rect 30616 27968 32597 27996
rect 30616 27956 30622 27968
rect 32585 27965 32597 27968
rect 32631 27965 32643 27999
rect 32585 27959 32643 27965
rect 46569 27999 46627 28005
rect 46569 27965 46581 27999
rect 46615 27996 46627 27999
rect 47394 27996 47400 28008
rect 46615 27968 47400 27996
rect 46615 27965 46627 27968
rect 46569 27959 46627 27965
rect 47394 27956 47400 27968
rect 47452 27956 47458 28008
rect 28534 27888 28540 27940
rect 28592 27928 28598 27940
rect 29181 27931 29239 27937
rect 29181 27928 29193 27931
rect 28592 27900 29193 27928
rect 28592 27888 28598 27900
rect 29181 27897 29193 27900
rect 29227 27897 29239 27931
rect 29181 27891 29239 27897
rect 31573 27931 31631 27937
rect 31573 27897 31585 27931
rect 31619 27928 31631 27931
rect 32030 27928 32036 27940
rect 31619 27900 32036 27928
rect 31619 27897 31631 27900
rect 31573 27891 31631 27897
rect 32030 27888 32036 27900
rect 32088 27888 32094 27940
rect 32398 27888 32404 27940
rect 32456 27928 32462 27940
rect 34330 27928 34336 27940
rect 32456 27900 34336 27928
rect 32456 27888 32462 27900
rect 34330 27888 34336 27900
rect 34388 27888 34394 27940
rect 35345 27931 35403 27937
rect 35345 27897 35357 27931
rect 35391 27928 35403 27931
rect 36078 27928 36084 27940
rect 35391 27900 36084 27928
rect 35391 27897 35403 27900
rect 35345 27891 35403 27897
rect 36078 27888 36084 27900
rect 36136 27888 36142 27940
rect 27614 27860 27620 27872
rect 26436 27832 27620 27860
rect 27614 27820 27620 27832
rect 27672 27820 27678 27872
rect 27982 27820 27988 27872
rect 28040 27860 28046 27872
rect 31846 27860 31852 27872
rect 28040 27832 31852 27860
rect 28040 27820 28046 27832
rect 31846 27820 31852 27832
rect 31904 27820 31910 27872
rect 31938 27820 31944 27872
rect 31996 27860 32002 27872
rect 32125 27863 32183 27869
rect 32125 27860 32137 27863
rect 31996 27832 32137 27860
rect 31996 27820 32002 27832
rect 32125 27829 32137 27832
rect 32171 27829 32183 27863
rect 32125 27823 32183 27829
rect 33318 27820 33324 27872
rect 33376 27860 33382 27872
rect 34422 27860 34428 27872
rect 33376 27832 34428 27860
rect 33376 27820 33382 27832
rect 34422 27820 34428 27832
rect 34480 27820 34486 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 3326 27616 3332 27668
rect 3384 27656 3390 27668
rect 21634 27656 21640 27668
rect 3384 27628 14596 27656
rect 21595 27628 21640 27656
rect 3384 27616 3390 27628
rect 12161 27591 12219 27597
rect 12161 27557 12173 27591
rect 12207 27588 12219 27591
rect 12434 27588 12440 27600
rect 12207 27560 12440 27588
rect 12207 27557 12219 27560
rect 12161 27551 12219 27557
rect 12434 27548 12440 27560
rect 12492 27548 12498 27600
rect 9401 27523 9459 27529
rect 9401 27489 9413 27523
rect 9447 27520 9459 27523
rect 11514 27520 11520 27532
rect 9447 27492 11520 27520
rect 9447 27489 9459 27492
rect 9401 27483 9459 27489
rect 11514 27480 11520 27492
rect 11572 27480 11578 27532
rect 14568 27529 14596 27628
rect 21634 27616 21640 27628
rect 21692 27656 21698 27668
rect 22278 27656 22284 27668
rect 21692 27628 22284 27656
rect 21692 27616 21698 27628
rect 22278 27616 22284 27628
rect 22336 27656 22342 27668
rect 22465 27659 22523 27665
rect 22465 27656 22477 27659
rect 22336 27628 22477 27656
rect 22336 27616 22342 27628
rect 22465 27625 22477 27628
rect 22511 27625 22523 27659
rect 22465 27619 22523 27625
rect 24762 27616 24768 27668
rect 24820 27656 24826 27668
rect 28074 27656 28080 27668
rect 24820 27628 28080 27656
rect 24820 27616 24826 27628
rect 28074 27616 28080 27628
rect 28132 27616 28138 27668
rect 28534 27656 28540 27668
rect 28184 27628 28540 27656
rect 18049 27591 18107 27597
rect 18049 27557 18061 27591
rect 18095 27588 18107 27591
rect 18322 27588 18328 27600
rect 18095 27560 18328 27588
rect 18095 27557 18107 27560
rect 18049 27551 18107 27557
rect 18322 27548 18328 27560
rect 18380 27548 18386 27600
rect 19242 27548 19248 27600
rect 19300 27588 19306 27600
rect 21913 27591 21971 27597
rect 21913 27588 21925 27591
rect 19300 27560 21925 27588
rect 19300 27548 19306 27560
rect 21913 27557 21925 27560
rect 21959 27588 21971 27591
rect 25774 27588 25780 27600
rect 21959 27560 25780 27588
rect 21959 27557 21971 27560
rect 21913 27551 21971 27557
rect 25774 27548 25780 27560
rect 25832 27548 25838 27600
rect 25958 27588 25964 27600
rect 25919 27560 25964 27588
rect 25958 27548 25964 27560
rect 26016 27548 26022 27600
rect 26326 27548 26332 27600
rect 26384 27588 26390 27600
rect 26970 27588 26976 27600
rect 26384 27560 26976 27588
rect 26384 27548 26390 27560
rect 26970 27548 26976 27560
rect 27028 27588 27034 27600
rect 27246 27588 27252 27600
rect 27028 27560 27252 27588
rect 27028 27548 27034 27560
rect 27246 27548 27252 27560
rect 27304 27548 27310 27600
rect 27430 27548 27436 27600
rect 27488 27588 27494 27600
rect 28184 27588 28212 27628
rect 28534 27616 28540 27628
rect 28592 27616 28598 27668
rect 30558 27616 30564 27668
rect 30616 27656 30622 27668
rect 30616 27628 31248 27656
rect 30616 27616 30622 27628
rect 27488 27560 28212 27588
rect 28353 27591 28411 27597
rect 27488 27548 27494 27560
rect 28353 27557 28365 27591
rect 28399 27588 28411 27591
rect 30282 27588 30288 27600
rect 28399 27560 30288 27588
rect 28399 27557 28411 27560
rect 28353 27551 28411 27557
rect 30282 27548 30288 27560
rect 30340 27548 30346 27600
rect 30374 27548 30380 27600
rect 30432 27588 30438 27600
rect 31220 27597 31248 27628
rect 31846 27616 31852 27668
rect 31904 27656 31910 27668
rect 33318 27656 33324 27668
rect 31904 27628 33324 27656
rect 31904 27616 31910 27628
rect 33318 27616 33324 27628
rect 33376 27616 33382 27668
rect 34958 27659 35016 27665
rect 34958 27656 34970 27659
rect 33796 27628 34970 27656
rect 30653 27591 30711 27597
rect 30653 27588 30665 27591
rect 30432 27560 30665 27588
rect 30432 27548 30438 27560
rect 30653 27557 30665 27560
rect 30699 27557 30711 27591
rect 30653 27551 30711 27557
rect 31205 27591 31263 27597
rect 31205 27557 31217 27591
rect 31251 27557 31263 27591
rect 31205 27551 31263 27557
rect 32585 27591 32643 27597
rect 32585 27557 32597 27591
rect 32631 27588 32643 27591
rect 33796 27588 33824 27628
rect 34958 27625 34970 27628
rect 35004 27625 35016 27659
rect 34958 27619 35016 27625
rect 36446 27588 36452 27600
rect 32631 27560 33824 27588
rect 36407 27560 36452 27588
rect 32631 27557 32643 27560
rect 32585 27551 32643 27557
rect 36446 27548 36452 27560
rect 36504 27548 36510 27600
rect 46934 27588 46940 27600
rect 46308 27560 46940 27588
rect 14553 27523 14611 27529
rect 14553 27489 14565 27523
rect 14599 27489 14611 27523
rect 14553 27483 14611 27489
rect 20993 27523 21051 27529
rect 20993 27489 21005 27523
rect 21039 27520 21051 27523
rect 21545 27523 21603 27529
rect 21545 27520 21557 27523
rect 21039 27492 21557 27520
rect 21039 27489 21051 27492
rect 20993 27483 21051 27489
rect 21545 27489 21557 27492
rect 21591 27520 21603 27523
rect 22554 27520 22560 27532
rect 21591 27492 22094 27520
rect 22515 27492 22560 27520
rect 21591 27489 21603 27492
rect 21545 27483 21603 27489
rect 12069 27455 12127 27461
rect 12069 27421 12081 27455
rect 12115 27452 12127 27455
rect 12526 27452 12532 27464
rect 12115 27424 12532 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 12526 27412 12532 27424
rect 12584 27412 12590 27464
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 13814 27452 13820 27464
rect 13403 27424 13820 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 14090 27452 14096 27464
rect 14051 27424 14096 27452
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 17586 27412 17592 27464
rect 17644 27452 17650 27464
rect 17957 27455 18015 27461
rect 17957 27452 17969 27455
rect 17644 27424 17969 27452
rect 17644 27412 17650 27424
rect 17957 27421 17969 27424
rect 18003 27421 18015 27455
rect 17957 27415 18015 27421
rect 20625 27455 20683 27461
rect 20625 27421 20637 27455
rect 20671 27452 20683 27455
rect 21266 27452 21272 27464
rect 20671 27424 21272 27452
rect 20671 27421 20683 27424
rect 20625 27415 20683 27421
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 21459 27455 21517 27461
rect 21459 27421 21471 27455
rect 21505 27454 21517 27455
rect 21634 27454 21640 27464
rect 21505 27426 21640 27454
rect 21505 27421 21517 27426
rect 21459 27415 21517 27421
rect 21634 27412 21640 27426
rect 21692 27412 21698 27464
rect 21729 27455 21787 27461
rect 21729 27421 21741 27455
rect 21775 27452 21787 27455
rect 21910 27452 21916 27464
rect 21775 27424 21916 27452
rect 21775 27421 21787 27424
rect 21729 27415 21787 27421
rect 21910 27412 21916 27424
rect 21968 27412 21974 27464
rect 22066 27452 22094 27492
rect 22554 27480 22560 27492
rect 22612 27480 22618 27532
rect 27338 27520 27344 27532
rect 25884 27492 27344 27520
rect 22462 27452 22468 27464
rect 22066 27424 22468 27452
rect 22462 27412 22468 27424
rect 22520 27412 22526 27464
rect 24854 27452 24860 27464
rect 24815 27424 24860 27452
rect 24854 27412 24860 27424
rect 24912 27412 24918 27464
rect 25884 27461 25912 27492
rect 27338 27480 27344 27492
rect 27396 27480 27402 27532
rect 29822 27520 29828 27532
rect 28552 27492 29828 27520
rect 25869 27455 25927 27461
rect 25869 27421 25881 27455
rect 25915 27421 25927 27455
rect 27062 27452 27068 27464
rect 27023 27424 27068 27452
rect 25869 27415 25927 27421
rect 27062 27412 27068 27424
rect 27120 27412 27126 27464
rect 28552 27461 28580 27492
rect 29822 27480 29828 27492
rect 29880 27480 29886 27532
rect 33410 27520 33416 27532
rect 30944 27492 33416 27520
rect 30944 27464 30972 27492
rect 33410 27480 33416 27492
rect 33468 27480 33474 27532
rect 34698 27520 34704 27532
rect 34659 27492 34704 27520
rect 34698 27480 34704 27492
rect 34756 27480 34762 27532
rect 46308 27529 46336 27560
rect 46934 27548 46940 27560
rect 46992 27548 46998 27600
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46293 27483 46351 27489
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 47670 27520 47676 27532
rect 46523 27492 47676 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 47670 27480 47676 27492
rect 47728 27480 47734 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27421 28595 27455
rect 28537 27415 28595 27421
rect 28721 27455 28779 27461
rect 28721 27421 28733 27455
rect 28767 27452 28779 27455
rect 29362 27452 29368 27464
rect 28767 27424 29368 27452
rect 28767 27421 28779 27424
rect 28721 27415 28779 27421
rect 29362 27412 29368 27424
rect 29420 27412 29426 27464
rect 29546 27412 29552 27464
rect 29604 27452 29610 27464
rect 29641 27455 29699 27461
rect 29641 27452 29653 27455
rect 29604 27424 29653 27452
rect 29604 27412 29610 27424
rect 29641 27421 29653 27424
rect 29687 27421 29699 27455
rect 29641 27415 29699 27421
rect 30561 27455 30619 27461
rect 30561 27421 30573 27455
rect 30607 27421 30619 27455
rect 30561 27415 30619 27421
rect 30745 27455 30803 27461
rect 30745 27421 30757 27455
rect 30791 27452 30803 27455
rect 30926 27452 30932 27464
rect 30791 27424 30932 27452
rect 30791 27421 30803 27424
rect 30745 27415 30803 27421
rect 9585 27387 9643 27393
rect 9585 27353 9597 27387
rect 9631 27384 9643 27387
rect 9766 27384 9772 27396
rect 9631 27356 9772 27384
rect 9631 27353 9643 27356
rect 9585 27347 9643 27353
rect 9766 27344 9772 27356
rect 9824 27344 9830 27396
rect 11241 27387 11299 27393
rect 11241 27384 11253 27387
rect 10980 27356 11253 27384
rect 7558 27276 7564 27328
rect 7616 27316 7622 27328
rect 10980 27316 11008 27356
rect 11241 27353 11253 27356
rect 11287 27353 11299 27387
rect 11241 27347 11299 27353
rect 13449 27387 13507 27393
rect 13449 27353 13461 27387
rect 13495 27384 13507 27387
rect 14277 27387 14335 27393
rect 14277 27384 14289 27387
rect 13495 27356 14289 27384
rect 13495 27353 13507 27356
rect 13449 27347 13507 27353
rect 14277 27353 14289 27356
rect 14323 27353 14335 27387
rect 20806 27384 20812 27396
rect 20767 27356 20812 27384
rect 14277 27347 14335 27353
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 28813 27387 28871 27393
rect 28813 27384 28825 27387
rect 20916 27356 28825 27384
rect 7616 27288 11008 27316
rect 7616 27276 7622 27288
rect 14366 27276 14372 27328
rect 14424 27316 14430 27328
rect 15470 27316 15476 27328
rect 14424 27288 15476 27316
rect 14424 27276 14430 27288
rect 15470 27276 15476 27288
rect 15528 27316 15534 27328
rect 20916 27316 20944 27356
rect 28813 27353 28825 27356
rect 28859 27353 28871 27387
rect 30576 27384 30604 27415
rect 30926 27412 30932 27424
rect 30984 27412 30990 27464
rect 31202 27452 31208 27464
rect 31163 27424 31208 27452
rect 31202 27412 31208 27424
rect 31260 27412 31266 27464
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27452 31447 27455
rect 31938 27452 31944 27464
rect 31435 27424 31754 27452
rect 31899 27424 31944 27452
rect 31435 27421 31447 27424
rect 31389 27415 31447 27421
rect 31726 27396 31754 27424
rect 31938 27412 31944 27424
rect 31996 27412 32002 27464
rect 32034 27455 32092 27461
rect 32034 27421 32046 27455
rect 32080 27421 32092 27455
rect 32034 27415 32092 27421
rect 31478 27384 31484 27396
rect 30576 27356 31484 27384
rect 28813 27347 28871 27353
rect 31478 27344 31484 27356
rect 31536 27344 31542 27396
rect 31726 27356 31760 27396
rect 31754 27344 31760 27356
rect 31812 27384 31818 27396
rect 32048 27384 32076 27415
rect 32214 27412 32220 27464
rect 32272 27452 32278 27464
rect 32490 27461 32496 27464
rect 32447 27455 32496 27461
rect 32272 27424 32317 27452
rect 32272 27412 32278 27424
rect 32447 27421 32459 27455
rect 32493 27421 32496 27455
rect 32447 27415 32496 27421
rect 32490 27412 32496 27415
rect 32548 27412 32554 27464
rect 36078 27412 36084 27464
rect 36136 27412 36142 27464
rect 45646 27452 45652 27464
rect 45607 27424 45652 27452
rect 45646 27412 45652 27424
rect 45704 27412 45710 27464
rect 31812 27356 32076 27384
rect 31812 27344 31818 27356
rect 22830 27316 22836 27328
rect 15528 27288 20944 27316
rect 22791 27288 22836 27316
rect 15528 27276 15534 27288
rect 22830 27276 22836 27288
rect 22888 27276 22894 27328
rect 24946 27316 24952 27328
rect 24907 27288 24952 27316
rect 24946 27276 24952 27288
rect 25004 27276 25010 27328
rect 27154 27276 27160 27328
rect 27212 27316 27218 27328
rect 29825 27319 29883 27325
rect 29825 27316 29837 27319
rect 27212 27288 29837 27316
rect 27212 27276 27218 27288
rect 29825 27285 29837 27288
rect 29871 27316 29883 27319
rect 32232 27316 32260 27412
rect 32306 27344 32312 27396
rect 32364 27384 32370 27396
rect 32766 27384 32772 27396
rect 32364 27356 32772 27384
rect 32364 27344 32370 27356
rect 32766 27344 32772 27356
rect 32824 27344 32830 27396
rect 45738 27316 45744 27328
rect 29871 27288 32260 27316
rect 45699 27288 45744 27316
rect 29871 27285 29883 27288
rect 29825 27279 29883 27285
rect 45738 27276 45744 27288
rect 45796 27276 45802 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 9766 27112 9772 27124
rect 9727 27084 9772 27112
rect 9766 27072 9772 27084
rect 9824 27072 9830 27124
rect 14458 27072 14464 27124
rect 14516 27112 14522 27124
rect 14645 27115 14703 27121
rect 14645 27112 14657 27115
rect 14516 27084 14657 27112
rect 14516 27072 14522 27084
rect 14645 27081 14657 27084
rect 14691 27081 14703 27115
rect 14645 27075 14703 27081
rect 14734 27072 14740 27124
rect 14792 27112 14798 27124
rect 15473 27115 15531 27121
rect 14792 27084 15424 27112
rect 14792 27072 14798 27084
rect 11882 27004 11888 27056
rect 11940 27044 11946 27056
rect 11940 27016 12282 27044
rect 11940 27004 11946 27016
rect 14090 27004 14096 27056
rect 14148 27044 14154 27056
rect 15396 27044 15424 27084
rect 15473 27081 15485 27115
rect 15519 27112 15531 27115
rect 15562 27112 15568 27124
rect 15519 27084 15568 27112
rect 15519 27081 15531 27084
rect 15473 27075 15531 27081
rect 15562 27072 15568 27084
rect 15620 27072 15626 27124
rect 17405 27115 17463 27121
rect 17405 27081 17417 27115
rect 17451 27112 17463 27115
rect 17954 27112 17960 27124
rect 17451 27084 17960 27112
rect 17451 27081 17463 27084
rect 17405 27075 17463 27081
rect 17954 27072 17960 27084
rect 18012 27072 18018 27124
rect 23109 27115 23167 27121
rect 23109 27112 23121 27115
rect 20824 27084 23121 27112
rect 14148 27016 15332 27044
rect 15396 27016 15608 27044
rect 14148 27004 14154 27016
rect 9674 26976 9680 26988
rect 9635 26948 9680 26976
rect 9674 26936 9680 26948
rect 9732 26936 9738 26988
rect 10778 26976 10784 26988
rect 10691 26948 10784 26976
rect 10778 26936 10784 26948
rect 10836 26976 10842 26988
rect 10962 26976 10968 26988
rect 10836 26948 10968 26976
rect 10836 26936 10842 26948
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 14461 26979 14519 26985
rect 14461 26945 14473 26979
rect 14507 26976 14519 26979
rect 14550 26976 14556 26988
rect 14507 26948 14556 26976
rect 14507 26945 14519 26948
rect 14461 26939 14519 26945
rect 14550 26936 14556 26948
rect 14608 26936 14614 26988
rect 15304 26985 15332 27016
rect 15289 26979 15347 26985
rect 15289 26945 15301 26979
rect 15335 26976 15347 26979
rect 15378 26976 15384 26988
rect 15335 26948 15384 26976
rect 15335 26945 15347 26948
rect 15289 26939 15347 26945
rect 15378 26936 15384 26948
rect 15436 26936 15442 26988
rect 15580 26985 15608 27016
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26945 15623 26979
rect 15565 26939 15623 26945
rect 17313 26979 17371 26985
rect 17313 26945 17325 26979
rect 17359 26976 17371 26979
rect 17402 26976 17408 26988
rect 17359 26948 17408 26976
rect 17359 26945 17371 26948
rect 17313 26939 17371 26945
rect 17402 26936 17408 26948
rect 17460 26936 17466 26988
rect 17954 26976 17960 26988
rect 17915 26948 17960 26976
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 20824 26985 20852 27084
rect 23109 27081 23121 27084
rect 23155 27081 23167 27115
rect 26329 27115 26387 27121
rect 26329 27112 26341 27115
rect 23109 27075 23167 27081
rect 24136 27084 26341 27112
rect 21174 27044 21180 27056
rect 20916 27016 21180 27044
rect 20916 26985 20944 27016
rect 21174 27004 21180 27016
rect 21232 27004 21238 27056
rect 21269 27047 21327 27053
rect 21269 27013 21281 27047
rect 21315 27044 21327 27047
rect 21315 27016 21864 27044
rect 21315 27013 21327 27016
rect 21269 27007 21327 27013
rect 20809 26979 20867 26985
rect 20809 26945 20821 26979
rect 20855 26945 20867 26979
rect 20809 26939 20867 26945
rect 20901 26979 20959 26985
rect 20901 26945 20913 26979
rect 20947 26945 20959 26979
rect 21082 26976 21088 26988
rect 21043 26948 21088 26976
rect 20901 26939 20959 26945
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 21836 26985 21864 27016
rect 22296 27016 23060 27044
rect 21821 26979 21879 26985
rect 21821 26945 21833 26979
rect 21867 26945 21879 26979
rect 22002 26976 22008 26988
rect 21963 26948 22008 26976
rect 21821 26939 21879 26945
rect 22002 26936 22008 26948
rect 22060 26936 22066 26988
rect 22186 26976 22192 26988
rect 22147 26948 22192 26976
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 10873 26911 10931 26917
rect 10873 26877 10885 26911
rect 10919 26908 10931 26911
rect 11517 26911 11575 26917
rect 11517 26908 11529 26911
rect 10919 26880 11529 26908
rect 10919 26877 10931 26880
rect 10873 26871 10931 26877
rect 11517 26877 11529 26880
rect 11563 26877 11575 26911
rect 11793 26911 11851 26917
rect 11793 26908 11805 26911
rect 11517 26871 11575 26877
rect 11624 26880 11805 26908
rect 11054 26800 11060 26852
rect 11112 26840 11118 26852
rect 11624 26840 11652 26880
rect 11793 26877 11805 26880
rect 11839 26877 11851 26911
rect 11793 26871 11851 26877
rect 14277 26911 14335 26917
rect 14277 26877 14289 26911
rect 14323 26908 14335 26911
rect 14826 26908 14832 26920
rect 14323 26880 14832 26908
rect 14323 26877 14335 26880
rect 14277 26871 14335 26877
rect 14826 26868 14832 26880
rect 14884 26868 14890 26920
rect 18138 26908 18144 26920
rect 18099 26880 18144 26908
rect 18138 26868 18144 26880
rect 18196 26868 18202 26920
rect 19797 26911 19855 26917
rect 19797 26877 19809 26911
rect 19843 26908 19855 26911
rect 20254 26908 20260 26920
rect 19843 26880 20260 26908
rect 19843 26877 19855 26880
rect 19797 26871 19855 26877
rect 20254 26868 20260 26880
rect 20312 26868 20318 26920
rect 21177 26911 21235 26917
rect 21177 26877 21189 26911
rect 21223 26908 21235 26911
rect 21450 26908 21456 26920
rect 21223 26880 21456 26908
rect 21223 26877 21235 26880
rect 21177 26871 21235 26877
rect 21450 26868 21456 26880
rect 21508 26868 21514 26920
rect 22097 26911 22155 26917
rect 22097 26877 22109 26911
rect 22143 26877 22155 26911
rect 22097 26871 22155 26877
rect 11112 26812 11652 26840
rect 11112 26800 11118 26812
rect 13814 26800 13820 26852
rect 13872 26840 13878 26852
rect 17586 26840 17592 26852
rect 13872 26812 17592 26840
rect 13872 26800 13878 26812
rect 17586 26800 17592 26812
rect 17644 26800 17650 26852
rect 21082 26800 21088 26852
rect 21140 26840 21146 26852
rect 22112 26840 22140 26871
rect 22296 26840 22324 27016
rect 23032 26985 23060 27016
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26974 22431 26979
rect 23017 26979 23075 26985
rect 22419 26946 22508 26974
rect 22419 26945 22431 26946
rect 22373 26939 22431 26945
rect 22480 26908 22508 26946
rect 23017 26945 23029 26979
rect 23063 26945 23075 26979
rect 23017 26939 23075 26945
rect 22738 26908 22744 26920
rect 22480 26880 22744 26908
rect 22738 26868 22744 26880
rect 22796 26908 22802 26920
rect 24136 26908 24164 27084
rect 26329 27081 26341 27084
rect 26375 27112 26387 27115
rect 26375 27084 27568 27112
rect 26375 27081 26387 27084
rect 26329 27075 26387 27081
rect 25774 27004 25780 27056
rect 25832 27044 25838 27056
rect 27154 27044 27160 27056
rect 25832 27016 27160 27044
rect 25832 27004 25838 27016
rect 27154 27004 27160 27016
rect 27212 27044 27218 27056
rect 27433 27047 27491 27053
rect 27433 27044 27445 27047
rect 27212 27016 27445 27044
rect 27212 27004 27218 27016
rect 27433 27013 27445 27016
rect 27479 27013 27491 27047
rect 27433 27007 27491 27013
rect 24210 26936 24216 26988
rect 24268 26976 24274 26988
rect 24268 26948 24313 26976
rect 24268 26936 24274 26948
rect 26050 26936 26056 26988
rect 26108 26976 26114 26988
rect 26145 26979 26203 26985
rect 26145 26976 26157 26979
rect 26108 26948 26157 26976
rect 26108 26936 26114 26948
rect 26145 26945 26157 26948
rect 26191 26945 26203 26979
rect 26145 26939 26203 26945
rect 22796 26880 24164 26908
rect 24489 26911 24547 26917
rect 22796 26868 22802 26880
rect 24489 26877 24501 26911
rect 24535 26908 24547 26911
rect 24854 26908 24860 26920
rect 24535 26880 24860 26908
rect 24535 26877 24547 26880
rect 24489 26871 24547 26877
rect 24854 26868 24860 26880
rect 24912 26868 24918 26920
rect 27540 26908 27568 27084
rect 27632 27084 28396 27112
rect 27632 27053 27660 27084
rect 28368 27053 28396 27084
rect 31754 27072 31760 27124
rect 31812 27112 31818 27124
rect 36446 27112 36452 27124
rect 31812 27084 36452 27112
rect 31812 27072 31818 27084
rect 36446 27072 36452 27084
rect 36504 27072 36510 27124
rect 46566 27112 46572 27124
rect 46527 27084 46572 27112
rect 46566 27072 46572 27084
rect 46624 27072 46630 27124
rect 27617 27047 27675 27053
rect 27617 27013 27629 27047
rect 27663 27013 27675 27047
rect 27617 27007 27675 27013
rect 28169 27047 28227 27053
rect 28169 27013 28181 27047
rect 28215 27013 28227 27047
rect 28368 27047 28443 27053
rect 28368 27016 28397 27047
rect 28169 27007 28227 27013
rect 28385 27013 28397 27016
rect 28431 27044 28443 27047
rect 29178 27044 29184 27056
rect 28431 27016 29184 27044
rect 28431 27013 28443 27016
rect 28385 27007 28443 27013
rect 28184 26976 28212 27007
rect 29178 27004 29184 27016
rect 29236 27004 29242 27056
rect 30377 27047 30435 27053
rect 30377 27013 30389 27047
rect 30423 27044 30435 27047
rect 32858 27044 32864 27056
rect 30423 27016 32864 27044
rect 30423 27013 30435 27016
rect 30377 27007 30435 27013
rect 32858 27004 32864 27016
rect 32916 27004 32922 27056
rect 29362 26976 29368 26988
rect 28184 26948 29368 26976
rect 29362 26936 29368 26948
rect 29420 26936 29426 26988
rect 30285 26979 30343 26985
rect 30285 26976 30297 26979
rect 29472 26948 30297 26976
rect 28994 26908 29000 26920
rect 27540 26880 29000 26908
rect 28994 26868 29000 26880
rect 29052 26868 29058 26920
rect 29178 26908 29184 26920
rect 29139 26880 29184 26908
rect 29178 26868 29184 26880
rect 29236 26868 29242 26920
rect 21140 26812 22324 26840
rect 21140 26800 21146 26812
rect 22830 26800 22836 26852
rect 22888 26840 22894 26852
rect 24305 26843 24363 26849
rect 24305 26840 24317 26843
rect 22888 26812 24317 26840
rect 22888 26800 22894 26812
rect 24305 26809 24317 26812
rect 24351 26840 24363 26843
rect 24670 26840 24676 26852
rect 24351 26812 24676 26840
rect 24351 26809 24363 26812
rect 24305 26803 24363 26809
rect 24670 26800 24676 26812
rect 24728 26800 24734 26852
rect 26142 26800 26148 26852
rect 26200 26840 26206 26852
rect 29472 26840 29500 26948
rect 30285 26945 30297 26948
rect 30331 26945 30343 26979
rect 30285 26939 30343 26945
rect 31018 26936 31024 26988
rect 31076 26976 31082 26988
rect 31113 26979 31171 26985
rect 31113 26976 31125 26979
rect 31076 26948 31125 26976
rect 31076 26936 31082 26948
rect 31113 26945 31125 26948
rect 31159 26945 31171 26979
rect 31113 26939 31171 26945
rect 45281 26979 45339 26985
rect 45281 26945 45293 26979
rect 45327 26976 45339 26979
rect 45646 26976 45652 26988
rect 45327 26948 45652 26976
rect 45327 26945 45339 26948
rect 45281 26939 45339 26945
rect 45646 26936 45652 26948
rect 45704 26936 45710 26988
rect 29733 26911 29791 26917
rect 29733 26877 29745 26911
rect 29779 26908 29791 26911
rect 29822 26908 29828 26920
rect 29779 26880 29828 26908
rect 29779 26877 29791 26880
rect 29733 26871 29791 26877
rect 29822 26868 29828 26880
rect 29880 26868 29886 26920
rect 30929 26911 30987 26917
rect 30929 26877 30941 26911
rect 30975 26908 30987 26911
rect 31846 26908 31852 26920
rect 30975 26880 31852 26908
rect 30975 26877 30987 26880
rect 30929 26871 30987 26877
rect 31846 26868 31852 26880
rect 31904 26868 31910 26920
rect 33042 26868 33048 26920
rect 33100 26908 33106 26920
rect 46382 26908 46388 26920
rect 33100 26880 46388 26908
rect 33100 26868 33106 26880
rect 46382 26868 46388 26880
rect 46440 26868 46446 26920
rect 26200 26812 29500 26840
rect 26200 26800 26206 26812
rect 29546 26800 29552 26852
rect 29604 26840 29610 26852
rect 29641 26843 29699 26849
rect 29641 26840 29653 26843
rect 29604 26812 29653 26840
rect 29604 26800 29610 26812
rect 29641 26809 29653 26812
rect 29687 26809 29699 26843
rect 29641 26803 29699 26809
rect 30466 26800 30472 26852
rect 30524 26840 30530 26852
rect 32766 26840 32772 26852
rect 30524 26812 32772 26840
rect 30524 26800 30530 26812
rect 32766 26800 32772 26812
rect 32824 26800 32830 26852
rect 13078 26732 13084 26784
rect 13136 26772 13142 26784
rect 13265 26775 13323 26781
rect 13265 26772 13277 26775
rect 13136 26744 13277 26772
rect 13136 26732 13142 26744
rect 13265 26741 13277 26744
rect 13311 26741 13323 26775
rect 15286 26772 15292 26784
rect 15247 26744 15292 26772
rect 13265 26735 13323 26741
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 20714 26772 20720 26784
rect 19484 26744 20720 26772
rect 19484 26732 19490 26744
rect 20714 26732 20720 26744
rect 20772 26732 20778 26784
rect 20990 26732 20996 26784
rect 21048 26772 21054 26784
rect 22557 26775 22615 26781
rect 22557 26772 22569 26775
rect 21048 26744 22569 26772
rect 21048 26732 21054 26744
rect 22557 26741 22569 26744
rect 22603 26741 22615 26775
rect 22557 26735 22615 26741
rect 24397 26775 24455 26781
rect 24397 26741 24409 26775
rect 24443 26772 24455 26775
rect 25130 26772 25136 26784
rect 24443 26744 25136 26772
rect 24443 26741 24455 26744
rect 24397 26735 24455 26741
rect 25130 26732 25136 26744
rect 25188 26732 25194 26784
rect 26050 26732 26056 26784
rect 26108 26772 26114 26784
rect 27890 26772 27896 26784
rect 26108 26744 27896 26772
rect 26108 26732 26114 26744
rect 27890 26732 27896 26744
rect 27948 26732 27954 26784
rect 28350 26772 28356 26784
rect 28311 26744 28356 26772
rect 28350 26732 28356 26744
rect 28408 26732 28414 26784
rect 28534 26772 28540 26784
rect 28495 26744 28540 26772
rect 28534 26732 28540 26744
rect 28592 26732 28598 26784
rect 30834 26732 30840 26784
rect 30892 26772 30898 26784
rect 31297 26775 31355 26781
rect 31297 26772 31309 26775
rect 30892 26744 31309 26772
rect 30892 26732 30898 26744
rect 31297 26741 31309 26744
rect 31343 26741 31355 26775
rect 31297 26735 31355 26741
rect 46658 26732 46664 26784
rect 46716 26772 46722 26784
rect 47765 26775 47823 26781
rect 47765 26772 47777 26775
rect 46716 26744 47777 26772
rect 46716 26732 46722 26744
rect 47765 26741 47777 26744
rect 47811 26741 47823 26775
rect 47765 26735 47823 26741
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 11054 26568 11060 26580
rect 11015 26540 11060 26568
rect 11054 26528 11060 26540
rect 11112 26528 11118 26580
rect 11882 26568 11888 26580
rect 11843 26540 11888 26568
rect 11882 26528 11888 26540
rect 11940 26528 11946 26580
rect 15378 26568 15384 26580
rect 14660 26540 15384 26568
rect 14660 26509 14688 26540
rect 15378 26528 15384 26540
rect 15436 26568 15442 26580
rect 17405 26571 17463 26577
rect 17405 26568 17417 26571
rect 15436 26540 17417 26568
rect 15436 26528 15442 26540
rect 17405 26537 17417 26540
rect 17451 26537 17463 26571
rect 17405 26531 17463 26537
rect 17957 26571 18015 26577
rect 17957 26537 17969 26571
rect 18003 26568 18015 26571
rect 18138 26568 18144 26580
rect 18003 26540 18144 26568
rect 18003 26537 18015 26540
rect 17957 26531 18015 26537
rect 18138 26528 18144 26540
rect 18196 26528 18202 26580
rect 19692 26571 19750 26577
rect 19692 26537 19704 26571
rect 19738 26568 19750 26571
rect 20990 26568 20996 26580
rect 19738 26540 20996 26568
rect 19738 26537 19750 26540
rect 19692 26531 19750 26537
rect 20990 26528 20996 26540
rect 21048 26528 21054 26580
rect 21082 26528 21088 26580
rect 21140 26568 21146 26580
rect 21177 26571 21235 26577
rect 21177 26568 21189 26571
rect 21140 26540 21189 26568
rect 21140 26528 21146 26540
rect 21177 26537 21189 26540
rect 21223 26537 21235 26571
rect 21177 26531 21235 26537
rect 21450 26528 21456 26580
rect 21508 26568 21514 26580
rect 22189 26571 22247 26577
rect 21508 26540 21864 26568
rect 21508 26528 21514 26540
rect 13081 26503 13139 26509
rect 13081 26500 13093 26503
rect 12544 26472 13093 26500
rect 12544 26376 12572 26472
rect 13081 26469 13093 26472
rect 13127 26469 13139 26503
rect 13081 26463 13139 26469
rect 14645 26503 14703 26509
rect 14645 26469 14657 26503
rect 14691 26469 14703 26503
rect 14645 26463 14703 26469
rect 20714 26460 20720 26512
rect 20772 26500 20778 26512
rect 21729 26503 21787 26509
rect 21729 26500 21741 26503
rect 20772 26472 21741 26500
rect 20772 26460 20778 26472
rect 21729 26469 21741 26472
rect 21775 26469 21787 26503
rect 21729 26463 21787 26469
rect 15197 26435 15255 26441
rect 15197 26401 15209 26435
rect 15243 26432 15255 26435
rect 15243 26404 18828 26432
rect 15243 26401 15255 26404
rect 15197 26395 15255 26401
rect 11054 26364 11060 26376
rect 11015 26336 11060 26364
rect 11054 26324 11060 26336
rect 11112 26324 11118 26376
rect 11238 26364 11244 26376
rect 11199 26336 11244 26364
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 11793 26367 11851 26373
rect 11793 26333 11805 26367
rect 11839 26364 11851 26367
rect 12526 26364 12532 26376
rect 11839 26336 12532 26364
rect 11839 26333 11851 26336
rect 11793 26327 11851 26333
rect 12526 26324 12532 26336
rect 12584 26324 12590 26376
rect 12897 26367 12955 26373
rect 12897 26333 12909 26367
rect 12943 26364 12955 26367
rect 13446 26364 13452 26376
rect 12943 26336 13452 26364
rect 12943 26333 12955 26336
rect 12897 26327 12955 26333
rect 13446 26324 13452 26336
rect 13504 26364 13510 26376
rect 14918 26364 14924 26376
rect 13504 26336 14924 26364
rect 13504 26324 13510 26336
rect 14918 26324 14924 26336
rect 14976 26324 14982 26376
rect 15654 26364 15660 26376
rect 15615 26336 15660 26364
rect 15654 26324 15660 26336
rect 15712 26324 15718 26376
rect 17586 26324 17592 26376
rect 17644 26364 17650 26376
rect 17865 26367 17923 26373
rect 17865 26364 17877 26367
rect 17644 26336 17877 26364
rect 17644 26324 17650 26336
rect 17865 26333 17877 26336
rect 17911 26333 17923 26367
rect 18800 26364 18828 26404
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19429 26435 19487 26441
rect 19429 26432 19441 26435
rect 19392 26404 19441 26432
rect 19392 26392 19398 26404
rect 19429 26401 19441 26404
rect 19475 26432 19487 26435
rect 20070 26432 20076 26444
rect 19475 26404 20076 26432
rect 19475 26401 19487 26404
rect 19429 26395 19487 26401
rect 20070 26392 20076 26404
rect 20128 26392 20134 26444
rect 21836 26364 21864 26540
rect 22189 26537 22201 26571
rect 22235 26568 22247 26571
rect 22462 26568 22468 26580
rect 22235 26540 22468 26568
rect 22235 26537 22247 26540
rect 22189 26531 22247 26537
rect 22462 26528 22468 26540
rect 22520 26528 22526 26580
rect 24210 26528 24216 26580
rect 24268 26568 24274 26580
rect 24765 26571 24823 26577
rect 24765 26568 24777 26571
rect 24268 26540 24777 26568
rect 24268 26528 24274 26540
rect 24765 26537 24777 26540
rect 24811 26568 24823 26571
rect 26510 26568 26516 26580
rect 24811 26540 26096 26568
rect 26471 26540 26516 26568
rect 24811 26537 24823 26540
rect 24765 26531 24823 26537
rect 25332 26512 25360 26540
rect 22094 26460 22100 26512
rect 22152 26500 22158 26512
rect 23845 26503 23903 26509
rect 23845 26500 23857 26503
rect 22152 26472 22416 26500
rect 22152 26460 22158 26472
rect 22278 26432 22284 26444
rect 22239 26404 22284 26432
rect 22278 26392 22284 26404
rect 22336 26392 22342 26444
rect 22388 26373 22416 26472
rect 22664 26472 23857 26500
rect 22005 26367 22063 26373
rect 22005 26364 22017 26367
rect 18800 26336 19334 26364
rect 21836 26336 22017 26364
rect 17865 26327 17923 26333
rect 14826 26296 14832 26308
rect 14787 26268 14832 26296
rect 14826 26256 14832 26268
rect 14884 26256 14890 26308
rect 15013 26299 15071 26305
rect 15013 26265 15025 26299
rect 15059 26296 15071 26299
rect 15562 26296 15568 26308
rect 15059 26268 15568 26296
rect 15059 26265 15071 26268
rect 15013 26259 15071 26265
rect 15562 26256 15568 26268
rect 15620 26256 15626 26308
rect 15930 26296 15936 26308
rect 15891 26268 15936 26296
rect 15930 26256 15936 26268
rect 15988 26256 15994 26308
rect 18782 26296 18788 26308
rect 17158 26268 18788 26296
rect 18782 26256 18788 26268
rect 18840 26256 18846 26308
rect 14550 26188 14556 26240
rect 14608 26228 14614 26240
rect 14921 26231 14979 26237
rect 14921 26228 14933 26231
rect 14608 26200 14933 26228
rect 14608 26188 14614 26200
rect 14921 26197 14933 26200
rect 14967 26197 14979 26231
rect 19306 26228 19334 26336
rect 22005 26333 22017 26336
rect 22051 26333 22063 26367
rect 22005 26327 22063 26333
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26364 22155 26367
rect 22373 26367 22431 26373
rect 22143 26336 22177 26364
rect 22143 26333 22155 26336
rect 22097 26327 22155 26333
rect 22373 26333 22385 26367
rect 22419 26333 22431 26367
rect 22373 26327 22431 26333
rect 20714 26256 20720 26308
rect 20772 26256 20778 26308
rect 21634 26256 21640 26308
rect 21692 26296 21698 26308
rect 22112 26296 22140 26327
rect 22664 26296 22692 26472
rect 23845 26469 23857 26472
rect 23891 26469 23903 26503
rect 23845 26463 23903 26469
rect 25041 26503 25099 26509
rect 25041 26469 25053 26503
rect 25087 26500 25099 26503
rect 25222 26500 25228 26512
rect 25087 26472 25228 26500
rect 25087 26469 25099 26472
rect 25041 26463 25099 26469
rect 25222 26460 25228 26472
rect 25280 26460 25286 26512
rect 25314 26460 25320 26512
rect 25372 26460 25378 26512
rect 26068 26500 26096 26540
rect 26510 26528 26516 26540
rect 26568 26528 26574 26580
rect 27338 26568 27344 26580
rect 26620 26540 27344 26568
rect 26620 26500 26648 26540
rect 27338 26528 27344 26540
rect 27396 26528 27402 26580
rect 27433 26571 27491 26577
rect 27433 26537 27445 26571
rect 27479 26568 27491 26571
rect 29822 26568 29828 26580
rect 27479 26540 29828 26568
rect 27479 26537 27491 26540
rect 27433 26531 27491 26537
rect 29822 26528 29828 26540
rect 29880 26528 29886 26580
rect 45462 26528 45468 26580
rect 45520 26568 45526 26580
rect 45520 26528 45554 26568
rect 45646 26528 45652 26580
rect 45704 26568 45710 26580
rect 45704 26540 45749 26568
rect 45704 26528 45710 26540
rect 26068 26472 26648 26500
rect 27062 26460 27068 26512
rect 27120 26460 27126 26512
rect 27617 26503 27675 26509
rect 27617 26469 27629 26503
rect 27663 26469 27675 26503
rect 27617 26463 27675 26469
rect 27080 26432 27108 26460
rect 27632 26432 27660 26463
rect 27798 26460 27804 26512
rect 27856 26500 27862 26512
rect 28718 26500 28724 26512
rect 27856 26472 28724 26500
rect 27856 26460 27862 26472
rect 28718 26460 28724 26472
rect 28776 26500 28782 26512
rect 29733 26503 29791 26509
rect 29733 26500 29745 26503
rect 28776 26472 29745 26500
rect 28776 26460 28782 26472
rect 29733 26469 29745 26472
rect 29779 26469 29791 26503
rect 29733 26463 29791 26469
rect 30282 26460 30288 26512
rect 30340 26500 30346 26512
rect 31757 26503 31815 26509
rect 31757 26500 31769 26503
rect 30340 26472 31769 26500
rect 30340 26460 30346 26472
rect 31757 26469 31769 26472
rect 31803 26469 31815 26503
rect 31757 26463 31815 26469
rect 31938 26460 31944 26512
rect 31996 26500 32002 26512
rect 45526 26500 45554 26528
rect 47578 26500 47584 26512
rect 31996 26472 33456 26500
rect 45526 26472 47584 26500
rect 31996 26460 32002 26472
rect 30466 26432 30472 26444
rect 23492 26404 24900 26432
rect 23492 26305 23520 26404
rect 24872 26376 24900 26404
rect 26436 26404 27660 26432
rect 28368 26404 30472 26432
rect 24670 26364 24676 26376
rect 24631 26336 24676 26364
rect 24670 26324 24676 26336
rect 24728 26324 24734 26376
rect 24854 26364 24860 26376
rect 24815 26336 24860 26364
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 26436 26373 26464 26404
rect 26421 26367 26479 26373
rect 26421 26333 26433 26367
rect 26467 26333 26479 26367
rect 26421 26327 26479 26333
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26364 27123 26367
rect 27154 26364 27160 26376
rect 27111 26336 27160 26364
rect 27111 26333 27123 26336
rect 27065 26327 27123 26333
rect 27154 26324 27160 26336
rect 27212 26324 27218 26376
rect 27430 26364 27436 26376
rect 27391 26336 27436 26364
rect 27430 26324 27436 26336
rect 27488 26324 27494 26376
rect 27614 26324 27620 26376
rect 27672 26364 27678 26376
rect 28368 26373 28396 26404
rect 30466 26392 30472 26404
rect 30524 26392 30530 26444
rect 32122 26432 32128 26444
rect 31726 26404 32128 26432
rect 28353 26367 28411 26373
rect 28353 26364 28365 26367
rect 27672 26336 28365 26364
rect 27672 26324 27678 26336
rect 28353 26333 28365 26336
rect 28399 26333 28411 26367
rect 28353 26327 28411 26333
rect 28534 26324 28540 26376
rect 28592 26364 28598 26376
rect 29549 26367 29607 26373
rect 29549 26364 29561 26367
rect 28592 26336 29561 26364
rect 28592 26324 28598 26336
rect 29549 26333 29561 26336
rect 29595 26364 29607 26367
rect 31330 26367 31388 26373
rect 31330 26364 31342 26367
rect 29595 26336 31342 26364
rect 29595 26333 29607 26336
rect 29549 26327 29607 26333
rect 31330 26333 31342 26336
rect 31376 26364 31388 26367
rect 31726 26364 31754 26404
rect 32122 26392 32128 26404
rect 32180 26392 32186 26444
rect 32309 26435 32367 26441
rect 32309 26401 32321 26435
rect 32355 26432 32367 26435
rect 33318 26432 33324 26444
rect 32355 26404 33324 26432
rect 32355 26401 32367 26404
rect 32309 26395 32367 26401
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 31846 26364 31852 26376
rect 31376 26336 31754 26364
rect 31807 26336 31852 26364
rect 31376 26333 31388 26336
rect 31330 26327 31388 26333
rect 31846 26324 31852 26336
rect 31904 26324 31910 26376
rect 32493 26367 32551 26373
rect 32493 26333 32505 26367
rect 32539 26333 32551 26367
rect 32493 26327 32551 26333
rect 21692 26268 22692 26296
rect 23477 26299 23535 26305
rect 21692 26256 21698 26268
rect 23477 26265 23489 26299
rect 23523 26265 23535 26299
rect 23477 26259 23535 26265
rect 23661 26299 23719 26305
rect 23661 26265 23673 26299
rect 23707 26296 23719 26299
rect 23750 26296 23756 26308
rect 23707 26268 23756 26296
rect 23707 26265 23719 26268
rect 23661 26259 23719 26265
rect 23750 26256 23756 26268
rect 23808 26296 23814 26308
rect 24397 26299 24455 26305
rect 24397 26296 24409 26299
rect 23808 26268 24409 26296
rect 23808 26256 23814 26268
rect 24397 26265 24409 26268
rect 24443 26265 24455 26299
rect 24688 26296 24716 26324
rect 25038 26296 25044 26308
rect 24688 26268 25044 26296
rect 24397 26259 24455 26265
rect 25038 26256 25044 26268
rect 25096 26256 25102 26308
rect 28169 26299 28227 26305
rect 28169 26265 28181 26299
rect 28215 26296 28227 26299
rect 28626 26296 28632 26308
rect 28215 26268 28632 26296
rect 28215 26265 28227 26268
rect 28169 26259 28227 26265
rect 21450 26228 21456 26240
rect 19306 26200 21456 26228
rect 14921 26191 14979 26197
rect 21450 26188 21456 26200
rect 21508 26188 21514 26240
rect 23290 26188 23296 26240
rect 23348 26228 23354 26240
rect 25406 26228 25412 26240
rect 23348 26200 25412 26228
rect 23348 26188 23354 26200
rect 25406 26188 25412 26200
rect 25464 26188 25470 26240
rect 26510 26188 26516 26240
rect 26568 26228 26574 26240
rect 28184 26228 28212 26259
rect 28626 26256 28632 26268
rect 28684 26256 28690 26308
rect 32508 26296 32536 26327
rect 32582 26324 32588 26376
rect 32640 26364 32646 26376
rect 32766 26364 32772 26376
rect 32640 26336 32685 26364
rect 32727 26336 32772 26364
rect 32640 26324 32646 26336
rect 32766 26324 32772 26336
rect 32824 26324 32830 26376
rect 32858 26324 32864 26376
rect 32916 26364 32922 26376
rect 33428 26373 33456 26472
rect 47578 26460 47584 26472
rect 47636 26460 47642 26512
rect 33781 26435 33839 26441
rect 33781 26401 33793 26435
rect 33827 26432 33839 26435
rect 40126 26432 40132 26444
rect 33827 26404 40132 26432
rect 33827 26401 33839 26404
rect 33781 26395 33839 26401
rect 40126 26392 40132 26404
rect 40184 26392 40190 26444
rect 45646 26432 45652 26444
rect 43548 26404 45652 26432
rect 33413 26367 33471 26373
rect 32916 26336 32961 26364
rect 32916 26324 32922 26336
rect 33413 26333 33425 26367
rect 33459 26333 33471 26367
rect 33413 26327 33471 26333
rect 33502 26324 33508 26376
rect 33560 26364 33566 26376
rect 33601 26367 33659 26373
rect 33601 26364 33613 26367
rect 33560 26336 33613 26364
rect 33560 26324 33566 26336
rect 33601 26333 33613 26336
rect 33647 26333 33659 26367
rect 33601 26327 33659 26333
rect 33698 26367 33756 26373
rect 33698 26333 33710 26367
rect 33744 26333 33756 26367
rect 33962 26364 33968 26376
rect 33923 26336 33968 26364
rect 33698 26327 33756 26333
rect 31404 26268 32536 26296
rect 31404 26240 31432 26268
rect 33226 26256 33232 26308
rect 33284 26296 33290 26308
rect 33713 26296 33741 26327
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 43548 26373 43576 26404
rect 45646 26392 45652 26404
rect 45704 26392 45710 26444
rect 47302 26432 47308 26444
rect 45940 26404 47308 26432
rect 43533 26367 43591 26373
rect 43533 26333 43545 26367
rect 43579 26333 43591 26367
rect 43533 26327 43591 26333
rect 43990 26324 43996 26376
rect 44048 26364 44054 26376
rect 44269 26367 44327 26373
rect 44269 26364 44281 26367
rect 44048 26336 44281 26364
rect 44048 26324 44054 26336
rect 44269 26333 44281 26336
rect 44315 26333 44327 26367
rect 45462 26364 45468 26376
rect 45423 26336 45468 26364
rect 44269 26327 44327 26333
rect 34146 26296 34152 26308
rect 33284 26268 33741 26296
rect 34107 26268 34152 26296
rect 33284 26256 33290 26268
rect 34146 26256 34152 26268
rect 34204 26256 34210 26308
rect 44284 26296 44312 26327
rect 45462 26324 45468 26336
rect 45520 26324 45526 26376
rect 45940 26296 45968 26404
rect 47302 26392 47308 26404
rect 47360 26392 47366 26444
rect 46014 26324 46020 26376
rect 46072 26364 46078 26376
rect 46293 26367 46351 26373
rect 46293 26364 46305 26367
rect 46072 26336 46305 26364
rect 46072 26324 46078 26336
rect 46293 26333 46305 26336
rect 46339 26333 46351 26367
rect 46293 26327 46351 26333
rect 44284 26268 45968 26296
rect 46477 26299 46535 26305
rect 46477 26265 46489 26299
rect 46523 26296 46535 26299
rect 47670 26296 47676 26308
rect 46523 26268 47676 26296
rect 46523 26265 46535 26268
rect 46477 26259 46535 26265
rect 47670 26256 47676 26268
rect 47728 26256 47734 26308
rect 48130 26296 48136 26308
rect 48091 26268 48136 26296
rect 48130 26256 48136 26268
rect 48188 26256 48194 26308
rect 26568 26200 28212 26228
rect 26568 26188 26574 26200
rect 30926 26188 30932 26240
rect 30984 26228 30990 26240
rect 31205 26231 31263 26237
rect 31205 26228 31217 26231
rect 30984 26200 31217 26228
rect 30984 26188 30990 26200
rect 31205 26197 31217 26200
rect 31251 26197 31263 26231
rect 31386 26228 31392 26240
rect 31347 26200 31392 26228
rect 31205 26191 31263 26197
rect 31386 26188 31392 26200
rect 31444 26188 31450 26240
rect 31478 26188 31484 26240
rect 31536 26228 31542 26240
rect 36538 26228 36544 26240
rect 31536 26200 36544 26228
rect 31536 26188 31542 26200
rect 36538 26188 36544 26200
rect 36596 26188 36602 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 2314 25984 2320 26036
rect 2372 26024 2378 26036
rect 13449 26027 13507 26033
rect 2372 25996 13400 26024
rect 2372 25984 2378 25996
rect 11514 25956 11520 25968
rect 11427 25928 11520 25956
rect 11514 25916 11520 25928
rect 11572 25956 11578 25968
rect 13078 25956 13084 25968
rect 11572 25928 13084 25956
rect 11572 25916 11578 25928
rect 13078 25916 13084 25928
rect 13136 25916 13142 25968
rect 13281 25959 13339 25965
rect 13281 25956 13293 25959
rect 13280 25925 13293 25956
rect 13327 25925 13339 25959
rect 13372 25956 13400 25996
rect 13449 25993 13461 26027
rect 13495 26024 13507 26027
rect 14826 26024 14832 26036
rect 13495 25996 14832 26024
rect 13495 25993 13507 25996
rect 13449 25987 13507 25993
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 15194 25984 15200 26036
rect 15252 26024 15258 26036
rect 15289 26027 15347 26033
rect 15289 26024 15301 26027
rect 15252 25996 15301 26024
rect 15252 25984 15258 25996
rect 15289 25993 15301 25996
rect 15335 26024 15347 26027
rect 15470 26024 15476 26036
rect 15335 25996 15476 26024
rect 15335 25993 15347 25996
rect 15289 25987 15347 25993
rect 15470 25984 15476 25996
rect 15528 25984 15534 26036
rect 15654 25984 15660 26036
rect 15712 26024 15718 26036
rect 16025 26027 16083 26033
rect 16025 26024 16037 26027
rect 15712 25996 16037 26024
rect 15712 25984 15718 25996
rect 16025 25993 16037 25996
rect 16071 25993 16083 26027
rect 16025 25987 16083 25993
rect 17402 25984 17408 26036
rect 17460 26024 17466 26036
rect 18782 26024 18788 26036
rect 17460 25996 18276 26024
rect 18743 25996 18788 26024
rect 17460 25984 17466 25996
rect 13372 25928 18184 25956
rect 13280 25919 13339 25925
rect 10137 25891 10195 25897
rect 10137 25857 10149 25891
rect 10183 25857 10195 25891
rect 10137 25851 10195 25857
rect 10152 25820 10180 25851
rect 11422 25848 11428 25900
rect 11480 25888 11486 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 11480 25860 11713 25888
rect 11480 25848 11486 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 11793 25891 11851 25897
rect 11793 25857 11805 25891
rect 11839 25888 11851 25891
rect 12066 25888 12072 25900
rect 11839 25860 12072 25888
rect 11839 25857 11851 25860
rect 11793 25851 11851 25857
rect 12066 25848 12072 25860
rect 12124 25848 12130 25900
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25888 12311 25891
rect 13170 25888 13176 25900
rect 12299 25860 13176 25888
rect 12299 25857 12311 25860
rect 12253 25851 12311 25857
rect 13170 25848 13176 25860
rect 13228 25848 13234 25900
rect 10778 25820 10784 25832
rect 10152 25792 10784 25820
rect 10778 25780 10784 25792
rect 10836 25820 10842 25832
rect 13280 25820 13308 25919
rect 14277 25891 14335 25897
rect 14277 25857 14289 25891
rect 14323 25888 14335 25891
rect 14642 25888 14648 25900
rect 14323 25860 14648 25888
rect 14323 25857 14335 25860
rect 14277 25851 14335 25857
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 15102 25848 15108 25900
rect 15160 25888 15166 25900
rect 15160 25860 15205 25888
rect 15160 25848 15166 25860
rect 15562 25848 15568 25900
rect 15620 25888 15626 25900
rect 15841 25891 15899 25897
rect 15841 25888 15853 25891
rect 15620 25860 15853 25888
rect 15620 25848 15626 25860
rect 15841 25857 15853 25860
rect 15887 25888 15899 25891
rect 16114 25888 16120 25900
rect 15887 25860 16120 25888
rect 15887 25857 15899 25860
rect 15841 25851 15899 25857
rect 16114 25848 16120 25860
rect 16172 25848 16178 25900
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 18049 25891 18107 25897
rect 18049 25857 18061 25891
rect 18095 25857 18107 25891
rect 18049 25851 18107 25857
rect 14366 25820 14372 25832
rect 10836 25792 12480 25820
rect 13280 25792 14372 25820
rect 10836 25780 10842 25792
rect 9674 25712 9680 25764
rect 9732 25752 9738 25764
rect 9732 25724 10364 25752
rect 9732 25712 9738 25724
rect 9858 25644 9864 25696
rect 9916 25684 9922 25696
rect 10229 25687 10287 25693
rect 10229 25684 10241 25687
rect 9916 25656 10241 25684
rect 9916 25644 9922 25656
rect 10229 25653 10241 25656
rect 10275 25653 10287 25687
rect 10336 25684 10364 25724
rect 11054 25712 11060 25764
rect 11112 25752 11118 25764
rect 12452 25761 12480 25792
rect 14366 25780 14372 25792
rect 14424 25780 14430 25832
rect 11517 25755 11575 25761
rect 11517 25752 11529 25755
rect 11112 25724 11529 25752
rect 11112 25712 11118 25724
rect 11517 25721 11529 25724
rect 11563 25721 11575 25755
rect 11517 25715 11575 25721
rect 12437 25755 12495 25761
rect 12437 25721 12449 25755
rect 12483 25721 12495 25755
rect 14461 25755 14519 25761
rect 14461 25752 14473 25755
rect 12437 25715 12495 25721
rect 13096 25724 14473 25752
rect 13096 25684 13124 25724
rect 14461 25721 14473 25724
rect 14507 25721 14519 25755
rect 14461 25715 14519 25721
rect 15010 25712 15016 25764
rect 15068 25752 15074 25764
rect 17052 25752 17080 25851
rect 15068 25724 17080 25752
rect 18064 25752 18092 25851
rect 18156 25820 18184 25928
rect 18248 25888 18276 25996
rect 18782 25984 18788 25996
rect 18840 25984 18846 26036
rect 20714 26024 20720 26036
rect 20675 25996 20720 26024
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 26050 26024 26056 26036
rect 23676 25996 26056 26024
rect 18693 25891 18751 25897
rect 18693 25888 18705 25891
rect 18248 25860 18705 25888
rect 18693 25857 18705 25860
rect 18739 25857 18751 25891
rect 20622 25888 20628 25900
rect 20583 25860 20628 25888
rect 18693 25851 18751 25857
rect 20622 25848 20628 25860
rect 20680 25888 20686 25900
rect 22186 25888 22192 25900
rect 20680 25860 22192 25888
rect 20680 25848 20686 25860
rect 22186 25848 22192 25860
rect 22244 25848 22250 25900
rect 23017 25891 23075 25897
rect 23017 25857 23029 25891
rect 23063 25888 23075 25891
rect 23063 25860 23520 25888
rect 23063 25857 23075 25860
rect 23017 25851 23075 25857
rect 18156 25792 23428 25820
rect 23290 25752 23296 25764
rect 18064 25724 23296 25752
rect 15068 25712 15074 25724
rect 23290 25712 23296 25724
rect 23348 25712 23354 25764
rect 13262 25684 13268 25696
rect 10336 25656 13124 25684
rect 13223 25656 13268 25684
rect 10229 25647 10287 25653
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 17221 25687 17279 25693
rect 17221 25653 17233 25687
rect 17267 25684 17279 25687
rect 17402 25684 17408 25696
rect 17267 25656 17408 25684
rect 17267 25653 17279 25656
rect 17221 25647 17279 25653
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 18138 25684 18144 25696
rect 18099 25656 18144 25684
rect 18138 25644 18144 25656
rect 18196 25644 18202 25696
rect 22370 25644 22376 25696
rect 22428 25684 22434 25696
rect 22833 25687 22891 25693
rect 22833 25684 22845 25687
rect 22428 25656 22845 25684
rect 22428 25644 22434 25656
rect 22833 25653 22845 25656
rect 22879 25653 22891 25687
rect 23400 25684 23428 25792
rect 23492 25761 23520 25860
rect 23676 25820 23704 25996
rect 26050 25984 26056 25996
rect 26108 25984 26114 26036
rect 26145 26027 26203 26033
rect 26145 25993 26157 26027
rect 26191 26024 26203 26027
rect 26602 26024 26608 26036
rect 26191 25996 26608 26024
rect 26191 25993 26203 25996
rect 26145 25987 26203 25993
rect 26602 25984 26608 25996
rect 26660 25984 26666 26036
rect 26973 26027 27031 26033
rect 26973 25993 26985 26027
rect 27019 25993 27031 26027
rect 26973 25987 27031 25993
rect 27341 26027 27399 26033
rect 27341 25993 27353 26027
rect 27387 26024 27399 26027
rect 28534 26024 28540 26036
rect 27387 25996 28540 26024
rect 27387 25993 27399 25996
rect 27341 25987 27399 25993
rect 23750 25916 23756 25968
rect 23808 25956 23814 25968
rect 26988 25956 27016 25987
rect 28534 25984 28540 25996
rect 28592 25984 28598 26036
rect 28813 26027 28871 26033
rect 28813 25993 28825 26027
rect 28859 26024 28871 26027
rect 31938 26024 31944 26036
rect 28859 25996 31944 26024
rect 28859 25993 28871 25996
rect 28813 25987 28871 25993
rect 31938 25984 31944 25996
rect 31996 25984 32002 26036
rect 32030 25984 32036 26036
rect 32088 26024 32094 26036
rect 32088 25996 33916 26024
rect 32088 25984 32094 25996
rect 23808 25928 25176 25956
rect 23808 25916 23814 25928
rect 23842 25888 23848 25900
rect 23803 25860 23848 25888
rect 23842 25848 23848 25860
rect 23900 25848 23906 25900
rect 23937 25891 23995 25897
rect 23937 25857 23949 25891
rect 23983 25888 23995 25891
rect 24673 25891 24731 25897
rect 24673 25888 24685 25891
rect 23983 25860 24685 25888
rect 23983 25857 23995 25860
rect 23937 25851 23995 25857
rect 24673 25857 24685 25860
rect 24719 25857 24731 25891
rect 24854 25888 24860 25900
rect 24815 25860 24860 25888
rect 24673 25851 24731 25857
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 25038 25888 25044 25900
rect 24999 25860 25044 25888
rect 25038 25848 25044 25860
rect 25096 25848 25102 25900
rect 25148 25897 25176 25928
rect 25976 25928 27016 25956
rect 25976 25897 26004 25928
rect 27890 25916 27896 25968
rect 27948 25956 27954 25968
rect 31478 25956 31484 25968
rect 27948 25928 31484 25956
rect 27948 25916 27954 25928
rect 31478 25916 31484 25928
rect 31536 25916 31542 25968
rect 25133 25891 25191 25897
rect 25133 25857 25145 25891
rect 25179 25857 25191 25891
rect 25133 25851 25191 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 25961 25851 26019 25857
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 24029 25823 24087 25829
rect 24029 25820 24041 25823
rect 23676 25792 24041 25820
rect 24029 25789 24041 25792
rect 24075 25789 24087 25823
rect 26252 25820 26280 25851
rect 26786 25848 26792 25900
rect 26844 25888 26850 25900
rect 28261 25891 28319 25897
rect 26844 25860 27752 25888
rect 26844 25848 26850 25860
rect 27448 25832 27476 25860
rect 27430 25820 27436 25832
rect 24029 25783 24087 25789
rect 24136 25792 26280 25820
rect 27391 25792 27436 25820
rect 23477 25755 23535 25761
rect 23477 25721 23489 25755
rect 23523 25721 23535 25755
rect 23477 25715 23535 25721
rect 24136 25684 24164 25792
rect 27430 25780 27436 25792
rect 27488 25780 27494 25832
rect 27614 25820 27620 25832
rect 27575 25792 27620 25820
rect 27614 25780 27620 25792
rect 27672 25780 27678 25832
rect 27724 25820 27752 25860
rect 28261 25857 28273 25891
rect 28307 25888 28319 25891
rect 28442 25888 28448 25900
rect 28307 25860 28448 25888
rect 28307 25857 28319 25860
rect 28261 25851 28319 25857
rect 28442 25848 28448 25860
rect 28500 25848 28506 25900
rect 28626 25888 28632 25900
rect 28587 25860 28632 25888
rect 28626 25848 28632 25860
rect 28684 25848 28690 25900
rect 29546 25888 29552 25900
rect 29507 25860 29552 25888
rect 29546 25848 29552 25860
rect 29604 25848 29610 25900
rect 30834 25888 30840 25900
rect 30795 25860 30840 25888
rect 30834 25848 30840 25860
rect 30892 25848 30898 25900
rect 30926 25848 30932 25900
rect 30984 25888 30990 25900
rect 31202 25888 31208 25900
rect 30984 25860 31029 25888
rect 31163 25860 31208 25888
rect 30984 25848 30990 25860
rect 31202 25848 31208 25860
rect 31260 25848 31266 25900
rect 32140 25897 32168 25996
rect 32858 25916 32864 25968
rect 32916 25916 32922 25968
rect 33888 25900 33916 25996
rect 36538 25984 36544 26036
rect 36596 26024 36602 26036
rect 45830 26024 45836 26036
rect 36596 25996 45836 26024
rect 36596 25984 36602 25996
rect 45830 25984 45836 25996
rect 45888 25984 45894 26036
rect 34698 25956 34704 25968
rect 34348 25928 34704 25956
rect 32125 25891 32183 25897
rect 32125 25857 32137 25891
rect 32171 25857 32183 25891
rect 32125 25851 32183 25857
rect 33870 25848 33876 25900
rect 33928 25888 33934 25900
rect 34348 25897 34376 25928
rect 34698 25916 34704 25928
rect 34756 25916 34762 25968
rect 35342 25916 35348 25968
rect 35400 25916 35406 25968
rect 45373 25959 45431 25965
rect 45373 25925 45385 25959
rect 45419 25956 45431 25959
rect 45738 25956 45744 25968
rect 45419 25928 45744 25956
rect 45419 25925 45431 25928
rect 45373 25919 45431 25925
rect 45738 25916 45744 25928
rect 45796 25916 45802 25968
rect 45922 25916 45928 25968
rect 45980 25956 45986 25968
rect 45980 25928 47624 25956
rect 45980 25916 45986 25928
rect 47596 25897 47624 25928
rect 34333 25891 34391 25897
rect 34333 25888 34345 25891
rect 33928 25860 34345 25888
rect 33928 25848 33934 25860
rect 34333 25857 34345 25860
rect 34379 25857 34391 25891
rect 34333 25851 34391 25857
rect 47581 25891 47639 25897
rect 47581 25857 47593 25891
rect 47627 25857 47639 25891
rect 47581 25851 47639 25857
rect 29733 25823 29791 25829
rect 29733 25820 29745 25823
rect 27724 25792 29745 25820
rect 29733 25789 29745 25792
rect 29779 25820 29791 25823
rect 30098 25820 30104 25832
rect 29779 25792 30104 25820
rect 29779 25789 29791 25792
rect 29733 25783 29791 25789
rect 30098 25780 30104 25792
rect 30156 25780 30162 25832
rect 30653 25823 30711 25829
rect 30653 25789 30665 25823
rect 30699 25820 30711 25823
rect 32401 25823 32459 25829
rect 32401 25820 32413 25823
rect 30699 25792 32413 25820
rect 30699 25789 30711 25792
rect 30653 25783 30711 25789
rect 32401 25789 32413 25792
rect 32447 25789 32459 25823
rect 32401 25783 32459 25789
rect 32766 25780 32772 25832
rect 32824 25820 32830 25832
rect 34606 25820 34612 25832
rect 32824 25792 33916 25820
rect 34567 25792 34612 25820
rect 32824 25780 32830 25792
rect 24949 25755 25007 25761
rect 24949 25721 24961 25755
rect 24995 25752 25007 25755
rect 25314 25752 25320 25764
rect 24995 25724 25320 25752
rect 24995 25721 25007 25724
rect 24949 25715 25007 25721
rect 25314 25712 25320 25724
rect 25372 25712 25378 25764
rect 26602 25712 26608 25764
rect 26660 25752 26666 25764
rect 32122 25752 32128 25764
rect 26660 25724 32128 25752
rect 26660 25712 26666 25724
rect 32122 25712 32128 25724
rect 32180 25712 32186 25764
rect 33888 25761 33916 25792
rect 34606 25780 34612 25792
rect 34664 25780 34670 25832
rect 45186 25820 45192 25832
rect 45147 25792 45192 25820
rect 45186 25780 45192 25792
rect 45244 25780 45250 25832
rect 46842 25820 46848 25832
rect 46803 25792 46848 25820
rect 46842 25780 46848 25792
rect 46900 25780 46906 25832
rect 33873 25755 33931 25761
rect 33873 25721 33885 25755
rect 33919 25721 33931 25755
rect 33873 25715 33931 25721
rect 23400 25656 24164 25684
rect 25777 25687 25835 25693
rect 22833 25647 22891 25653
rect 25777 25653 25789 25687
rect 25823 25684 25835 25687
rect 25866 25684 25872 25696
rect 25823 25656 25872 25684
rect 25823 25653 25835 25656
rect 25777 25647 25835 25653
rect 25866 25644 25872 25656
rect 25924 25644 25930 25696
rect 28350 25684 28356 25696
rect 28311 25656 28356 25684
rect 28350 25644 28356 25656
rect 28408 25644 28414 25696
rect 31113 25687 31171 25693
rect 31113 25653 31125 25687
rect 31159 25684 31171 25687
rect 31294 25684 31300 25696
rect 31159 25656 31300 25684
rect 31159 25653 31171 25656
rect 31113 25647 31171 25653
rect 31294 25644 31300 25656
rect 31352 25644 31358 25696
rect 31478 25644 31484 25696
rect 31536 25684 31542 25696
rect 33778 25684 33784 25696
rect 31536 25656 33784 25684
rect 31536 25644 31542 25656
rect 33778 25644 33784 25656
rect 33836 25644 33842 25696
rect 36078 25684 36084 25696
rect 36039 25656 36084 25684
rect 36078 25644 36084 25656
rect 36136 25644 36142 25696
rect 46290 25644 46296 25696
rect 46348 25684 46354 25696
rect 47673 25687 47731 25693
rect 47673 25684 47685 25687
rect 46348 25656 47685 25684
rect 46348 25644 46354 25656
rect 47673 25653 47685 25656
rect 47719 25653 47731 25687
rect 47673 25647 47731 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 11422 25440 11428 25492
rect 11480 25480 11486 25492
rect 13262 25480 13268 25492
rect 11480 25452 13268 25480
rect 11480 25440 11486 25452
rect 13262 25440 13268 25452
rect 13320 25440 13326 25492
rect 14277 25483 14335 25489
rect 14277 25449 14289 25483
rect 14323 25480 14335 25483
rect 14366 25480 14372 25492
rect 14323 25452 14372 25480
rect 14323 25449 14335 25452
rect 14277 25443 14335 25449
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 15105 25483 15163 25489
rect 15105 25449 15117 25483
rect 15151 25480 15163 25483
rect 15562 25480 15568 25492
rect 15151 25452 15568 25480
rect 15151 25449 15163 25452
rect 15105 25443 15163 25449
rect 15562 25440 15568 25452
rect 15620 25440 15626 25492
rect 15657 25483 15715 25489
rect 15657 25449 15669 25483
rect 15703 25480 15715 25483
rect 15930 25480 15936 25492
rect 15703 25452 15936 25480
rect 15703 25449 15715 25452
rect 15657 25443 15715 25449
rect 15930 25440 15936 25452
rect 15988 25440 15994 25492
rect 17586 25480 17592 25492
rect 17547 25452 17592 25480
rect 17586 25440 17592 25452
rect 17644 25440 17650 25492
rect 23750 25440 23756 25492
rect 23808 25480 23814 25492
rect 23845 25483 23903 25489
rect 23845 25480 23857 25483
rect 23808 25452 23857 25480
rect 23808 25440 23814 25452
rect 23845 25449 23857 25452
rect 23891 25449 23903 25483
rect 26602 25480 26608 25492
rect 26563 25452 26608 25480
rect 23845 25443 23903 25449
rect 26602 25440 26608 25452
rect 26660 25440 26666 25492
rect 28074 25440 28080 25492
rect 28132 25480 28138 25492
rect 28905 25483 28963 25489
rect 28905 25480 28917 25483
rect 28132 25452 28917 25480
rect 28132 25440 28138 25452
rect 28905 25449 28917 25452
rect 28951 25449 28963 25483
rect 28905 25443 28963 25449
rect 28994 25440 29000 25492
rect 29052 25480 29058 25492
rect 31202 25480 31208 25492
rect 29052 25452 31208 25480
rect 29052 25440 29058 25452
rect 31202 25440 31208 25452
rect 31260 25440 31266 25492
rect 31386 25480 31392 25492
rect 31347 25452 31392 25480
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 31846 25440 31852 25492
rect 31904 25480 31910 25492
rect 32125 25483 32183 25489
rect 32125 25480 32137 25483
rect 31904 25452 32137 25480
rect 31904 25440 31910 25452
rect 32125 25449 32137 25452
rect 32171 25480 32183 25483
rect 32858 25480 32864 25492
rect 32171 25452 32444 25480
rect 32819 25452 32864 25480
rect 32171 25449 32183 25452
rect 32125 25443 32183 25449
rect 9858 25344 9864 25356
rect 9819 25316 9864 25344
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 15102 25344 15108 25356
rect 14108 25316 15108 25344
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25276 12127 25279
rect 12526 25276 12532 25288
rect 12115 25248 12532 25276
rect 12115 25245 12127 25248
rect 12069 25239 12127 25245
rect 12526 25236 12532 25248
rect 12584 25236 12590 25288
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 10134 25208 10140 25220
rect 10095 25180 10140 25208
rect 10134 25168 10140 25180
rect 10192 25168 10198 25220
rect 14108 25217 14136 25316
rect 15102 25304 15108 25316
rect 15160 25344 15166 25356
rect 19242 25344 19248 25356
rect 15160 25316 19248 25344
rect 15160 25304 15166 25316
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 22370 25344 22376 25356
rect 22331 25316 22376 25344
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 26620 25344 26648 25440
rect 29730 25372 29736 25424
rect 29788 25412 29794 25424
rect 32309 25415 32367 25421
rect 32309 25412 32321 25415
rect 29788 25384 32321 25412
rect 29788 25372 29794 25384
rect 32309 25381 32321 25384
rect 32355 25381 32367 25415
rect 32309 25375 32367 25381
rect 32416 25412 32444 25452
rect 32858 25440 32864 25452
rect 32916 25440 32922 25492
rect 34149 25483 34207 25489
rect 34149 25449 34161 25483
rect 34195 25480 34207 25483
rect 34606 25480 34612 25492
rect 34195 25452 34612 25480
rect 34195 25449 34207 25452
rect 34149 25443 34207 25449
rect 34606 25440 34612 25452
rect 34664 25440 34670 25492
rect 34885 25483 34943 25489
rect 34885 25449 34897 25483
rect 34931 25480 34943 25483
rect 35342 25480 35348 25492
rect 34931 25452 35348 25480
rect 34931 25449 34943 25452
rect 34885 25443 34943 25449
rect 35342 25440 35348 25452
rect 35400 25440 35406 25492
rect 44453 25483 44511 25489
rect 44453 25449 44465 25483
rect 44499 25480 44511 25483
rect 46014 25480 46020 25492
rect 44499 25452 46020 25480
rect 44499 25449 44511 25452
rect 44453 25443 44511 25449
rect 46014 25440 46020 25452
rect 46072 25440 46078 25492
rect 32766 25412 32772 25424
rect 32416 25384 32772 25412
rect 25148 25316 26648 25344
rect 14921 25279 14979 25285
rect 14921 25276 14933 25279
rect 14200 25248 14933 25276
rect 12161 25211 12219 25217
rect 12161 25208 12173 25211
rect 11362 25180 12173 25208
rect 12161 25177 12173 25180
rect 12207 25177 12219 25211
rect 12161 25171 12219 25177
rect 14093 25211 14151 25217
rect 14093 25177 14105 25211
rect 14139 25177 14151 25211
rect 14093 25171 14151 25177
rect 1946 25140 1952 25152
rect 1907 25112 1952 25140
rect 1946 25100 1952 25112
rect 2004 25100 2010 25152
rect 11514 25100 11520 25152
rect 11572 25140 11578 25152
rect 11609 25143 11667 25149
rect 11609 25140 11621 25143
rect 11572 25112 11621 25140
rect 11572 25100 11578 25112
rect 11609 25109 11621 25112
rect 11655 25109 11667 25143
rect 11609 25103 11667 25109
rect 13170 25100 13176 25152
rect 13228 25140 13234 25152
rect 13722 25140 13728 25152
rect 13228 25112 13728 25140
rect 13228 25100 13234 25112
rect 13722 25100 13728 25112
rect 13780 25140 13786 25152
rect 14200 25140 14228 25248
rect 14921 25245 14933 25248
rect 14967 25245 14979 25279
rect 14921 25239 14979 25245
rect 15286 25236 15292 25288
rect 15344 25276 15350 25288
rect 15657 25279 15715 25285
rect 15657 25276 15669 25279
rect 15344 25248 15669 25276
rect 15344 25236 15350 25248
rect 15657 25245 15669 25248
rect 15703 25245 15715 25279
rect 15838 25276 15844 25288
rect 15799 25248 15844 25276
rect 15657 25239 15715 25245
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 17405 25279 17463 25285
rect 17405 25245 17417 25279
rect 17451 25276 17463 25279
rect 18138 25276 18144 25288
rect 17451 25248 18144 25276
rect 17451 25245 17463 25248
rect 17405 25239 17463 25245
rect 14309 25211 14367 25217
rect 14309 25177 14321 25211
rect 14355 25208 14367 25211
rect 14550 25208 14556 25220
rect 14355 25180 14556 25208
rect 14355 25177 14367 25180
rect 14309 25171 14367 25177
rect 14550 25168 14556 25180
rect 14608 25168 14614 25220
rect 14642 25168 14648 25220
rect 14700 25208 14706 25220
rect 17420 25208 17448 25239
rect 18138 25236 18144 25248
rect 18196 25236 18202 25288
rect 20070 25236 20076 25288
rect 20128 25276 20134 25288
rect 22097 25279 22155 25285
rect 22097 25276 22109 25279
rect 20128 25248 22109 25276
rect 20128 25236 20134 25248
rect 22097 25245 22109 25248
rect 22143 25245 22155 25279
rect 22097 25239 22155 25245
rect 24949 25279 25007 25285
rect 24949 25245 24961 25279
rect 24995 25276 25007 25279
rect 25038 25276 25044 25288
rect 24995 25248 25044 25276
rect 24995 25245 25007 25248
rect 24949 25239 25007 25245
rect 14700 25180 17448 25208
rect 14700 25168 14706 25180
rect 14458 25140 14464 25152
rect 13780 25112 14228 25140
rect 14419 25112 14464 25140
rect 13780 25100 13786 25112
rect 14458 25100 14464 25112
rect 14516 25100 14522 25152
rect 22112 25140 22140 25239
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 25148 25285 25176 25316
rect 27154 25304 27160 25356
rect 27212 25344 27218 25356
rect 31478 25344 31484 25356
rect 27212 25316 31484 25344
rect 27212 25304 27218 25316
rect 31478 25304 31484 25316
rect 31536 25304 31542 25356
rect 31754 25304 31760 25356
rect 31812 25344 31818 25356
rect 31941 25347 31999 25353
rect 31941 25344 31953 25347
rect 31812 25316 31953 25344
rect 31812 25304 31818 25316
rect 31941 25313 31953 25316
rect 31987 25313 31999 25347
rect 32416 25344 32444 25384
rect 32766 25372 32772 25384
rect 32824 25372 32830 25424
rect 33778 25372 33784 25424
rect 33836 25412 33842 25424
rect 45186 25412 45192 25424
rect 33836 25384 45192 25412
rect 33836 25372 33842 25384
rect 45186 25372 45192 25384
rect 45244 25372 45250 25424
rect 31941 25307 31999 25313
rect 32048 25316 32444 25344
rect 25133 25279 25191 25285
rect 25133 25245 25145 25279
rect 25179 25245 25191 25279
rect 25133 25239 25191 25245
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25276 25283 25279
rect 25590 25276 25596 25288
rect 25271 25248 25596 25276
rect 25271 25245 25283 25248
rect 25225 25239 25283 25245
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 26418 25276 26424 25288
rect 26379 25248 26424 25276
rect 26418 25236 26424 25248
rect 26476 25236 26482 25288
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25276 28779 25279
rect 29362 25276 29368 25288
rect 28767 25248 29368 25276
rect 28767 25245 28779 25248
rect 28721 25239 28779 25245
rect 29362 25236 29368 25248
rect 29420 25236 29426 25288
rect 29825 25279 29883 25285
rect 29825 25245 29837 25279
rect 29871 25245 29883 25279
rect 29825 25239 29883 25245
rect 22646 25168 22652 25220
rect 22704 25208 22710 25220
rect 22704 25180 22862 25208
rect 22704 25168 22710 25180
rect 25774 25168 25780 25220
rect 25832 25208 25838 25220
rect 27430 25208 27436 25220
rect 25832 25180 27436 25208
rect 25832 25168 25838 25180
rect 27430 25168 27436 25180
rect 27488 25168 27494 25220
rect 29840 25208 29868 25239
rect 29914 25236 29920 25288
rect 29972 25276 29978 25288
rect 30098 25276 30104 25288
rect 29972 25248 30017 25276
rect 30059 25248 30104 25276
rect 29972 25236 29978 25248
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 30193 25279 30251 25285
rect 30193 25245 30205 25279
rect 30239 25276 30251 25279
rect 31110 25276 31116 25288
rect 30239 25248 31116 25276
rect 30239 25245 30251 25248
rect 30193 25239 30251 25245
rect 31110 25236 31116 25248
rect 31168 25236 31174 25288
rect 31205 25279 31263 25285
rect 31205 25245 31217 25279
rect 31251 25276 31263 25279
rect 32048 25276 32076 25316
rect 32582 25304 32588 25356
rect 32640 25344 32646 25356
rect 33689 25347 33747 25353
rect 33689 25344 33701 25347
rect 32640 25316 33701 25344
rect 32640 25304 32646 25316
rect 33689 25313 33701 25316
rect 33735 25344 33747 25347
rect 36078 25344 36084 25356
rect 33735 25316 36084 25344
rect 33735 25313 33747 25316
rect 33689 25307 33747 25313
rect 36078 25304 36084 25316
rect 36136 25304 36142 25356
rect 46290 25344 46296 25356
rect 46251 25316 46296 25344
rect 46290 25304 46296 25316
rect 46348 25304 46354 25356
rect 47946 25344 47952 25356
rect 47907 25316 47952 25344
rect 47946 25304 47952 25316
rect 48004 25304 48010 25356
rect 31251 25248 32076 25276
rect 32125 25279 32183 25285
rect 31251 25245 31263 25248
rect 31205 25239 31263 25245
rect 32125 25245 32137 25279
rect 32171 25276 32183 25279
rect 32600 25276 32628 25304
rect 32766 25276 32772 25288
rect 32171 25248 32628 25276
rect 32727 25248 32772 25276
rect 32171 25245 32183 25248
rect 32125 25239 32183 25245
rect 32766 25236 32772 25248
rect 32824 25236 32830 25288
rect 33318 25236 33324 25288
rect 33376 25276 33382 25288
rect 33413 25279 33471 25285
rect 33413 25276 33425 25279
rect 33376 25248 33425 25276
rect 33376 25236 33382 25248
rect 33413 25245 33425 25248
rect 33459 25245 33471 25279
rect 33413 25239 33471 25245
rect 33502 25236 33508 25288
rect 33560 25276 33566 25288
rect 33597 25279 33655 25285
rect 33597 25276 33609 25279
rect 33560 25248 33609 25276
rect 33560 25236 33566 25248
rect 33597 25245 33609 25248
rect 33643 25245 33655 25279
rect 33597 25239 33655 25245
rect 33778 25236 33784 25288
rect 33836 25276 33842 25288
rect 33836 25248 33881 25276
rect 33836 25236 33842 25248
rect 33962 25236 33968 25288
rect 34020 25276 34026 25288
rect 34020 25248 34065 25276
rect 34020 25236 34026 25248
rect 34698 25236 34704 25288
rect 34756 25276 34762 25288
rect 34793 25279 34851 25285
rect 34793 25276 34805 25279
rect 34756 25248 34805 25276
rect 34756 25236 34762 25248
rect 34793 25245 34805 25248
rect 34839 25245 34851 25279
rect 45462 25276 45468 25288
rect 45423 25248 45468 25276
rect 34793 25239 34851 25245
rect 45462 25236 45468 25248
rect 45520 25236 45526 25288
rect 45922 25236 45928 25288
rect 45980 25276 45986 25288
rect 46109 25279 46167 25285
rect 46109 25276 46121 25279
rect 45980 25248 46121 25276
rect 45980 25236 45986 25248
rect 46109 25245 46121 25248
rect 46155 25245 46167 25279
rect 46109 25239 46167 25245
rect 31018 25208 31024 25220
rect 29840 25180 30788 25208
rect 30979 25180 31024 25208
rect 22738 25140 22744 25152
rect 22112 25112 22744 25140
rect 22738 25100 22744 25112
rect 22796 25100 22802 25152
rect 24762 25140 24768 25152
rect 24723 25112 24768 25140
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 29641 25143 29699 25149
rect 29641 25109 29653 25143
rect 29687 25140 29699 25143
rect 30466 25140 30472 25152
rect 29687 25112 30472 25140
rect 29687 25109 29699 25112
rect 29641 25103 29699 25109
rect 30466 25100 30472 25112
rect 30524 25100 30530 25152
rect 30760 25140 30788 25180
rect 31018 25168 31024 25180
rect 31076 25168 31082 25220
rect 31846 25208 31852 25220
rect 31312 25180 31524 25208
rect 31807 25180 31852 25208
rect 31312 25140 31340 25180
rect 30760 25112 31340 25140
rect 31496 25140 31524 25180
rect 31846 25168 31852 25180
rect 31904 25168 31910 25220
rect 32214 25140 32220 25152
rect 31496 25112 32220 25140
rect 32214 25100 32220 25112
rect 32272 25100 32278 25152
rect 45554 25100 45560 25152
rect 45612 25140 45618 25152
rect 45612 25112 45657 25140
rect 45612 25100 45618 25112
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 28169 24939 28227 24945
rect 28169 24905 28181 24939
rect 28215 24936 28227 24939
rect 28350 24936 28356 24948
rect 28215 24908 28356 24936
rect 28215 24905 28227 24908
rect 28169 24899 28227 24905
rect 28350 24896 28356 24908
rect 28408 24896 28414 24948
rect 29457 24939 29515 24945
rect 29457 24936 29469 24939
rect 29012 24908 29469 24936
rect 11514 24868 11520 24880
rect 11475 24840 11520 24868
rect 11514 24828 11520 24840
rect 11572 24828 11578 24880
rect 11717 24871 11775 24877
rect 11717 24868 11729 24871
rect 11716 24837 11729 24868
rect 11763 24837 11775 24871
rect 14458 24868 14464 24880
rect 11716 24831 11775 24837
rect 13832 24840 14464 24868
rect 11716 24800 11744 24831
rect 11974 24800 11980 24812
rect 11716 24772 11980 24800
rect 11974 24760 11980 24772
rect 12032 24760 12038 24812
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24800 12495 24803
rect 12710 24800 12716 24812
rect 12483 24772 12716 24800
rect 12483 24769 12495 24772
rect 12437 24763 12495 24769
rect 12710 24760 12716 24772
rect 12768 24800 12774 24812
rect 13832 24800 13860 24840
rect 14458 24828 14464 24840
rect 14516 24828 14522 24880
rect 18064 24840 18460 24868
rect 12768 24772 13860 24800
rect 12768 24760 12774 24772
rect 15838 24760 15844 24812
rect 15896 24800 15902 24812
rect 18064 24800 18092 24840
rect 15896 24772 18092 24800
rect 18141 24803 18199 24809
rect 15896 24760 15902 24772
rect 18141 24769 18153 24803
rect 18187 24769 18199 24803
rect 18322 24800 18328 24812
rect 18283 24772 18328 24800
rect 18141 24763 18199 24769
rect 8570 24732 8576 24744
rect 8531 24704 8576 24732
rect 8570 24692 8576 24704
rect 8628 24692 8634 24744
rect 8757 24735 8815 24741
rect 8757 24701 8769 24735
rect 8803 24732 8815 24735
rect 8938 24732 8944 24744
rect 8803 24704 8944 24732
rect 8803 24701 8815 24704
rect 8757 24695 8815 24701
rect 8938 24692 8944 24704
rect 8996 24692 9002 24744
rect 9033 24735 9091 24741
rect 9033 24701 9045 24735
rect 9079 24701 9091 24735
rect 9033 24695 9091 24701
rect 13817 24735 13875 24741
rect 13817 24701 13829 24735
rect 13863 24701 13875 24735
rect 13817 24695 13875 24701
rect 14001 24735 14059 24741
rect 14001 24701 14013 24735
rect 14047 24732 14059 24735
rect 14182 24732 14188 24744
rect 14047 24704 14188 24732
rect 14047 24701 14059 24704
rect 14001 24695 14059 24701
rect 3602 24556 3608 24608
rect 3660 24596 3666 24608
rect 9048 24596 9076 24695
rect 11422 24624 11428 24676
rect 11480 24664 11486 24676
rect 11885 24667 11943 24673
rect 11885 24664 11897 24667
rect 11480 24636 11897 24664
rect 11480 24624 11486 24636
rect 11885 24633 11897 24636
rect 11931 24633 11943 24667
rect 13832 24664 13860 24695
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14458 24732 14464 24744
rect 14419 24704 14464 24732
rect 14458 24692 14464 24704
rect 14516 24692 14522 24744
rect 18156 24732 18184 24763
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 18432 24809 18460 24840
rect 23474 24828 23480 24880
rect 23532 24828 23538 24880
rect 26418 24828 26424 24880
rect 26476 24868 26482 24880
rect 29012 24868 29040 24908
rect 29457 24905 29469 24908
rect 29503 24936 29515 24939
rect 29914 24936 29920 24948
rect 29503 24908 29920 24936
rect 29503 24905 29515 24908
rect 29457 24899 29515 24905
rect 29914 24896 29920 24908
rect 29972 24896 29978 24948
rect 31018 24896 31024 24948
rect 31076 24936 31082 24948
rect 31389 24939 31447 24945
rect 31389 24936 31401 24939
rect 31076 24908 31401 24936
rect 31076 24896 31082 24908
rect 31389 24905 31401 24908
rect 31435 24905 31447 24939
rect 31389 24899 31447 24905
rect 32214 24896 32220 24948
rect 32272 24936 32278 24948
rect 44082 24936 44088 24948
rect 32272 24908 44088 24936
rect 32272 24896 32278 24908
rect 44082 24896 44088 24908
rect 44140 24896 44146 24948
rect 29362 24868 29368 24880
rect 26476 24840 29040 24868
rect 29323 24840 29368 24868
rect 26476 24828 26482 24840
rect 29362 24828 29368 24840
rect 29420 24868 29426 24880
rect 30374 24868 30380 24880
rect 29420 24840 30380 24868
rect 29420 24828 29426 24840
rect 30374 24828 30380 24840
rect 30432 24868 30438 24880
rect 31205 24871 31263 24877
rect 31205 24868 31217 24871
rect 30432 24840 31217 24868
rect 30432 24828 30438 24840
rect 31205 24837 31217 24840
rect 31251 24837 31263 24871
rect 31205 24831 31263 24837
rect 34790 24828 34796 24880
rect 34848 24828 34854 24880
rect 45020 24840 45876 24868
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24800 18475 24803
rect 19334 24800 19340 24812
rect 18463 24772 19340 24800
rect 18463 24769 18475 24772
rect 18417 24763 18475 24769
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 21266 24800 21272 24812
rect 21227 24772 21272 24800
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 24949 24803 25007 24809
rect 22152 24772 22197 24800
rect 22152 24760 22158 24772
rect 24949 24769 24961 24803
rect 24995 24769 25007 24803
rect 25130 24800 25136 24812
rect 25091 24772 25136 24800
rect 24949 24763 25007 24769
rect 18506 24732 18512 24744
rect 18156 24704 18512 24732
rect 18506 24692 18512 24704
rect 18564 24732 18570 24744
rect 19429 24735 19487 24741
rect 19429 24732 19441 24735
rect 18564 24704 19441 24732
rect 18564 24692 18570 24704
rect 19429 24701 19441 24704
rect 19475 24701 19487 24735
rect 19429 24695 19487 24701
rect 19613 24735 19671 24741
rect 19613 24701 19625 24735
rect 19659 24732 19671 24735
rect 19978 24732 19984 24744
rect 19659 24704 19984 24732
rect 19659 24701 19671 24704
rect 19613 24695 19671 24701
rect 19978 24692 19984 24704
rect 20036 24692 20042 24744
rect 22738 24732 22744 24744
rect 22699 24704 22744 24732
rect 22738 24692 22744 24704
rect 22796 24692 22802 24744
rect 23017 24735 23075 24741
rect 23017 24701 23029 24735
rect 23063 24732 23075 24735
rect 24762 24732 24768 24744
rect 23063 24704 24768 24732
rect 23063 24701 23075 24704
rect 23017 24695 23075 24701
rect 24762 24692 24768 24704
rect 24820 24692 24826 24744
rect 24964 24732 24992 24763
rect 25130 24760 25136 24772
rect 25188 24760 25194 24812
rect 25222 24760 25228 24812
rect 25280 24800 25286 24812
rect 28353 24803 28411 24809
rect 25280 24772 25325 24800
rect 25280 24760 25286 24772
rect 28353 24769 28365 24803
rect 28399 24800 28411 24803
rect 28534 24800 28540 24812
rect 28399 24772 28540 24800
rect 28399 24769 28411 24772
rect 28353 24763 28411 24769
rect 28534 24760 28540 24772
rect 28592 24760 28598 24812
rect 30466 24800 30472 24812
rect 30427 24772 30472 24800
rect 30466 24760 30472 24772
rect 30524 24760 30530 24812
rect 31478 24760 31484 24812
rect 31536 24800 31542 24812
rect 33870 24800 33876 24812
rect 31536 24772 31581 24800
rect 33831 24772 33876 24800
rect 31536 24760 31542 24772
rect 33870 24760 33876 24772
rect 33928 24760 33934 24812
rect 40034 24760 40040 24812
rect 40092 24800 40098 24812
rect 40313 24803 40371 24809
rect 40313 24800 40325 24803
rect 40092 24772 40325 24800
rect 40092 24760 40098 24772
rect 40313 24769 40325 24772
rect 40359 24800 40371 24803
rect 44266 24800 44272 24812
rect 40359 24772 44272 24800
rect 40359 24769 40371 24772
rect 40313 24763 40371 24769
rect 44266 24760 44272 24772
rect 44324 24760 44330 24812
rect 44637 24803 44695 24809
rect 44637 24769 44649 24803
rect 44683 24800 44695 24803
rect 45020 24800 45048 24840
rect 44683 24772 45048 24800
rect 44683 24769 44695 24772
rect 44637 24763 44695 24769
rect 45094 24760 45100 24812
rect 45152 24800 45158 24812
rect 45152 24772 45197 24800
rect 45152 24760 45158 24772
rect 45646 24760 45652 24812
rect 45704 24800 45710 24812
rect 45741 24803 45799 24809
rect 45741 24800 45753 24803
rect 45704 24772 45753 24800
rect 45704 24760 45710 24772
rect 45741 24769 45753 24772
rect 45787 24769 45799 24803
rect 45848 24800 45876 24840
rect 46382 24800 46388 24812
rect 45848 24772 46388 24800
rect 45741 24763 45799 24769
rect 46382 24760 46388 24772
rect 46440 24760 46446 24812
rect 46569 24803 46627 24809
rect 46569 24769 46581 24803
rect 46615 24800 46627 24803
rect 47486 24800 47492 24812
rect 46615 24772 47492 24800
rect 46615 24769 46627 24772
rect 46569 24763 46627 24769
rect 47486 24760 47492 24772
rect 47544 24760 47550 24812
rect 47581 24803 47639 24809
rect 47581 24769 47593 24803
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 28074 24732 28080 24744
rect 24964 24704 28080 24732
rect 28074 24692 28080 24704
rect 28132 24692 28138 24744
rect 28626 24732 28632 24744
rect 28587 24704 28632 24732
rect 28626 24692 28632 24704
rect 28684 24692 28690 24744
rect 30285 24735 30343 24741
rect 30285 24701 30297 24735
rect 30331 24732 30343 24735
rect 30650 24732 30656 24744
rect 30331 24704 30656 24732
rect 30331 24701 30343 24704
rect 30285 24695 30343 24701
rect 30650 24692 30656 24704
rect 30708 24692 30714 24744
rect 30745 24735 30803 24741
rect 30745 24701 30757 24735
rect 30791 24732 30803 24735
rect 31754 24732 31760 24744
rect 30791 24704 31760 24732
rect 30791 24701 30803 24704
rect 30745 24695 30803 24701
rect 31754 24692 31760 24704
rect 31812 24692 31818 24744
rect 34146 24732 34152 24744
rect 34107 24704 34152 24732
rect 34146 24692 34152 24704
rect 34204 24692 34210 24744
rect 46198 24732 46204 24744
rect 35176 24704 46204 24732
rect 13906 24664 13912 24676
rect 13832 24636 13912 24664
rect 11885 24627 11943 24633
rect 13906 24624 13912 24636
rect 13964 24624 13970 24676
rect 16114 24624 16120 24676
rect 16172 24664 16178 24676
rect 22189 24667 22247 24673
rect 16172 24636 22094 24664
rect 16172 24624 16178 24636
rect 11698 24596 11704 24608
rect 3660 24568 9076 24596
rect 11659 24568 11704 24596
rect 3660 24556 3666 24568
rect 11698 24556 11704 24568
rect 11756 24556 11762 24608
rect 12066 24556 12072 24608
rect 12124 24596 12130 24608
rect 12529 24599 12587 24605
rect 12529 24596 12541 24599
rect 12124 24568 12541 24596
rect 12124 24556 12130 24568
rect 12529 24565 12541 24568
rect 12575 24565 12587 24599
rect 12529 24559 12587 24565
rect 17770 24556 17776 24608
rect 17828 24596 17834 24608
rect 18141 24599 18199 24605
rect 18141 24596 18153 24599
rect 17828 24568 18153 24596
rect 17828 24556 17834 24568
rect 18141 24565 18153 24568
rect 18187 24565 18199 24599
rect 22066 24596 22094 24636
rect 22189 24633 22201 24667
rect 22235 24664 22247 24667
rect 22646 24664 22652 24676
rect 22235 24636 22652 24664
rect 22235 24633 22247 24636
rect 22189 24627 22247 24633
rect 22646 24624 22652 24636
rect 22704 24624 22710 24676
rect 24489 24667 24547 24673
rect 24489 24633 24501 24667
rect 24535 24664 24547 24667
rect 24854 24664 24860 24676
rect 24535 24636 24860 24664
rect 24535 24633 24547 24636
rect 24489 24627 24547 24633
rect 24854 24624 24860 24636
rect 24912 24624 24918 24676
rect 24949 24667 25007 24673
rect 24949 24633 24961 24667
rect 24995 24664 25007 24667
rect 25038 24664 25044 24676
rect 24995 24636 25044 24664
rect 24995 24633 25007 24636
rect 24949 24627 25007 24633
rect 25038 24624 25044 24636
rect 25096 24624 25102 24676
rect 27706 24624 27712 24676
rect 27764 24664 27770 24676
rect 27764 24636 31754 24664
rect 27764 24624 27770 24636
rect 25498 24596 25504 24608
rect 22066 24568 25504 24596
rect 18141 24559 18199 24565
rect 25498 24556 25504 24568
rect 25556 24556 25562 24608
rect 27982 24556 27988 24608
rect 28040 24596 28046 24608
rect 28537 24599 28595 24605
rect 28537 24596 28549 24599
rect 28040 24568 28549 24596
rect 28040 24556 28046 24568
rect 28537 24565 28549 24568
rect 28583 24565 28595 24599
rect 28537 24559 28595 24565
rect 29638 24556 29644 24608
rect 29696 24596 29702 24608
rect 30653 24599 30711 24605
rect 30653 24596 30665 24599
rect 29696 24568 30665 24596
rect 29696 24556 29702 24568
rect 30653 24565 30665 24568
rect 30699 24565 30711 24599
rect 30653 24559 30711 24565
rect 31110 24556 31116 24608
rect 31168 24596 31174 24608
rect 31205 24599 31263 24605
rect 31205 24596 31217 24599
rect 31168 24568 31217 24596
rect 31168 24556 31174 24568
rect 31205 24565 31217 24568
rect 31251 24565 31263 24599
rect 31726 24596 31754 24636
rect 35176 24596 35204 24704
rect 46198 24692 46204 24704
rect 46256 24692 46262 24744
rect 47394 24692 47400 24744
rect 47452 24732 47458 24744
rect 47596 24732 47624 24763
rect 47670 24760 47676 24812
rect 47728 24800 47734 24812
rect 47728 24772 47773 24800
rect 47728 24760 47734 24772
rect 47452 24704 47624 24732
rect 47452 24692 47458 24704
rect 44453 24667 44511 24673
rect 44453 24633 44465 24667
rect 44499 24664 44511 24667
rect 45646 24664 45652 24676
rect 44499 24636 45652 24664
rect 44499 24633 44511 24636
rect 44453 24627 44511 24633
rect 45646 24624 45652 24636
rect 45704 24624 45710 24676
rect 35618 24596 35624 24608
rect 31726 24568 35204 24596
rect 35579 24568 35624 24596
rect 31205 24559 31263 24565
rect 35618 24556 35624 24568
rect 35676 24556 35682 24608
rect 40402 24596 40408 24608
rect 40363 24568 40408 24596
rect 40402 24556 40408 24568
rect 40460 24556 40466 24608
rect 45189 24599 45247 24605
rect 45189 24565 45201 24599
rect 45235 24596 45247 24599
rect 46474 24596 46480 24608
rect 45235 24568 46480 24596
rect 45235 24565 45247 24568
rect 45189 24559 45247 24565
rect 46474 24556 46480 24568
rect 46532 24556 46538 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 10134 24352 10140 24404
rect 10192 24392 10198 24404
rect 10505 24395 10563 24401
rect 10505 24392 10517 24395
rect 10192 24364 10517 24392
rect 10192 24352 10198 24364
rect 10505 24361 10517 24364
rect 10551 24361 10563 24395
rect 10505 24355 10563 24361
rect 11974 24352 11980 24404
rect 12032 24392 12038 24404
rect 12713 24395 12771 24401
rect 12713 24392 12725 24395
rect 12032 24364 12725 24392
rect 12032 24352 12038 24364
rect 12713 24361 12725 24364
rect 12759 24361 12771 24395
rect 14182 24392 14188 24404
rect 14143 24364 14188 24392
rect 12713 24355 12771 24361
rect 14182 24352 14188 24364
rect 14240 24352 14246 24404
rect 23385 24395 23443 24401
rect 23385 24361 23397 24395
rect 23431 24392 23443 24395
rect 23474 24392 23480 24404
rect 23431 24364 23480 24392
rect 23431 24361 23443 24364
rect 23385 24355 23443 24361
rect 23474 24352 23480 24364
rect 23532 24352 23538 24404
rect 26602 24352 26608 24404
rect 26660 24392 26666 24404
rect 28537 24395 28595 24401
rect 28537 24392 28549 24395
rect 26660 24364 28549 24392
rect 26660 24352 26666 24364
rect 28537 24361 28549 24364
rect 28583 24392 28595 24395
rect 28626 24392 28632 24404
rect 28583 24364 28632 24392
rect 28583 24361 28595 24364
rect 28537 24355 28595 24361
rect 28626 24352 28632 24364
rect 28684 24352 28690 24404
rect 30193 24395 30251 24401
rect 30193 24361 30205 24395
rect 30239 24392 30251 24395
rect 31478 24392 31484 24404
rect 30239 24364 31484 24392
rect 30239 24361 30251 24364
rect 30193 24355 30251 24361
rect 31478 24352 31484 24364
rect 31536 24352 31542 24404
rect 34790 24392 34796 24404
rect 34751 24364 34796 24392
rect 34790 24352 34796 24364
rect 34848 24352 34854 24404
rect 8570 24284 8576 24336
rect 8628 24324 8634 24336
rect 11057 24327 11115 24333
rect 11057 24324 11069 24327
rect 8628 24296 11069 24324
rect 8628 24284 8634 24296
rect 11057 24293 11069 24296
rect 11103 24324 11115 24327
rect 11514 24324 11520 24336
rect 11103 24296 11520 24324
rect 11103 24293 11115 24296
rect 11057 24287 11115 24293
rect 11514 24284 11520 24296
rect 11572 24284 11578 24336
rect 12897 24327 12955 24333
rect 12897 24324 12909 24327
rect 12406 24296 12909 24324
rect 11149 24259 11207 24265
rect 11149 24225 11161 24259
rect 11195 24256 11207 24259
rect 12406 24256 12434 24296
rect 12897 24293 12909 24296
rect 12943 24293 12955 24327
rect 15838 24324 15844 24336
rect 12897 24287 12955 24293
rect 15120 24296 15844 24324
rect 15120 24265 15148 24296
rect 15838 24284 15844 24296
rect 15896 24284 15902 24336
rect 33226 24324 33232 24336
rect 22112 24296 28488 24324
rect 11195 24228 12434 24256
rect 15105 24259 15163 24265
rect 11195 24225 11207 24228
rect 11149 24219 11207 24225
rect 11532 24200 11560 24228
rect 15105 24225 15117 24259
rect 15151 24225 15163 24259
rect 15105 24219 15163 24225
rect 15381 24259 15439 24265
rect 15381 24225 15393 24259
rect 15427 24256 15439 24259
rect 15654 24256 15660 24268
rect 15427 24228 15660 24256
rect 15427 24225 15439 24228
rect 15381 24219 15439 24225
rect 15654 24216 15660 24228
rect 15712 24216 15718 24268
rect 17586 24216 17592 24268
rect 17644 24256 17650 24268
rect 17644 24228 18460 24256
rect 17644 24216 17650 24228
rect 10686 24191 10744 24197
rect 10686 24157 10698 24191
rect 10732 24188 10744 24191
rect 11422 24188 11428 24200
rect 10732 24160 11428 24188
rect 10732 24157 10744 24160
rect 10686 24151 10744 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11514 24148 11520 24200
rect 11572 24148 11578 24200
rect 11698 24148 11704 24200
rect 11756 24188 11762 24200
rect 11793 24191 11851 24197
rect 11793 24188 11805 24191
rect 11756 24160 11805 24188
rect 11756 24148 11762 24160
rect 11793 24157 11805 24160
rect 11839 24157 11851 24191
rect 12066 24188 12072 24200
rect 12027 24160 12072 24188
rect 11793 24151 11851 24157
rect 11808 24120 11836 24151
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 13357 24191 13415 24197
rect 13357 24157 13369 24191
rect 13403 24188 13415 24191
rect 13814 24188 13820 24200
rect 13403 24160 13820 24188
rect 13403 24157 13415 24160
rect 13357 24151 13415 24157
rect 13814 24148 13820 24160
rect 13872 24188 13878 24200
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 13872 24160 14105 24188
rect 13872 24148 13878 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 15013 24191 15071 24197
rect 15013 24157 15025 24191
rect 15059 24157 15071 24191
rect 15013 24151 15071 24157
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24188 16083 24191
rect 16666 24188 16672 24200
rect 16071 24160 16672 24188
rect 16071 24157 16083 24160
rect 16025 24151 16083 24157
rect 12529 24123 12587 24129
rect 12529 24120 12541 24123
rect 11808 24092 12541 24120
rect 12529 24089 12541 24092
rect 12575 24120 12587 24123
rect 13170 24120 13176 24132
rect 12575 24092 13176 24120
rect 12575 24089 12587 24092
rect 12529 24083 12587 24089
rect 13170 24080 13176 24092
rect 13228 24080 13234 24132
rect 13906 24080 13912 24132
rect 13964 24120 13970 24132
rect 15028 24120 15056 24151
rect 16666 24148 16672 24160
rect 16724 24148 16730 24200
rect 16942 24188 16948 24200
rect 16903 24160 16948 24188
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 18432 24188 18460 24228
rect 18690 24216 18696 24268
rect 18748 24256 18754 24268
rect 22112 24265 22140 24296
rect 20257 24259 20315 24265
rect 20257 24256 20269 24259
rect 18748 24228 20269 24256
rect 18748 24216 18754 24228
rect 20257 24225 20269 24228
rect 20303 24225 20315 24259
rect 20257 24219 20315 24225
rect 22097 24259 22155 24265
rect 22097 24225 22109 24259
rect 22143 24225 22155 24259
rect 26697 24259 26755 24265
rect 22097 24219 22155 24225
rect 25424 24228 26648 24256
rect 25424 24197 25452 24228
rect 26620 24200 26648 24228
rect 26697 24225 26709 24259
rect 26743 24256 26755 24259
rect 27982 24256 27988 24268
rect 26743 24228 27988 24256
rect 26743 24225 26755 24228
rect 26697 24219 26755 24225
rect 27982 24216 27988 24228
rect 28040 24216 28046 24268
rect 28350 24256 28356 24268
rect 28311 24228 28356 24256
rect 28350 24216 28356 24228
rect 28408 24216 28414 24268
rect 25700 24197 25820 24198
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 18432 24160 19257 24188
rect 19245 24157 19257 24160
rect 19291 24157 19303 24191
rect 23293 24191 23351 24197
rect 23293 24188 23305 24191
rect 19245 24151 19303 24157
rect 22112 24160 23305 24188
rect 22112 24132 22140 24160
rect 23293 24157 23305 24160
rect 23339 24157 23351 24191
rect 23293 24151 23351 24157
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24157 25467 24191
rect 25700 24191 25835 24197
rect 25700 24188 25789 24191
rect 25409 24151 25467 24157
rect 25516 24170 25789 24188
rect 25516 24160 25728 24170
rect 16850 24120 16856 24132
rect 13964 24092 16856 24120
rect 13964 24080 13970 24092
rect 16850 24080 16856 24092
rect 16908 24080 16914 24132
rect 17218 24120 17224 24132
rect 17179 24092 17224 24120
rect 17218 24080 17224 24092
rect 17276 24080 17282 24132
rect 19337 24123 19395 24129
rect 19337 24120 19349 24123
rect 18446 24092 19349 24120
rect 19337 24089 19349 24092
rect 19383 24089 19395 24123
rect 19337 24083 19395 24089
rect 20441 24123 20499 24129
rect 20441 24089 20453 24123
rect 20487 24120 20499 24123
rect 20622 24120 20628 24132
rect 20487 24092 20628 24120
rect 20487 24089 20499 24092
rect 20441 24083 20499 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 22094 24080 22100 24132
rect 22152 24080 22158 24132
rect 25130 24080 25136 24132
rect 25188 24120 25194 24132
rect 25516 24120 25544 24160
rect 25777 24157 25789 24170
rect 25823 24157 25835 24191
rect 25777 24151 25835 24157
rect 26418 24148 26424 24200
rect 26476 24148 26482 24200
rect 26602 24188 26608 24200
rect 26563 24160 26608 24188
rect 26602 24148 26608 24160
rect 26660 24148 26666 24200
rect 27614 24148 27620 24200
rect 27672 24188 27678 24200
rect 28074 24188 28080 24200
rect 27672 24160 28080 24188
rect 27672 24148 27678 24160
rect 28074 24148 28080 24160
rect 28132 24188 28138 24200
rect 28261 24191 28319 24197
rect 28261 24188 28273 24191
rect 28132 24160 28273 24188
rect 28132 24148 28138 24160
rect 28261 24157 28273 24160
rect 28307 24157 28319 24191
rect 28261 24151 28319 24157
rect 25188 24092 25544 24120
rect 25593 24123 25651 24129
rect 25188 24080 25194 24092
rect 25593 24089 25605 24123
rect 25639 24089 25651 24123
rect 25593 24083 25651 24089
rect 25685 24123 25743 24129
rect 25685 24089 25697 24123
rect 25731 24120 25743 24123
rect 26436 24120 26464 24148
rect 25731 24092 26464 24120
rect 28460 24120 28488 24296
rect 28966 24296 33232 24324
rect 28534 24197 28540 24200
rect 28530 24151 28540 24197
rect 28592 24188 28598 24200
rect 28966 24188 28994 24296
rect 33226 24284 33232 24296
rect 33284 24284 33290 24336
rect 34054 24284 34060 24336
rect 34112 24324 34118 24336
rect 34112 24296 40724 24324
rect 34112 24284 34118 24296
rect 31018 24216 31024 24268
rect 31076 24256 31082 24268
rect 31113 24259 31171 24265
rect 31113 24256 31125 24259
rect 31076 24228 31125 24256
rect 31076 24216 31082 24228
rect 31113 24225 31125 24228
rect 31159 24225 31171 24259
rect 33244 24256 33272 24284
rect 35618 24256 35624 24268
rect 33244 24228 35624 24256
rect 31113 24219 31171 24225
rect 35618 24216 35624 24228
rect 35676 24216 35682 24268
rect 40402 24256 40408 24268
rect 40363 24228 40408 24256
rect 40402 24216 40408 24228
rect 40460 24216 40466 24268
rect 40696 24265 40724 24296
rect 40681 24259 40739 24265
rect 40681 24225 40693 24259
rect 40727 24225 40739 24259
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 40681 24219 40739 24225
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48133 24259 48191 24265
rect 48133 24225 48145 24259
rect 48179 24256 48191 24259
rect 48222 24256 48228 24268
rect 48179 24228 48228 24256
rect 48179 24225 48191 24228
rect 48133 24219 48191 24225
rect 48222 24216 48228 24228
rect 48280 24216 48286 24268
rect 28592 24160 28994 24188
rect 30101 24191 30159 24197
rect 28534 24148 28540 24151
rect 28592 24148 28598 24160
rect 30101 24157 30113 24191
rect 30147 24157 30159 24191
rect 30101 24151 30159 24157
rect 30285 24191 30343 24197
rect 30285 24157 30297 24191
rect 30331 24188 30343 24191
rect 34698 24188 34704 24200
rect 30331 24160 30972 24188
rect 34659 24160 34704 24188
rect 30331 24157 30343 24160
rect 30285 24151 30343 24157
rect 30116 24120 30144 24151
rect 30558 24120 30564 24132
rect 28460 24092 28856 24120
rect 30116 24092 30564 24120
rect 25731 24089 25743 24092
rect 25685 24083 25743 24089
rect 10689 24055 10747 24061
rect 10689 24021 10701 24055
rect 10735 24052 10747 24055
rect 11146 24052 11152 24064
rect 10735 24024 11152 24052
rect 10735 24021 10747 24024
rect 10689 24015 10747 24021
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 11609 24055 11667 24061
rect 11609 24021 11621 24055
rect 11655 24052 11667 24055
rect 11790 24052 11796 24064
rect 11655 24024 11796 24052
rect 11655 24021 11667 24024
rect 11609 24015 11667 24021
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 11974 24052 11980 24064
rect 11935 24024 11980 24052
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 12710 24012 12716 24064
rect 12768 24061 12774 24064
rect 12768 24055 12787 24061
rect 12775 24021 12787 24055
rect 12768 24015 12787 24021
rect 13449 24055 13507 24061
rect 13449 24021 13461 24055
rect 13495 24052 13507 24055
rect 14090 24052 14096 24064
rect 13495 24024 14096 24052
rect 13495 24021 13507 24024
rect 13449 24015 13507 24021
rect 12768 24012 12774 24015
rect 14090 24012 14096 24024
rect 14148 24012 14154 24064
rect 15378 24012 15384 24064
rect 15436 24052 15442 24064
rect 16025 24055 16083 24061
rect 16025 24052 16037 24055
rect 15436 24024 16037 24052
rect 15436 24012 15442 24024
rect 16025 24021 16037 24024
rect 16071 24021 16083 24055
rect 16025 24015 16083 24021
rect 18506 24012 18512 24064
rect 18564 24052 18570 24064
rect 18693 24055 18751 24061
rect 18693 24052 18705 24055
rect 18564 24024 18705 24052
rect 18564 24012 18570 24024
rect 18693 24021 18705 24024
rect 18739 24021 18751 24055
rect 25608 24052 25636 24083
rect 25774 24052 25780 24064
rect 25608 24024 25780 24052
rect 18693 24015 18751 24021
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 25961 24055 26019 24061
rect 25961 24021 25973 24055
rect 26007 24052 26019 24055
rect 26142 24052 26148 24064
rect 26007 24024 26148 24052
rect 26007 24021 26019 24024
rect 25961 24015 26019 24021
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 26418 24012 26424 24064
rect 26476 24052 26482 24064
rect 26973 24055 27031 24061
rect 26973 24052 26985 24055
rect 26476 24024 26985 24052
rect 26476 24012 26482 24024
rect 26973 24021 26985 24024
rect 27019 24021 27031 24055
rect 26973 24015 27031 24021
rect 28442 24012 28448 24064
rect 28500 24052 28506 24064
rect 28718 24052 28724 24064
rect 28500 24024 28724 24052
rect 28500 24012 28506 24024
rect 28718 24012 28724 24024
rect 28776 24012 28782 24064
rect 28828 24052 28856 24092
rect 30558 24080 30564 24092
rect 30616 24120 30622 24132
rect 30944 24129 30972 24160
rect 34698 24148 34704 24160
rect 34756 24148 34762 24200
rect 40218 24188 40224 24200
rect 40179 24160 40224 24188
rect 40218 24148 40224 24160
rect 40276 24148 40282 24200
rect 43346 24188 43352 24200
rect 43307 24160 43352 24188
rect 43346 24148 43352 24160
rect 43404 24148 43410 24200
rect 43530 24188 43536 24200
rect 43491 24160 43536 24188
rect 43530 24148 43536 24160
rect 43588 24148 43594 24200
rect 43993 24191 44051 24197
rect 43993 24157 44005 24191
rect 44039 24188 44051 24191
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44039 24160 45201 24188
rect 44039 24157 44051 24160
rect 43993 24151 44051 24157
rect 45189 24157 45201 24160
rect 45235 24188 45247 24191
rect 45462 24188 45468 24200
rect 45235 24160 45468 24188
rect 45235 24157 45247 24160
rect 45189 24151 45247 24157
rect 45462 24148 45468 24160
rect 45520 24148 45526 24200
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 46293 24191 46351 24197
rect 46293 24188 46305 24191
rect 45612 24160 46305 24188
rect 45612 24148 45618 24160
rect 46293 24157 46305 24160
rect 46339 24157 46351 24191
rect 46293 24151 46351 24157
rect 30745 24123 30803 24129
rect 30745 24120 30757 24123
rect 30616 24092 30757 24120
rect 30616 24080 30622 24092
rect 30745 24089 30757 24092
rect 30791 24089 30803 24123
rect 30745 24083 30803 24089
rect 30929 24123 30987 24129
rect 30929 24089 30941 24123
rect 30975 24120 30987 24123
rect 31754 24120 31760 24132
rect 30975 24092 31760 24120
rect 30975 24089 30987 24092
rect 30929 24083 30987 24089
rect 31754 24080 31760 24092
rect 31812 24120 31818 24132
rect 32950 24120 32956 24132
rect 31812 24092 32956 24120
rect 31812 24080 31818 24092
rect 32950 24080 32956 24092
rect 33008 24080 33014 24132
rect 44266 24120 44272 24132
rect 44179 24092 44272 24120
rect 44266 24080 44272 24092
rect 44324 24120 44330 24132
rect 45094 24120 45100 24132
rect 44324 24092 45100 24120
rect 44324 24080 44330 24092
rect 45094 24080 45100 24092
rect 45152 24080 45158 24132
rect 45741 24123 45799 24129
rect 45741 24089 45753 24123
rect 45787 24120 45799 24123
rect 46014 24120 46020 24132
rect 45787 24092 46020 24120
rect 45787 24089 45799 24092
rect 45741 24083 45799 24089
rect 46014 24080 46020 24092
rect 46072 24120 46078 24132
rect 46474 24120 46480 24132
rect 46072 24092 46480 24120
rect 46072 24080 46078 24092
rect 46474 24080 46480 24092
rect 46532 24080 46538 24132
rect 37274 24052 37280 24064
rect 28828 24024 37280 24052
rect 37274 24012 37280 24024
rect 37332 24012 37338 24064
rect 43533 24055 43591 24061
rect 43533 24021 43545 24055
rect 43579 24052 43591 24055
rect 43806 24052 43812 24064
rect 43579 24024 43812 24052
rect 43579 24021 43591 24024
rect 43533 24015 43591 24021
rect 43806 24012 43812 24024
rect 43864 24012 43870 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 8938 23848 8944 23860
rect 8899 23820 8944 23848
rect 8938 23808 8944 23820
rect 8996 23808 9002 23860
rect 11146 23808 11152 23860
rect 11204 23848 11210 23860
rect 12066 23848 12072 23860
rect 11204 23820 12072 23848
rect 11204 23808 11210 23820
rect 12066 23808 12072 23820
rect 12124 23808 12130 23860
rect 17218 23808 17224 23860
rect 17276 23848 17282 23860
rect 17865 23851 17923 23857
rect 17865 23848 17877 23851
rect 17276 23820 17877 23848
rect 17276 23808 17282 23820
rect 17865 23817 17877 23820
rect 17911 23817 17923 23851
rect 17865 23811 17923 23817
rect 18627 23851 18685 23857
rect 18627 23817 18639 23851
rect 18673 23848 18685 23851
rect 19334 23848 19340 23860
rect 18673 23820 19340 23848
rect 18673 23817 18685 23820
rect 18627 23811 18685 23817
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 19978 23848 19984 23860
rect 19939 23820 19984 23848
rect 19978 23808 19984 23820
rect 20036 23808 20042 23860
rect 20622 23848 20628 23860
rect 20583 23820 20628 23848
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 26329 23851 26387 23857
rect 26329 23817 26341 23851
rect 26375 23848 26387 23851
rect 27798 23848 27804 23860
rect 26375 23820 27804 23848
rect 26375 23817 26387 23820
rect 26329 23811 26387 23817
rect 27798 23808 27804 23820
rect 27856 23808 27862 23860
rect 27982 23808 27988 23860
rect 28040 23848 28046 23860
rect 28442 23848 28448 23860
rect 28040 23820 28448 23848
rect 28040 23808 28046 23820
rect 28442 23808 28448 23820
rect 28500 23808 28506 23860
rect 30190 23848 30196 23860
rect 29564 23820 30196 23848
rect 11514 23780 11520 23792
rect 11475 23752 11520 23780
rect 11514 23740 11520 23752
rect 11572 23740 11578 23792
rect 14090 23780 14096 23792
rect 14051 23752 14096 23780
rect 14090 23740 14096 23752
rect 14148 23740 14154 23792
rect 18414 23780 18420 23792
rect 18375 23752 18420 23780
rect 18414 23740 18420 23752
rect 18472 23740 18478 23792
rect 28074 23780 28080 23792
rect 28035 23752 28080 23780
rect 28074 23740 28080 23752
rect 28132 23740 28138 23792
rect 1394 23712 1400 23724
rect 1355 23684 1400 23712
rect 1394 23672 1400 23684
rect 1452 23672 1458 23724
rect 8849 23715 8907 23721
rect 8849 23681 8861 23715
rect 8895 23712 8907 23715
rect 8938 23712 8944 23724
rect 8895 23684 8944 23712
rect 8895 23681 8907 23684
rect 8849 23675 8907 23681
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23712 11023 23715
rect 13906 23712 13912 23724
rect 11011 23684 12020 23712
rect 13867 23684 13912 23712
rect 11011 23681 11023 23684
rect 10965 23675 11023 23681
rect 11992 23653 12020 23684
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23712 16727 23715
rect 17402 23712 17408 23724
rect 16715 23684 17408 23712
rect 16715 23681 16727 23684
rect 16669 23675 16727 23681
rect 17402 23672 17408 23684
rect 17460 23672 17466 23724
rect 17770 23712 17776 23724
rect 17731 23684 17776 23712
rect 17770 23672 17776 23684
rect 17828 23672 17834 23724
rect 17957 23715 18015 23721
rect 17957 23681 17969 23715
rect 18003 23712 18015 23715
rect 18782 23712 18788 23724
rect 18003 23684 18788 23712
rect 18003 23681 18015 23684
rect 17957 23675 18015 23681
rect 18782 23672 18788 23684
rect 18840 23672 18846 23724
rect 19889 23715 19947 23721
rect 19889 23681 19901 23715
rect 19935 23712 19947 23715
rect 20533 23715 20591 23721
rect 20533 23712 20545 23715
rect 19935 23684 20545 23712
rect 19935 23681 19947 23684
rect 19889 23675 19947 23681
rect 20533 23681 20545 23684
rect 20579 23712 20591 23715
rect 20714 23712 20720 23724
rect 20579 23684 20720 23712
rect 20579 23681 20591 23684
rect 20533 23675 20591 23681
rect 20714 23672 20720 23684
rect 20772 23672 20778 23724
rect 21821 23715 21879 23721
rect 21821 23681 21833 23715
rect 21867 23712 21879 23715
rect 22094 23712 22100 23724
rect 21867 23684 22100 23712
rect 21867 23681 21879 23684
rect 21821 23675 21879 23681
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 26142 23712 26148 23724
rect 26103 23684 26148 23712
rect 26142 23672 26148 23684
rect 26200 23672 26206 23724
rect 26418 23672 26424 23724
rect 26476 23712 26482 23724
rect 28261 23715 28319 23721
rect 26476 23684 26521 23712
rect 26476 23672 26482 23684
rect 28261 23681 28273 23715
rect 28307 23712 28319 23715
rect 28350 23712 28356 23724
rect 28307 23684 28356 23712
rect 28307 23681 28319 23684
rect 28261 23675 28319 23681
rect 28350 23672 28356 23684
rect 28408 23672 28414 23724
rect 28718 23672 28724 23724
rect 28776 23712 28782 23724
rect 29564 23721 29592 23820
rect 30190 23808 30196 23820
rect 30248 23808 30254 23860
rect 30558 23848 30564 23860
rect 30519 23820 30564 23848
rect 30558 23808 30564 23820
rect 30616 23848 30622 23860
rect 31205 23851 31263 23857
rect 31205 23848 31217 23851
rect 30616 23820 31217 23848
rect 30616 23808 30622 23820
rect 31205 23817 31217 23820
rect 31251 23817 31263 23851
rect 31205 23811 31263 23817
rect 34057 23851 34115 23857
rect 34057 23817 34069 23851
rect 34103 23848 34115 23851
rect 34698 23848 34704 23860
rect 34103 23820 34704 23848
rect 34103 23817 34115 23820
rect 34057 23811 34115 23817
rect 29641 23783 29699 23789
rect 29641 23749 29653 23783
rect 29687 23780 29699 23783
rect 30377 23783 30435 23789
rect 29687 23752 30052 23780
rect 29687 23749 29699 23752
rect 29641 23743 29699 23749
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 28776 23684 29561 23712
rect 28776 23672 28782 23684
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29730 23712 29736 23724
rect 29691 23684 29736 23712
rect 29549 23675 29607 23681
rect 29730 23672 29736 23684
rect 29788 23672 29794 23724
rect 11977 23647 12035 23653
rect 11624 23616 11928 23644
rect 1581 23579 1639 23585
rect 1581 23545 1593 23579
rect 1627 23576 1639 23579
rect 11624 23576 11652 23616
rect 11790 23576 11796 23588
rect 1627 23548 11652 23576
rect 11751 23548 11796 23576
rect 1627 23545 1639 23548
rect 1581 23539 1639 23545
rect 11790 23536 11796 23548
rect 11848 23536 11854 23588
rect 11900 23576 11928 23616
rect 11977 23613 11989 23647
rect 12023 23613 12035 23647
rect 11977 23607 12035 23613
rect 14182 23604 14188 23656
rect 14240 23644 14246 23656
rect 14369 23647 14427 23653
rect 14369 23644 14381 23647
rect 14240 23616 14381 23644
rect 14240 23604 14246 23616
rect 14369 23613 14381 23616
rect 14415 23613 14427 23647
rect 30024 23644 30052 23752
rect 30377 23749 30389 23783
rect 30423 23780 30435 23783
rect 30466 23780 30472 23792
rect 30423 23752 30472 23780
rect 30423 23749 30435 23752
rect 30377 23743 30435 23749
rect 30466 23740 30472 23752
rect 30524 23740 30530 23792
rect 32766 23780 32772 23792
rect 32679 23752 32772 23780
rect 30190 23672 30196 23724
rect 30248 23712 30254 23724
rect 30248 23684 30293 23712
rect 30248 23672 30254 23684
rect 30926 23672 30932 23724
rect 30984 23712 30990 23724
rect 32692 23721 32720 23752
rect 32766 23740 32772 23752
rect 32824 23780 32830 23792
rect 33410 23780 33416 23792
rect 32824 23752 33416 23780
rect 32824 23740 32830 23752
rect 33410 23740 33416 23752
rect 33468 23780 33474 23792
rect 34072 23780 34100 23811
rect 34698 23808 34704 23820
rect 34756 23808 34762 23860
rect 40218 23808 40224 23860
rect 40276 23848 40282 23860
rect 41509 23851 41567 23857
rect 41509 23848 41521 23851
rect 40276 23820 41521 23848
rect 40276 23808 40282 23820
rect 41509 23817 41521 23820
rect 41555 23817 41567 23851
rect 41509 23811 41567 23817
rect 43165 23851 43223 23857
rect 43165 23817 43177 23851
rect 43211 23848 43223 23851
rect 43346 23848 43352 23860
rect 43211 23820 43352 23848
rect 43211 23817 43223 23820
rect 43165 23811 43223 23817
rect 43346 23808 43352 23820
rect 43404 23808 43410 23860
rect 44177 23851 44235 23857
rect 44177 23817 44189 23851
rect 44223 23848 44235 23851
rect 45554 23848 45560 23860
rect 44223 23820 45560 23848
rect 44223 23817 44235 23820
rect 44177 23811 44235 23817
rect 45554 23808 45560 23820
rect 45612 23808 45618 23860
rect 42794 23780 42800 23792
rect 33468 23752 34100 23780
rect 42755 23752 42800 23780
rect 33468 23740 33474 23752
rect 42794 23740 42800 23752
rect 42852 23740 42858 23792
rect 42981 23783 43039 23789
rect 42981 23749 42993 23783
rect 43027 23780 43039 23783
rect 44358 23780 44364 23792
rect 43027 23752 44364 23780
rect 43027 23749 43039 23752
rect 42981 23743 43039 23749
rect 44358 23740 44364 23752
rect 44416 23740 44422 23792
rect 45002 23740 45008 23792
rect 45060 23780 45066 23792
rect 45189 23783 45247 23789
rect 45189 23780 45201 23783
rect 45060 23752 45201 23780
rect 45060 23740 45066 23752
rect 45189 23749 45201 23752
rect 45235 23780 45247 23783
rect 45370 23780 45376 23792
rect 45235 23752 45376 23780
rect 45235 23749 45247 23752
rect 45189 23743 45247 23749
rect 45370 23740 45376 23752
rect 45428 23740 45434 23792
rect 31021 23715 31079 23721
rect 31021 23712 31033 23715
rect 30984 23684 31033 23712
rect 30984 23672 30990 23684
rect 31021 23681 31033 23684
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 31297 23715 31355 23721
rect 31297 23681 31309 23715
rect 31343 23681 31355 23715
rect 31297 23675 31355 23681
rect 32677 23715 32735 23721
rect 32677 23681 32689 23715
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 33873 23715 33931 23721
rect 33873 23681 33885 23715
rect 33919 23712 33931 23715
rect 34422 23712 34428 23724
rect 33919 23684 34428 23712
rect 33919 23681 33931 23684
rect 33873 23675 33931 23681
rect 31312 23644 31340 23675
rect 34422 23672 34428 23684
rect 34480 23672 34486 23724
rect 38378 23672 38384 23724
rect 38436 23712 38442 23724
rect 40129 23715 40187 23721
rect 40129 23712 40141 23715
rect 38436 23684 40141 23712
rect 38436 23672 38442 23684
rect 40129 23681 40141 23684
rect 40175 23681 40187 23715
rect 40129 23675 40187 23681
rect 41141 23715 41199 23721
rect 41141 23681 41153 23715
rect 41187 23712 41199 23715
rect 42610 23712 42616 23724
rect 41187 23684 42616 23712
rect 41187 23681 41199 23684
rect 41141 23675 41199 23681
rect 42610 23672 42616 23684
rect 42668 23672 42674 23724
rect 43806 23712 43812 23724
rect 43767 23684 43812 23712
rect 43806 23672 43812 23684
rect 43864 23672 43870 23724
rect 44913 23715 44971 23721
rect 44913 23681 44925 23715
rect 44959 23712 44971 23715
rect 45462 23712 45468 23724
rect 44959 23684 45468 23712
rect 44959 23681 44971 23684
rect 44913 23675 44971 23681
rect 45462 23672 45468 23684
rect 45520 23712 45526 23724
rect 45925 23715 45983 23721
rect 45925 23712 45937 23715
rect 45520 23684 45937 23712
rect 45520 23672 45526 23684
rect 45925 23681 45937 23684
rect 45971 23681 45983 23715
rect 47581 23715 47639 23721
rect 47581 23712 47593 23715
rect 45925 23675 45983 23681
rect 46308 23684 47593 23712
rect 46308 23656 46336 23684
rect 47581 23681 47593 23684
rect 47627 23681 47639 23715
rect 47581 23675 47639 23681
rect 30024 23616 31340 23644
rect 40221 23647 40279 23653
rect 14369 23607 14427 23613
rect 40221 23613 40233 23647
rect 40267 23613 40279 23647
rect 41049 23647 41107 23653
rect 41049 23644 41061 23647
rect 40221 23607 40279 23613
rect 40512 23616 41061 23644
rect 33594 23576 33600 23588
rect 11900 23548 33600 23576
rect 33594 23536 33600 23548
rect 33652 23536 33658 23588
rect 10781 23511 10839 23517
rect 10781 23477 10793 23511
rect 10827 23508 10839 23511
rect 11698 23508 11704 23520
rect 10827 23480 11704 23508
rect 10827 23477 10839 23480
rect 10781 23471 10839 23477
rect 11698 23468 11704 23480
rect 11756 23468 11762 23520
rect 16758 23508 16764 23520
rect 16719 23480 16764 23508
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 18322 23508 18328 23520
rect 16908 23480 18328 23508
rect 16908 23468 16914 23480
rect 18322 23468 18328 23480
rect 18380 23508 18386 23520
rect 18601 23511 18659 23517
rect 18601 23508 18613 23511
rect 18380 23480 18613 23508
rect 18380 23468 18386 23480
rect 18601 23477 18613 23480
rect 18647 23477 18659 23511
rect 18782 23508 18788 23520
rect 18743 23480 18788 23508
rect 18601 23471 18659 23477
rect 18782 23468 18788 23480
rect 18840 23468 18846 23520
rect 21910 23508 21916 23520
rect 21871 23480 21916 23508
rect 21910 23468 21916 23480
rect 21968 23468 21974 23520
rect 25314 23468 25320 23520
rect 25372 23508 25378 23520
rect 25961 23511 26019 23517
rect 25961 23508 25973 23511
rect 25372 23480 25973 23508
rect 25372 23468 25378 23480
rect 25961 23477 25973 23480
rect 26007 23477 26019 23511
rect 25961 23471 26019 23477
rect 26970 23468 26976 23520
rect 27028 23508 27034 23520
rect 28074 23508 28080 23520
rect 27028 23480 28080 23508
rect 27028 23468 27034 23480
rect 28074 23468 28080 23480
rect 28132 23508 28138 23520
rect 30926 23508 30932 23520
rect 28132 23480 30932 23508
rect 28132 23468 28138 23480
rect 30926 23468 30932 23480
rect 30984 23468 30990 23520
rect 31021 23511 31079 23517
rect 31021 23477 31033 23511
rect 31067 23508 31079 23511
rect 31202 23508 31208 23520
rect 31067 23480 31208 23508
rect 31067 23477 31079 23480
rect 31021 23471 31079 23477
rect 31202 23468 31208 23480
rect 31260 23468 31266 23520
rect 32766 23508 32772 23520
rect 32727 23480 32772 23508
rect 32766 23468 32772 23480
rect 32824 23468 32830 23520
rect 40236 23508 40264 23607
rect 40512 23585 40540 23616
rect 41049 23613 41061 23616
rect 41095 23613 41107 23647
rect 43714 23644 43720 23656
rect 43675 23616 43720 23644
rect 41049 23607 41107 23613
rect 43714 23604 43720 23616
rect 43772 23604 43778 23656
rect 46290 23644 46296 23656
rect 46251 23616 46296 23644
rect 46290 23604 46296 23616
rect 46348 23604 46354 23656
rect 40497 23579 40555 23585
rect 40497 23545 40509 23579
rect 40543 23545 40555 23579
rect 48038 23576 48044 23588
rect 40497 23539 40555 23545
rect 41386 23548 48044 23576
rect 41386 23508 41414 23548
rect 48038 23536 48044 23548
rect 48096 23536 48102 23588
rect 47670 23508 47676 23520
rect 40236 23480 41414 23508
rect 47631 23480 47676 23508
rect 47670 23468 47676 23480
rect 47728 23468 47734 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 16942 23264 16948 23316
rect 17000 23304 17006 23316
rect 17773 23307 17831 23313
rect 17773 23304 17785 23307
rect 17000 23276 17785 23304
rect 17000 23264 17006 23276
rect 17773 23273 17785 23276
rect 17819 23273 17831 23307
rect 17773 23267 17831 23273
rect 26602 23264 26608 23316
rect 26660 23304 26666 23316
rect 26789 23307 26847 23313
rect 26789 23304 26801 23307
rect 26660 23276 26801 23304
rect 26660 23264 26666 23276
rect 26789 23273 26801 23276
rect 26835 23273 26847 23307
rect 32950 23304 32956 23316
rect 32911 23276 32956 23304
rect 26789 23267 26847 23273
rect 32950 23264 32956 23276
rect 33008 23264 33014 23316
rect 42610 23264 42616 23316
rect 42668 23304 42674 23316
rect 43717 23307 43775 23313
rect 43717 23304 43729 23307
rect 42668 23276 43729 23304
rect 42668 23264 42674 23276
rect 43717 23273 43729 23276
rect 43763 23273 43775 23307
rect 43717 23267 43775 23273
rect 16850 23196 16856 23248
rect 16908 23236 16914 23248
rect 17129 23239 17187 23245
rect 17129 23236 17141 23239
rect 16908 23208 17141 23236
rect 16908 23196 16914 23208
rect 17129 23205 17141 23208
rect 17175 23205 17187 23239
rect 17129 23199 17187 23205
rect 28261 23239 28319 23245
rect 28261 23205 28273 23239
rect 28307 23236 28319 23239
rect 28810 23236 28816 23248
rect 28307 23208 28816 23236
rect 28307 23205 28319 23208
rect 28261 23199 28319 23205
rect 28810 23196 28816 23208
rect 28868 23196 28874 23248
rect 42794 23196 42800 23248
rect 42852 23236 42858 23248
rect 46658 23236 46664 23248
rect 42852 23208 44220 23236
rect 42852 23196 42858 23208
rect 11698 23168 11704 23180
rect 11659 23140 11704 23168
rect 11698 23128 11704 23140
rect 11756 23128 11762 23180
rect 15378 23168 15384 23180
rect 15339 23140 15384 23168
rect 15378 23128 15384 23140
rect 15436 23128 15442 23180
rect 15654 23168 15660 23180
rect 15615 23140 15660 23168
rect 15654 23128 15660 23140
rect 15712 23128 15718 23180
rect 16666 23128 16672 23180
rect 16724 23168 16730 23180
rect 20349 23171 20407 23177
rect 16724 23140 17724 23168
rect 16724 23128 16730 23140
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23069 10839 23103
rect 11422 23100 11428 23112
rect 11383 23072 11428 23100
rect 10781 23063 10839 23069
rect 10796 23032 10824 23063
rect 11422 23060 11428 23072
rect 11480 23060 11486 23112
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14642 23100 14648 23112
rect 14323 23072 14648 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14642 23060 14648 23072
rect 14700 23100 14706 23112
rect 15010 23100 15016 23112
rect 14700 23072 15016 23100
rect 14700 23060 14706 23072
rect 15010 23060 15016 23072
rect 15068 23060 15074 23112
rect 16758 23060 16764 23112
rect 16816 23060 16822 23112
rect 17696 23109 17724 23140
rect 20349 23137 20361 23171
rect 20395 23168 20407 23171
rect 20898 23168 20904 23180
rect 20395 23140 20904 23168
rect 20395 23137 20407 23140
rect 20349 23131 20407 23137
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 22738 23128 22744 23180
rect 22796 23168 22802 23180
rect 24946 23168 24952 23180
rect 22796 23140 24952 23168
rect 22796 23128 22802 23140
rect 24946 23128 24952 23140
rect 25004 23168 25010 23180
rect 25041 23171 25099 23177
rect 25041 23168 25053 23171
rect 25004 23140 25053 23168
rect 25004 23128 25010 23140
rect 25041 23137 25053 23140
rect 25087 23168 25099 23171
rect 25406 23168 25412 23180
rect 25087 23140 25412 23168
rect 25087 23137 25099 23140
rect 25041 23131 25099 23137
rect 25406 23128 25412 23140
rect 25464 23128 25470 23180
rect 27709 23171 27767 23177
rect 27709 23137 27721 23171
rect 27755 23168 27767 23171
rect 27755 23140 28580 23168
rect 27755 23137 27767 23140
rect 27709 23131 27767 23137
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23069 17739 23103
rect 19242 23100 19248 23112
rect 19203 23072 19248 23100
rect 17681 23063 17739 23069
rect 19242 23060 19248 23072
rect 19300 23060 19306 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23069 20131 23103
rect 20073 23063 20131 23069
rect 11330 23032 11336 23044
rect 10796 23004 11336 23032
rect 11330 22992 11336 23004
rect 11388 22992 11394 23044
rect 12434 22992 12440 23044
rect 12492 22992 12498 23044
rect 20088 23032 20116 23063
rect 23198 23060 23204 23112
rect 23256 23100 23262 23112
rect 23385 23103 23443 23109
rect 23385 23100 23397 23103
rect 23256 23072 23397 23100
rect 23256 23060 23262 23072
rect 23385 23069 23397 23072
rect 23431 23069 23443 23103
rect 27614 23100 27620 23112
rect 27575 23072 27620 23100
rect 23385 23063 23443 23069
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 27801 23103 27859 23109
rect 27801 23069 27813 23103
rect 27847 23100 27859 23103
rect 28350 23100 28356 23112
rect 27847 23072 28356 23100
rect 27847 23069 27859 23072
rect 27801 23063 27859 23069
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 28552 23109 28580 23140
rect 30374 23128 30380 23180
rect 30432 23128 30438 23180
rect 31205 23171 31263 23177
rect 31205 23137 31217 23171
rect 31251 23168 31263 23171
rect 32030 23168 32036 23180
rect 31251 23140 32036 23168
rect 31251 23137 31263 23140
rect 31205 23131 31263 23137
rect 32030 23128 32036 23140
rect 32088 23128 32094 23180
rect 40218 23128 40224 23180
rect 40276 23168 40282 23180
rect 40773 23171 40831 23177
rect 40773 23168 40785 23171
rect 40276 23140 40785 23168
rect 40276 23128 40282 23140
rect 40773 23137 40785 23140
rect 40819 23137 40831 23171
rect 41414 23168 41420 23180
rect 41375 23140 41420 23168
rect 40773 23131 40831 23137
rect 41414 23128 41420 23140
rect 41472 23128 41478 23180
rect 43346 23128 43352 23180
rect 43404 23168 43410 23180
rect 43441 23171 43499 23177
rect 43441 23168 43453 23171
rect 43404 23140 43453 23168
rect 43404 23128 43410 23140
rect 43441 23137 43453 23140
rect 43487 23137 43499 23171
rect 43441 23131 43499 23137
rect 28537 23103 28595 23109
rect 28537 23069 28549 23103
rect 28583 23069 28595 23103
rect 28537 23063 28595 23069
rect 29730 23060 29736 23112
rect 29788 23100 29794 23112
rect 30190 23100 30196 23112
rect 29788 23072 30196 23100
rect 29788 23060 29794 23072
rect 30190 23060 30196 23072
rect 30248 23060 30254 23112
rect 30392 23100 30420 23128
rect 30469 23103 30527 23109
rect 30469 23100 30481 23103
rect 30392 23072 30481 23100
rect 30469 23069 30481 23072
rect 30515 23069 30527 23103
rect 30469 23063 30527 23069
rect 30561 23103 30619 23109
rect 30561 23069 30573 23103
rect 30607 23100 30619 23103
rect 30742 23100 30748 23112
rect 30607 23072 30748 23100
rect 30607 23069 30619 23072
rect 30561 23063 30619 23069
rect 30742 23060 30748 23072
rect 30800 23060 30806 23112
rect 33410 23100 33416 23112
rect 33371 23072 33416 23100
rect 33410 23060 33416 23072
rect 33468 23060 33474 23112
rect 40313 23103 40371 23109
rect 40313 23069 40325 23103
rect 40359 23100 40371 23103
rect 40678 23100 40684 23112
rect 40359 23072 40684 23100
rect 40359 23069 40371 23072
rect 40313 23063 40371 23069
rect 40678 23060 40684 23072
rect 40736 23060 40742 23112
rect 43070 23060 43076 23112
rect 43128 23100 43134 23112
rect 43533 23103 43591 23109
rect 43533 23100 43545 23103
rect 43128 23072 43545 23100
rect 43128 23060 43134 23072
rect 43533 23069 43545 23072
rect 43579 23100 43591 23103
rect 43714 23100 43720 23112
rect 43579 23072 43720 23100
rect 43579 23069 43591 23072
rect 43533 23063 43591 23069
rect 43714 23060 43720 23072
rect 43772 23060 43778 23112
rect 44192 23109 44220 23208
rect 46308 23208 46664 23236
rect 46308 23177 46336 23208
rect 46658 23196 46664 23208
rect 46716 23196 46722 23248
rect 46293 23171 46351 23177
rect 46293 23137 46305 23171
rect 46339 23137 46351 23171
rect 46293 23131 46351 23137
rect 46477 23171 46535 23177
rect 46477 23137 46489 23171
rect 46523 23168 46535 23171
rect 47670 23168 47676 23180
rect 46523 23140 47676 23168
rect 46523 23137 46535 23140
rect 46477 23131 46535 23137
rect 47670 23128 47676 23140
rect 47728 23128 47734 23180
rect 48130 23168 48136 23180
rect 48091 23140 48136 23168
rect 48130 23128 48136 23140
rect 48188 23128 48194 23180
rect 44177 23103 44235 23109
rect 44177 23069 44189 23103
rect 44223 23069 44235 23103
rect 44358 23100 44364 23112
rect 44319 23072 44364 23100
rect 44177 23063 44235 23069
rect 44358 23060 44364 23072
rect 44416 23060 44422 23112
rect 45373 23103 45431 23109
rect 45373 23069 45385 23103
rect 45419 23100 45431 23103
rect 45462 23100 45468 23112
rect 45419 23072 45468 23100
rect 45419 23069 45431 23072
rect 45373 23063 45431 23069
rect 45462 23060 45468 23072
rect 45520 23060 45526 23112
rect 21910 23032 21916 23044
rect 20088 23004 20300 23032
rect 21574 23004 21916 23032
rect 10226 22924 10232 22976
rect 10284 22964 10290 22976
rect 10781 22967 10839 22973
rect 10781 22964 10793 22967
rect 10284 22936 10793 22964
rect 10284 22924 10290 22936
rect 10781 22933 10793 22936
rect 10827 22933 10839 22967
rect 13170 22964 13176 22976
rect 13131 22936 13176 22964
rect 10781 22927 10839 22933
rect 13170 22924 13176 22936
rect 13228 22924 13234 22976
rect 13906 22924 13912 22976
rect 13964 22964 13970 22976
rect 14461 22967 14519 22973
rect 14461 22964 14473 22967
rect 13964 22936 14473 22964
rect 13964 22924 13970 22936
rect 14461 22933 14473 22936
rect 14507 22933 14519 22967
rect 14461 22927 14519 22933
rect 19613 22967 19671 22973
rect 19613 22933 19625 22967
rect 19659 22964 19671 22967
rect 20162 22964 20168 22976
rect 19659 22936 20168 22964
rect 19659 22933 19671 22936
rect 19613 22927 19671 22933
rect 20162 22924 20168 22936
rect 20220 22924 20226 22976
rect 20272 22964 20300 23004
rect 21910 22992 21916 23004
rect 21968 22992 21974 23044
rect 25314 23032 25320 23044
rect 25275 23004 25320 23032
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 27706 23032 27712 23044
rect 26542 23004 27712 23032
rect 27706 22992 27712 23004
rect 27764 22992 27770 23044
rect 28074 22992 28080 23044
rect 28132 23032 28138 23044
rect 28261 23035 28319 23041
rect 28261 23032 28273 23035
rect 28132 23004 28273 23032
rect 28132 22992 28138 23004
rect 28261 23001 28273 23004
rect 28307 23001 28319 23035
rect 28368 23032 28396 23060
rect 28718 23032 28724 23044
rect 28368 23004 28724 23032
rect 28261 22995 28319 23001
rect 28718 22992 28724 23004
rect 28776 22992 28782 23044
rect 30282 22992 30288 23044
rect 30340 23032 30346 23044
rect 30377 23035 30435 23041
rect 30377 23032 30389 23035
rect 30340 23004 30389 23032
rect 30340 22992 30346 23004
rect 30377 23001 30389 23004
rect 30423 23001 30435 23035
rect 30377 22995 30435 23001
rect 30650 22992 30656 23044
rect 30708 23032 30714 23044
rect 31481 23035 31539 23041
rect 31481 23032 31493 23035
rect 30708 23004 31493 23032
rect 30708 22992 30714 23004
rect 31481 23001 31493 23004
rect 31527 23001 31539 23035
rect 32766 23032 32772 23044
rect 32706 23004 32772 23032
rect 31481 22995 31539 23001
rect 32766 22992 32772 23004
rect 32824 22992 32830 23044
rect 40957 23035 41015 23041
rect 40957 23001 40969 23035
rect 41003 23001 41015 23035
rect 40957 22995 41015 23001
rect 45649 23035 45707 23041
rect 45649 23001 45661 23035
rect 45695 23032 45707 23035
rect 45830 23032 45836 23044
rect 45695 23004 45836 23032
rect 45695 23001 45707 23004
rect 45649 22995 45707 23001
rect 20622 22964 20628 22976
rect 20272 22936 20628 22964
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 21818 22964 21824 22976
rect 21779 22936 21824 22964
rect 21818 22924 21824 22936
rect 21876 22924 21882 22976
rect 23474 22964 23480 22976
rect 23435 22936 23480 22964
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 28442 22964 28448 22976
rect 28403 22936 28448 22964
rect 28442 22924 28448 22936
rect 28500 22924 28506 22976
rect 30745 22967 30803 22973
rect 30745 22933 30757 22967
rect 30791 22964 30803 22967
rect 31018 22964 31024 22976
rect 30791 22936 31024 22964
rect 30791 22933 30803 22936
rect 30745 22927 30803 22933
rect 31018 22924 31024 22936
rect 31076 22924 31082 22976
rect 33502 22964 33508 22976
rect 33463 22936 33508 22964
rect 33502 22924 33508 22936
rect 33560 22924 33566 22976
rect 40129 22967 40187 22973
rect 40129 22933 40141 22967
rect 40175 22964 40187 22967
rect 40972 22964 41000 22995
rect 45830 22992 45836 23004
rect 45888 22992 45894 23044
rect 40175 22936 41000 22964
rect 43073 22967 43131 22973
rect 40175 22933 40187 22936
rect 40129 22927 40187 22933
rect 43073 22933 43085 22967
rect 43119 22964 43131 22967
rect 43530 22964 43536 22976
rect 43119 22936 43536 22964
rect 43119 22933 43131 22936
rect 43073 22927 43131 22933
rect 43530 22924 43536 22936
rect 43588 22964 43594 22976
rect 44269 22967 44327 22973
rect 44269 22964 44281 22967
rect 43588 22936 44281 22964
rect 43588 22924 43594 22936
rect 44269 22933 44281 22936
rect 44315 22933 44327 22967
rect 44269 22927 44327 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 11422 22720 11428 22772
rect 11480 22760 11486 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 11480 22732 11713 22760
rect 11480 22720 11486 22732
rect 11701 22729 11713 22732
rect 11747 22729 11759 22763
rect 11701 22723 11759 22729
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12529 22763 12587 22769
rect 12529 22760 12541 22763
rect 12492 22732 12541 22760
rect 12492 22720 12498 22732
rect 12529 22729 12541 22732
rect 12575 22729 12587 22763
rect 12529 22723 12587 22729
rect 18414 22720 18420 22772
rect 18472 22760 18478 22772
rect 18969 22763 19027 22769
rect 18969 22760 18981 22763
rect 18472 22732 18981 22760
rect 18472 22720 18478 22732
rect 18969 22729 18981 22732
rect 19015 22729 19027 22763
rect 19242 22760 19248 22772
rect 19203 22732 19248 22760
rect 18969 22723 19027 22729
rect 19242 22720 19248 22732
rect 19300 22720 19306 22772
rect 27706 22760 27712 22772
rect 27667 22732 27712 22760
rect 27706 22720 27712 22732
rect 27764 22720 27770 22772
rect 30190 22720 30196 22772
rect 30248 22760 30254 22772
rect 30466 22760 30472 22772
rect 30248 22732 30472 22760
rect 30248 22720 30254 22732
rect 30466 22720 30472 22732
rect 30524 22760 30530 22772
rect 31846 22760 31852 22772
rect 30524 22732 31852 22760
rect 30524 22720 30530 22732
rect 31846 22720 31852 22732
rect 31904 22760 31910 22772
rect 33873 22763 33931 22769
rect 33873 22760 33885 22763
rect 31904 22732 33885 22760
rect 31904 22720 31910 22732
rect 33873 22729 33885 22732
rect 33919 22729 33931 22763
rect 33873 22723 33931 22729
rect 39758 22720 39764 22772
rect 39816 22760 39822 22772
rect 39853 22763 39911 22769
rect 39853 22760 39865 22763
rect 39816 22732 39865 22760
rect 39816 22720 39822 22732
rect 39853 22729 39865 22732
rect 39899 22729 39911 22763
rect 40678 22760 40684 22772
rect 40639 22732 40684 22760
rect 39853 22723 39911 22729
rect 40678 22720 40684 22732
rect 40736 22720 40742 22772
rect 45646 22720 45652 22772
rect 45704 22760 45710 22772
rect 47578 22760 47584 22772
rect 45704 22732 47584 22760
rect 45704 22720 45710 22732
rect 47578 22720 47584 22732
rect 47636 22760 47642 22772
rect 47765 22763 47823 22769
rect 47765 22760 47777 22763
rect 47636 22732 47777 22760
rect 47636 22720 47642 22732
rect 47765 22729 47777 22732
rect 47811 22729 47823 22763
rect 47765 22723 47823 22729
rect 3510 22652 3516 22704
rect 3568 22692 3574 22704
rect 20809 22695 20867 22701
rect 3568 22664 19196 22692
rect 3568 22652 3574 22664
rect 9950 22624 9956 22636
rect 9911 22596 9956 22624
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 10827 22596 11284 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 10045 22559 10103 22565
rect 10045 22525 10057 22559
rect 10091 22556 10103 22559
rect 11146 22556 11152 22568
rect 10091 22528 11152 22556
rect 10091 22525 10103 22528
rect 10045 22519 10103 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 11256 22488 11284 22596
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 11388 22596 11529 22624
rect 11388 22584 11394 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 11517 22587 11575 22593
rect 11532 22556 11560 22587
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 12492 22596 12537 22624
rect 12492 22584 12498 22596
rect 13170 22584 13176 22636
rect 13228 22624 13234 22636
rect 13633 22627 13691 22633
rect 13633 22624 13645 22627
rect 13228 22596 13645 22624
rect 13228 22584 13234 22596
rect 13633 22593 13645 22596
rect 13679 22593 13691 22627
rect 17402 22624 17408 22636
rect 17363 22596 17408 22624
rect 13633 22587 13691 22593
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18472 22596 18889 22624
rect 18472 22584 18478 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 19061 22627 19119 22633
rect 19061 22593 19073 22627
rect 19107 22593 19119 22627
rect 19061 22587 19119 22593
rect 12802 22556 12808 22568
rect 11532 22528 12808 22556
rect 12802 22516 12808 22528
rect 12860 22516 12866 22568
rect 13814 22556 13820 22568
rect 13775 22528 13820 22556
rect 13814 22516 13820 22528
rect 13872 22516 13878 22568
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22556 15531 22559
rect 15562 22556 15568 22568
rect 15519 22528 15568 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 15562 22516 15568 22528
rect 15620 22516 15626 22568
rect 18690 22556 18696 22568
rect 18651 22528 18696 22556
rect 18690 22516 18696 22528
rect 18748 22516 18754 22568
rect 12434 22488 12440 22500
rect 11256 22460 12440 22488
rect 12434 22448 12440 22460
rect 12492 22448 12498 22500
rect 18322 22448 18328 22500
rect 18380 22488 18386 22500
rect 19076 22488 19104 22587
rect 18380 22460 19104 22488
rect 19168 22488 19196 22664
rect 20809 22661 20821 22695
rect 20855 22692 20867 22695
rect 22005 22695 22063 22701
rect 22005 22692 22017 22695
rect 20855 22664 22017 22692
rect 20855 22661 20867 22664
rect 20809 22655 20867 22661
rect 22005 22661 22017 22664
rect 22051 22661 22063 22695
rect 22005 22655 22063 22661
rect 23661 22695 23719 22701
rect 23661 22661 23673 22695
rect 23707 22692 23719 22695
rect 27890 22692 27896 22704
rect 23707 22664 27896 22692
rect 23707 22661 23719 22664
rect 23661 22655 23719 22661
rect 27890 22652 27896 22664
rect 27948 22652 27954 22704
rect 28905 22695 28963 22701
rect 28905 22661 28917 22695
rect 28951 22692 28963 22695
rect 29546 22692 29552 22704
rect 28951 22664 29552 22692
rect 28951 22661 28963 22664
rect 28905 22655 28963 22661
rect 29546 22652 29552 22664
rect 29604 22692 29610 22704
rect 30282 22692 30288 22704
rect 29604 22664 30288 22692
rect 29604 22652 29610 22664
rect 30282 22652 30288 22664
rect 30340 22652 30346 22704
rect 31018 22692 31024 22704
rect 30979 22664 31024 22692
rect 31018 22652 31024 22664
rect 31076 22652 31082 22704
rect 31202 22692 31208 22704
rect 31163 22664 31208 22692
rect 31202 22652 31208 22664
rect 31260 22652 31266 22704
rect 48133 22695 48191 22701
rect 48133 22692 48145 22695
rect 41386 22664 48145 22692
rect 20714 22624 20720 22636
rect 20675 22596 20720 22624
rect 20714 22584 20720 22596
rect 20772 22584 20778 22636
rect 26973 22627 27031 22633
rect 26973 22593 26985 22627
rect 27019 22624 27031 22627
rect 27430 22624 27436 22636
rect 27019 22596 27436 22624
rect 27019 22593 27031 22596
rect 26973 22587 27031 22593
rect 27430 22584 27436 22596
rect 27488 22624 27494 22636
rect 27617 22627 27675 22633
rect 27617 22624 27629 22627
rect 27488 22596 27629 22624
rect 27488 22584 27494 22596
rect 27617 22593 27629 22596
rect 27663 22593 27675 22627
rect 28718 22624 28724 22636
rect 28679 22596 28724 22624
rect 27617 22587 27675 22593
rect 28718 22584 28724 22596
rect 28776 22584 28782 22636
rect 28997 22627 29055 22633
rect 28997 22593 29009 22627
rect 29043 22593 29055 22627
rect 28997 22587 29055 22593
rect 21821 22559 21879 22565
rect 21821 22525 21833 22559
rect 21867 22556 21879 22559
rect 22002 22556 22008 22568
rect 21867 22528 22008 22556
rect 21867 22525 21879 22528
rect 21821 22519 21879 22525
rect 22002 22516 22008 22528
rect 22060 22516 22066 22568
rect 24118 22556 24124 22568
rect 24079 22528 24124 22556
rect 24118 22516 24124 22528
rect 24176 22516 24182 22568
rect 24302 22556 24308 22568
rect 24263 22528 24308 22556
rect 24302 22516 24308 22528
rect 24360 22516 24366 22568
rect 24581 22559 24639 22565
rect 24581 22525 24593 22559
rect 24627 22525 24639 22559
rect 29012 22556 29040 22587
rect 29086 22584 29092 22636
rect 29144 22624 29150 22636
rect 30009 22627 30067 22633
rect 30009 22624 30021 22627
rect 29144 22596 29189 22624
rect 29288 22596 30021 22624
rect 29144 22584 29150 22596
rect 29288 22556 29316 22596
rect 30009 22593 30021 22596
rect 30055 22624 30067 22627
rect 30374 22624 30380 22636
rect 30055 22596 30380 22624
rect 30055 22593 30067 22596
rect 30009 22587 30067 22593
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 32030 22584 32036 22636
rect 32088 22624 32094 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 32088 22596 32137 22624
rect 32088 22584 32094 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 33502 22584 33508 22636
rect 33560 22584 33566 22636
rect 40126 22584 40132 22636
rect 40184 22624 40190 22636
rect 40221 22627 40279 22633
rect 40221 22624 40233 22627
rect 40184 22596 40233 22624
rect 40184 22584 40190 22596
rect 40221 22593 40233 22596
rect 40267 22624 40279 22627
rect 41386 22624 41414 22664
rect 48133 22661 48145 22664
rect 48179 22661 48191 22695
rect 48133 22655 48191 22661
rect 40267 22596 41414 22624
rect 44913 22627 44971 22633
rect 40267 22593 40279 22596
rect 40221 22587 40279 22593
rect 44913 22593 44925 22627
rect 44959 22593 44971 22627
rect 44913 22587 44971 22593
rect 29730 22556 29736 22568
rect 29012 22528 29316 22556
rect 29691 22528 29736 22556
rect 24581 22519 24639 22525
rect 24596 22488 24624 22519
rect 29730 22516 29736 22528
rect 29788 22516 29794 22568
rect 31754 22516 31760 22568
rect 31812 22556 31818 22568
rect 32401 22559 32459 22565
rect 32401 22556 32413 22559
rect 31812 22528 32413 22556
rect 31812 22516 31818 22528
rect 32401 22525 32413 22528
rect 32447 22525 32459 22559
rect 44928 22556 44956 22587
rect 45278 22584 45284 22636
rect 45336 22624 45342 22636
rect 45373 22627 45431 22633
rect 45373 22624 45385 22627
rect 45336 22596 45385 22624
rect 45336 22584 45342 22596
rect 45373 22593 45385 22596
rect 45419 22593 45431 22627
rect 45373 22587 45431 22593
rect 45557 22627 45615 22633
rect 45557 22593 45569 22627
rect 45603 22624 45615 22627
rect 45646 22624 45652 22636
rect 45603 22596 45652 22624
rect 45603 22593 45615 22596
rect 45557 22587 45615 22593
rect 45646 22584 45652 22596
rect 45704 22584 45710 22636
rect 47854 22624 47860 22636
rect 47815 22596 47860 22624
rect 47854 22584 47860 22596
rect 47912 22584 47918 22636
rect 47949 22627 48007 22633
rect 47949 22593 47961 22627
rect 47995 22624 48007 22627
rect 48038 22624 48044 22636
rect 47995 22596 48044 22624
rect 47995 22593 48007 22596
rect 47949 22587 48007 22593
rect 48038 22584 48044 22596
rect 48096 22584 48102 22636
rect 46014 22556 46020 22568
rect 44928 22528 46020 22556
rect 32401 22519 32459 22525
rect 46014 22516 46020 22528
rect 46072 22516 46078 22568
rect 46198 22556 46204 22568
rect 46159 22528 46204 22556
rect 46198 22516 46204 22528
rect 46256 22516 46262 22568
rect 46477 22559 46535 22565
rect 46477 22525 46489 22559
rect 46523 22525 46535 22559
rect 46477 22519 46535 22525
rect 47581 22559 47639 22565
rect 47581 22525 47593 22559
rect 47627 22556 47639 22559
rect 47762 22556 47768 22568
rect 47627 22528 47768 22556
rect 47627 22525 47639 22528
rect 47581 22519 47639 22525
rect 19168 22460 24624 22488
rect 18380 22448 18386 22460
rect 44266 22448 44272 22500
rect 44324 22488 44330 22500
rect 46492 22488 46520 22519
rect 47762 22516 47768 22528
rect 47820 22516 47826 22568
rect 44324 22460 46520 22488
rect 44324 22448 44330 22460
rect 10318 22420 10324 22432
rect 10279 22392 10324 22420
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 10873 22423 10931 22429
rect 10873 22389 10885 22423
rect 10919 22420 10931 22423
rect 11054 22420 11060 22432
rect 10919 22392 11060 22420
rect 10919 22389 10931 22392
rect 10873 22383 10931 22389
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 17497 22423 17555 22429
rect 17497 22389 17509 22423
rect 17543 22420 17555 22423
rect 17954 22420 17960 22432
rect 17543 22392 17960 22420
rect 17543 22389 17555 22392
rect 17497 22383 17555 22389
rect 17954 22380 17960 22392
rect 18012 22380 18018 22432
rect 27062 22420 27068 22432
rect 27023 22392 27068 22420
rect 27062 22380 27068 22392
rect 27120 22380 27126 22432
rect 29270 22420 29276 22432
rect 29231 22392 29276 22420
rect 29270 22380 29276 22392
rect 29328 22380 29334 22432
rect 31389 22423 31447 22429
rect 31389 22389 31401 22423
rect 31435 22420 31447 22423
rect 31938 22420 31944 22432
rect 31435 22392 31944 22420
rect 31435 22389 31447 22392
rect 31389 22383 31447 22389
rect 31938 22380 31944 22392
rect 31996 22380 32002 22432
rect 39758 22380 39764 22432
rect 39816 22420 39822 22432
rect 40310 22420 40316 22432
rect 39816 22392 40316 22420
rect 39816 22380 39822 22392
rect 40310 22380 40316 22392
rect 40368 22380 40374 22432
rect 44729 22423 44787 22429
rect 44729 22389 44741 22423
rect 44775 22420 44787 22423
rect 45646 22420 45652 22432
rect 44775 22392 45652 22420
rect 44775 22389 44787 22392
rect 44729 22383 44787 22389
rect 45646 22380 45652 22392
rect 45704 22380 45710 22432
rect 45738 22380 45744 22432
rect 45796 22420 45802 22432
rect 45796 22392 45841 22420
rect 45796 22380 45802 22392
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 10318 22176 10324 22228
rect 10376 22216 10382 22228
rect 10486 22219 10544 22225
rect 10486 22216 10498 22219
rect 10376 22188 10498 22216
rect 10376 22176 10382 22188
rect 10486 22185 10498 22188
rect 10532 22185 10544 22219
rect 10486 22179 10544 22185
rect 16840 22219 16898 22225
rect 16840 22185 16852 22219
rect 16886 22216 16898 22219
rect 18046 22216 18052 22228
rect 16886 22188 18052 22216
rect 16886 22185 16898 22188
rect 16840 22179 16898 22185
rect 18046 22176 18052 22188
rect 18104 22176 18110 22228
rect 25764 22219 25822 22225
rect 25764 22185 25776 22219
rect 25810 22216 25822 22219
rect 25866 22216 25872 22228
rect 25810 22188 25872 22216
rect 25810 22185 25822 22188
rect 25764 22179 25822 22185
rect 25866 22176 25872 22188
rect 25924 22176 25930 22228
rect 43070 22216 43076 22228
rect 38626 22188 41414 22216
rect 43031 22188 43076 22216
rect 9950 22108 9956 22160
rect 10008 22148 10014 22160
rect 12713 22151 12771 22157
rect 10008 22120 10364 22148
rect 10008 22108 10014 22120
rect 10226 22080 10232 22092
rect 10187 22052 10232 22080
rect 10226 22040 10232 22052
rect 10284 22040 10290 22092
rect 10336 22080 10364 22120
rect 12713 22117 12725 22151
rect 12759 22148 12771 22151
rect 12802 22148 12808 22160
rect 12759 22120 12808 22148
rect 12759 22117 12771 22120
rect 12713 22111 12771 22117
rect 12802 22108 12808 22120
rect 12860 22108 12866 22160
rect 29086 22108 29092 22160
rect 29144 22148 29150 22160
rect 38626 22148 38654 22188
rect 29144 22120 38654 22148
rect 41386 22148 41414 22188
rect 43070 22176 43076 22188
rect 43128 22176 43134 22228
rect 42886 22148 42892 22160
rect 41386 22120 42892 22148
rect 29144 22108 29150 22120
rect 42886 22108 42892 22120
rect 42944 22108 42950 22160
rect 11974 22080 11980 22092
rect 10336 22052 11980 22080
rect 11974 22040 11980 22052
rect 12032 22040 12038 22092
rect 13449 22083 13507 22089
rect 13449 22049 13461 22083
rect 13495 22080 13507 22083
rect 13814 22080 13820 22092
rect 13495 22052 13820 22080
rect 13495 22049 13507 22052
rect 13449 22043 13507 22049
rect 13814 22040 13820 22052
rect 13872 22040 13878 22092
rect 16114 22080 16120 22092
rect 16075 22052 16120 22080
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 18414 22040 18420 22092
rect 18472 22080 18478 22092
rect 20898 22080 20904 22092
rect 18472 22052 19656 22080
rect 20859 22052 20904 22080
rect 18472 22040 18478 22052
rect 8938 22012 8944 22024
rect 8851 21984 8944 22012
rect 8938 21972 8944 21984
rect 8996 22012 9002 22024
rect 9585 22015 9643 22021
rect 9585 22012 9597 22015
rect 8996 21984 9597 22012
rect 8996 21972 9002 21984
rect 9585 21981 9597 21984
rect 9631 22012 9643 22015
rect 12526 22012 12532 22024
rect 9631 21984 10088 22012
rect 12487 21984 12532 22012
rect 9631 21981 9643 21984
rect 9585 21975 9643 21981
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 9033 21879 9091 21885
rect 9033 21876 9045 21879
rect 8904 21848 9045 21876
rect 8904 21836 8910 21848
rect 9033 21845 9045 21848
rect 9079 21845 9091 21879
rect 9033 21839 9091 21845
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 9677 21879 9735 21885
rect 9677 21876 9689 21879
rect 9180 21848 9689 21876
rect 9180 21836 9186 21848
rect 9677 21845 9689 21848
rect 9723 21845 9735 21879
rect 10060 21876 10088 21984
rect 12526 21972 12532 21984
rect 12584 21972 12590 22024
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 22012 13415 22015
rect 13906 22012 13912 22024
rect 13403 21984 13912 22012
rect 13403 21981 13415 21984
rect 13357 21975 13415 21981
rect 11054 21904 11060 21956
rect 11112 21904 11118 21956
rect 13372 21944 13400 21975
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14274 22012 14280 22024
rect 14235 21984 14280 22012
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 16574 22012 16580 22024
rect 16535 21984 16580 22012
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 17954 21972 17960 22024
rect 18012 21972 18018 22024
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 18782 22012 18788 22024
rect 18380 21984 18788 22012
rect 18380 21972 18386 21984
rect 18782 21972 18788 21984
rect 18840 22012 18846 22024
rect 19521 22015 19579 22021
rect 19521 22012 19533 22015
rect 18840 21984 19533 22012
rect 18840 21972 18846 21984
rect 19521 21981 19533 21984
rect 19567 21981 19579 22015
rect 19521 21975 19579 21981
rect 12406 21916 13400 21944
rect 14461 21947 14519 21953
rect 12406 21876 12434 21916
rect 14461 21913 14473 21947
rect 14507 21944 14519 21947
rect 14642 21944 14648 21956
rect 14507 21916 14648 21944
rect 14507 21913 14519 21916
rect 14461 21907 14519 21913
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 18690 21904 18696 21956
rect 18748 21944 18754 21956
rect 19242 21944 19248 21956
rect 18748 21916 19248 21944
rect 18748 21904 18754 21916
rect 19242 21904 19248 21916
rect 19300 21904 19306 21956
rect 19429 21947 19487 21953
rect 19429 21913 19441 21947
rect 19475 21944 19487 21947
rect 19628 21944 19656 22052
rect 20898 22040 20904 22052
rect 20956 22040 20962 22092
rect 23293 22083 23351 22089
rect 23293 22049 23305 22083
rect 23339 22080 23351 22083
rect 24302 22080 24308 22092
rect 23339 22052 24308 22080
rect 23339 22049 23351 22052
rect 23293 22043 23351 22049
rect 24302 22040 24308 22052
rect 24360 22040 24366 22092
rect 27249 22083 27307 22089
rect 27249 22049 27261 22083
rect 27295 22080 27307 22083
rect 27614 22080 27620 22092
rect 27295 22052 27620 22080
rect 27295 22049 27307 22052
rect 27249 22043 27307 22049
rect 27614 22040 27620 22052
rect 27672 22040 27678 22092
rect 28997 22083 29055 22089
rect 28997 22080 29009 22083
rect 28184 22052 29009 22080
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 22012 20867 22015
rect 21450 22012 21456 22024
rect 20855 21984 21456 22012
rect 20855 21981 20867 21984
rect 20809 21975 20867 21981
rect 21450 21972 21456 21984
rect 21508 21972 21514 22024
rect 23198 22012 23204 22024
rect 23159 21984 23204 22012
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 25498 22012 25504 22024
rect 25459 21984 25504 22012
rect 25498 21972 25504 21984
rect 25556 21972 25562 22024
rect 28184 22021 28212 22052
rect 28997 22049 29009 22052
rect 29043 22049 29055 22083
rect 28997 22043 29055 22049
rect 45554 22040 45560 22092
rect 45612 22080 45618 22092
rect 45741 22083 45799 22089
rect 45741 22080 45753 22083
rect 45612 22052 45753 22080
rect 45612 22040 45618 22052
rect 45741 22049 45753 22052
rect 45787 22049 45799 22083
rect 46934 22080 46940 22092
rect 46895 22052 46940 22080
rect 45741 22043 45799 22049
rect 46934 22040 46940 22052
rect 46992 22040 46998 22092
rect 28169 22015 28227 22021
rect 28169 21981 28181 22015
rect 28215 21981 28227 22015
rect 28169 21975 28227 21981
rect 28629 22015 28687 22021
rect 28629 21981 28641 22015
rect 28675 22012 28687 22015
rect 29270 22012 29276 22024
rect 28675 21984 29276 22012
rect 28675 21981 28687 21984
rect 28629 21975 28687 21981
rect 29270 21972 29276 21984
rect 29328 21972 29334 22024
rect 31938 22012 31944 22024
rect 31899 21984 31944 22012
rect 31938 21972 31944 21984
rect 31996 21972 32002 22024
rect 33870 21972 33876 22024
rect 33928 22012 33934 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 33928 21984 34897 22012
rect 33928 21972 33934 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 40126 22012 40132 22024
rect 40087 21984 40132 22012
rect 34885 21975 34943 21981
rect 40126 21972 40132 21984
rect 40184 21972 40190 22024
rect 40310 22012 40316 22024
rect 40271 21984 40316 22012
rect 40310 21972 40316 21984
rect 40368 21972 40374 22024
rect 43349 22015 43407 22021
rect 43349 21981 43361 22015
rect 43395 22012 43407 22015
rect 43438 22012 43444 22024
rect 43395 21984 43444 22012
rect 43395 21981 43407 21984
rect 43349 21975 43407 21981
rect 43438 21972 43444 21984
rect 43496 21972 43502 22024
rect 45097 22015 45155 22021
rect 45097 21981 45109 22015
rect 45143 22012 45155 22015
rect 45186 22012 45192 22024
rect 45143 21984 45192 22012
rect 45143 21981 45155 21984
rect 45097 21975 45155 21981
rect 45186 21972 45192 21984
rect 45244 21972 45250 22024
rect 45281 22015 45339 22021
rect 45281 21981 45293 22015
rect 45327 22012 45339 22015
rect 45327 21984 45600 22012
rect 45327 21981 45339 21984
rect 45281 21975 45339 21981
rect 27062 21944 27068 21956
rect 19475 21916 19656 21944
rect 27002 21916 27068 21944
rect 19475 21913 19487 21916
rect 19429 21907 19487 21913
rect 27062 21904 27068 21916
rect 27120 21904 27126 21956
rect 28810 21944 28816 21956
rect 28771 21916 28816 21944
rect 28810 21904 28816 21916
rect 28868 21904 28874 21956
rect 40497 21947 40555 21953
rect 40497 21913 40509 21947
rect 40543 21944 40555 21947
rect 40586 21944 40592 21956
rect 40543 21916 40592 21944
rect 40543 21913 40555 21916
rect 40497 21907 40555 21913
rect 40586 21904 40592 21916
rect 40644 21904 40650 21956
rect 43070 21944 43076 21956
rect 43031 21916 43076 21944
rect 43070 21904 43076 21916
rect 43128 21904 43134 21956
rect 10060 21848 12434 21876
rect 18325 21879 18383 21885
rect 9677 21839 9735 21845
rect 18325 21845 18337 21879
rect 18371 21876 18383 21879
rect 18414 21876 18420 21888
rect 18371 21848 18420 21876
rect 18371 21845 18383 21848
rect 18325 21839 18383 21845
rect 18414 21836 18420 21848
rect 18472 21836 18478 21888
rect 18506 21836 18512 21888
rect 18564 21876 18570 21888
rect 19343 21879 19401 21885
rect 19343 21876 19355 21879
rect 18564 21848 19355 21876
rect 18564 21836 18570 21848
rect 19343 21845 19355 21848
rect 19389 21845 19401 21879
rect 19343 21839 19401 21845
rect 27706 21836 27712 21888
rect 27764 21876 27770 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 27764 21848 27997 21876
rect 27764 21836 27770 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 31754 21876 31760 21888
rect 31715 21848 31760 21876
rect 27985 21839 28043 21845
rect 31754 21836 31760 21848
rect 31812 21836 31818 21888
rect 34514 21836 34520 21888
rect 34572 21876 34578 21888
rect 34701 21879 34759 21885
rect 34701 21876 34713 21879
rect 34572 21848 34713 21876
rect 34572 21836 34578 21848
rect 34701 21845 34713 21848
rect 34747 21845 34759 21879
rect 34701 21839 34759 21845
rect 43257 21879 43315 21885
rect 43257 21845 43269 21879
rect 43303 21876 43315 21879
rect 43346 21876 43352 21888
rect 43303 21848 43352 21876
rect 43303 21845 43315 21848
rect 43257 21839 43315 21845
rect 43346 21836 43352 21848
rect 43404 21836 43410 21888
rect 45278 21876 45284 21888
rect 45239 21848 45284 21876
rect 45278 21836 45284 21848
rect 45336 21836 45342 21888
rect 45462 21836 45468 21888
rect 45520 21876 45526 21888
rect 45572 21876 45600 21984
rect 45646 21904 45652 21956
rect 45704 21944 45710 21956
rect 45925 21947 45983 21953
rect 45925 21944 45937 21947
rect 45704 21916 45937 21944
rect 45704 21904 45710 21916
rect 45925 21913 45937 21916
rect 45971 21913 45983 21947
rect 45925 21907 45983 21913
rect 47762 21876 47768 21888
rect 45520 21848 47768 21876
rect 45520 21836 45526 21848
rect 47762 21836 47768 21848
rect 47820 21836 47826 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 10962 21672 10968 21684
rect 8680 21644 10968 21672
rect 14 21564 20 21616
rect 72 21604 78 21616
rect 72 21576 2774 21604
rect 72 21564 78 21576
rect 2746 21400 2774 21576
rect 8680 21545 8708 21644
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 14642 21672 14648 21684
rect 14603 21644 14648 21672
rect 14642 21632 14648 21644
rect 14700 21632 14706 21684
rect 16666 21632 16672 21684
rect 16724 21672 16730 21684
rect 16853 21675 16911 21681
rect 16853 21672 16865 21675
rect 16724 21644 16865 21672
rect 16724 21632 16730 21644
rect 16853 21641 16865 21644
rect 16899 21641 16911 21675
rect 16853 21635 16911 21641
rect 17144 21644 20944 21672
rect 8846 21604 8852 21616
rect 8807 21576 8852 21604
rect 8846 21564 8852 21576
rect 8904 21564 8910 21616
rect 12526 21564 12532 21616
rect 12584 21604 12590 21616
rect 13722 21604 13728 21616
rect 12584 21576 13728 21604
rect 12584 21564 12590 21576
rect 13722 21564 13728 21576
rect 13780 21604 13786 21616
rect 13780 21576 16712 21604
rect 13780 21564 13786 21576
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 13906 21496 13912 21548
rect 13964 21536 13970 21548
rect 16684 21545 16712 21576
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 13964 21508 14565 21536
rect 13964 21496 13970 21508
rect 14553 21505 14565 21508
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 17144 21536 17172 21644
rect 18414 21604 18420 21616
rect 17604 21576 18420 21604
rect 17604 21545 17632 21576
rect 18414 21564 18420 21576
rect 18472 21564 18478 21616
rect 20916 21613 20944 21644
rect 28718 21632 28724 21684
rect 28776 21672 28782 21684
rect 29181 21675 29239 21681
rect 29181 21672 29193 21675
rect 28776 21644 29193 21672
rect 28776 21632 28782 21644
rect 29181 21641 29193 21644
rect 29227 21641 29239 21675
rect 33870 21672 33876 21684
rect 33831 21644 33876 21672
rect 29181 21635 29239 21641
rect 33870 21632 33876 21644
rect 33928 21632 33934 21684
rect 42886 21632 42892 21684
rect 42944 21672 42950 21684
rect 42944 21644 45876 21672
rect 42944 21632 42950 21644
rect 20901 21607 20959 21613
rect 20901 21573 20913 21607
rect 20947 21604 20959 21607
rect 21818 21604 21824 21616
rect 20947 21576 21824 21604
rect 20947 21573 20959 21576
rect 20901 21567 20959 21573
rect 21818 21564 21824 21576
rect 21876 21564 21882 21616
rect 23201 21607 23259 21613
rect 23201 21573 23213 21607
rect 23247 21604 23259 21607
rect 23474 21604 23480 21616
rect 23247 21576 23480 21604
rect 23247 21573 23259 21576
rect 23201 21567 23259 21573
rect 23474 21564 23480 21576
rect 23532 21564 23538 21616
rect 27706 21604 27712 21616
rect 27667 21576 27712 21604
rect 27706 21564 27712 21576
rect 27764 21564 27770 21616
rect 28166 21564 28172 21616
rect 28224 21564 28230 21616
rect 34422 21604 34428 21616
rect 34383 21576 34428 21604
rect 34422 21564 34428 21576
rect 34480 21564 34486 21616
rect 34514 21564 34520 21616
rect 34572 21604 34578 21616
rect 42521 21607 42579 21613
rect 34572 21576 34617 21604
rect 34572 21564 34578 21576
rect 42521 21573 42533 21607
rect 42567 21604 42579 21607
rect 43070 21604 43076 21616
rect 42567 21576 43076 21604
rect 42567 21573 42579 21576
rect 42521 21567 42579 21573
rect 43070 21564 43076 21576
rect 43128 21564 43134 21616
rect 45554 21604 45560 21616
rect 44836 21576 45560 21604
rect 16715 21508 17172 21536
rect 17589 21539 17647 21545
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 17589 21505 17601 21539
rect 17635 21505 17647 21539
rect 18322 21536 18328 21548
rect 17589 21499 17647 21505
rect 17696 21508 18328 21536
rect 17696 21477 17724 21508
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 18506 21536 18512 21548
rect 18467 21508 18512 21536
rect 18506 21496 18512 21508
rect 18564 21496 18570 21548
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 20162 21536 20168 21548
rect 18739 21508 20168 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 20162 21496 20168 21508
rect 20220 21496 20226 21548
rect 22189 21539 22247 21545
rect 22189 21505 22201 21539
rect 22235 21536 22247 21539
rect 22235 21508 23060 21536
rect 22235 21505 22247 21508
rect 22189 21499 22247 21505
rect 23032 21480 23060 21508
rect 25498 21496 25504 21548
rect 25556 21536 25562 21548
rect 27433 21539 27491 21545
rect 27433 21536 27445 21539
rect 25556 21508 27445 21536
rect 25556 21496 25562 21508
rect 27433 21505 27445 21508
rect 27479 21505 27491 21539
rect 27433 21499 27491 21505
rect 33413 21539 33471 21545
rect 33413 21505 33425 21539
rect 33459 21505 33471 21539
rect 33413 21499 33471 21505
rect 9125 21471 9183 21477
rect 9125 21437 9137 21471
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 17681 21471 17739 21477
rect 17681 21437 17693 21471
rect 17727 21437 17739 21471
rect 17681 21431 17739 21437
rect 17957 21471 18015 21477
rect 17957 21437 17969 21471
rect 18003 21468 18015 21471
rect 18046 21468 18052 21480
rect 18003 21440 18052 21468
rect 18003 21437 18015 21440
rect 17957 21431 18015 21437
rect 9140 21400 9168 21431
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 22278 21468 22284 21480
rect 22239 21440 22284 21468
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 23014 21468 23020 21480
rect 22975 21440 23020 21468
rect 23014 21428 23020 21440
rect 23072 21428 23078 21480
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21437 23535 21471
rect 23477 21431 23535 21437
rect 23492 21400 23520 21431
rect 2746 21372 9168 21400
rect 12406 21372 23520 21400
rect 33428 21400 33456 21499
rect 42334 21496 42340 21548
rect 42392 21536 42398 21548
rect 42429 21539 42487 21545
rect 42429 21536 42441 21539
rect 42392 21508 42441 21536
rect 42392 21496 42398 21508
rect 42429 21505 42441 21508
rect 42475 21505 42487 21539
rect 42429 21499 42487 21505
rect 42613 21539 42671 21545
rect 42613 21505 42625 21539
rect 42659 21505 42671 21539
rect 42613 21499 42671 21505
rect 42628 21468 42656 21499
rect 42702 21496 42708 21548
rect 42760 21536 42766 21548
rect 43993 21539 44051 21545
rect 43993 21536 44005 21539
rect 42760 21508 44005 21536
rect 42760 21496 42766 21508
rect 43993 21505 44005 21508
rect 44039 21505 44051 21539
rect 43993 21499 44051 21505
rect 44174 21496 44180 21548
rect 44232 21536 44238 21548
rect 44836 21545 44864 21576
rect 45554 21564 45560 21576
rect 45612 21564 45618 21616
rect 45848 21604 45876 21644
rect 46014 21632 46020 21684
rect 46072 21672 46078 21684
rect 48133 21675 48191 21681
rect 48133 21672 48145 21675
rect 46072 21644 48145 21672
rect 46072 21632 46078 21644
rect 48133 21641 48145 21644
rect 48179 21641 48191 21675
rect 48133 21635 48191 21641
rect 45848 21576 46520 21604
rect 44821 21539 44879 21545
rect 44232 21508 44325 21536
rect 44232 21496 44238 21508
rect 44821 21505 44833 21539
rect 44867 21505 44879 21539
rect 44821 21499 44879 21505
rect 45186 21496 45192 21548
rect 45244 21536 45250 21548
rect 45281 21539 45339 21545
rect 45281 21536 45293 21539
rect 45244 21508 45293 21536
rect 45244 21496 45250 21508
rect 45281 21505 45293 21508
rect 45327 21505 45339 21539
rect 46198 21536 46204 21548
rect 46159 21508 46204 21536
rect 45281 21499 45339 21505
rect 44192 21468 44220 21496
rect 42628 21440 44220 21468
rect 45296 21468 45324 21499
rect 46198 21496 46204 21508
rect 46256 21496 46262 21548
rect 46492 21545 46520 21576
rect 46477 21539 46535 21545
rect 46477 21505 46489 21539
rect 46523 21505 46535 21539
rect 47578 21536 47584 21548
rect 47539 21508 47584 21536
rect 46477 21499 46535 21505
rect 47578 21496 47584 21508
rect 47636 21496 47642 21548
rect 48038 21536 48044 21548
rect 47688 21508 48044 21536
rect 47688 21468 47716 21508
rect 48038 21496 48044 21508
rect 48096 21496 48102 21548
rect 47854 21468 47860 21480
rect 45296 21440 47716 21468
rect 47815 21440 47860 21468
rect 47854 21428 47860 21440
rect 47912 21428 47918 21480
rect 34977 21403 35035 21409
rect 33428 21372 34652 21400
rect 3786 21292 3792 21344
rect 3844 21332 3850 21344
rect 12406 21332 12434 21372
rect 18506 21332 18512 21344
rect 3844 21304 12434 21332
rect 18467 21304 18512 21332
rect 3844 21292 3850 21304
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 20990 21332 20996 21344
rect 20951 21304 20996 21332
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 22370 21292 22376 21344
rect 22428 21332 22434 21344
rect 22557 21335 22615 21341
rect 22557 21332 22569 21335
rect 22428 21304 22569 21332
rect 22428 21292 22434 21304
rect 22557 21301 22569 21304
rect 22603 21301 22615 21335
rect 22557 21295 22615 21301
rect 33689 21335 33747 21341
rect 33689 21301 33701 21335
rect 33735 21332 33747 21335
rect 34238 21332 34244 21344
rect 33735 21304 34244 21332
rect 33735 21301 33747 21304
rect 33689 21295 33747 21301
rect 34238 21292 34244 21304
rect 34296 21292 34302 21344
rect 34624 21332 34652 21372
rect 34977 21369 34989 21403
rect 35023 21400 35035 21403
rect 35802 21400 35808 21412
rect 35023 21372 35808 21400
rect 35023 21369 35035 21372
rect 34977 21363 35035 21369
rect 35802 21360 35808 21372
rect 35860 21400 35866 21412
rect 42794 21400 42800 21412
rect 35860 21372 42800 21400
rect 35860 21360 35866 21372
rect 42794 21360 42800 21372
rect 42852 21360 42858 21412
rect 43346 21400 43352 21412
rect 43307 21372 43352 21400
rect 43346 21360 43352 21372
rect 43404 21400 43410 21412
rect 44085 21403 44143 21409
rect 44085 21400 44097 21403
rect 43404 21372 44097 21400
rect 43404 21360 43410 21372
rect 44085 21369 44097 21372
rect 44131 21369 44143 21403
rect 44085 21363 44143 21369
rect 45278 21360 45284 21412
rect 45336 21400 45342 21412
rect 45336 21372 47716 21400
rect 45336 21360 45342 21372
rect 35894 21332 35900 21344
rect 34624 21304 35900 21332
rect 35894 21292 35900 21304
rect 35952 21292 35958 21344
rect 43530 21332 43536 21344
rect 43491 21304 43536 21332
rect 43530 21292 43536 21304
rect 43588 21292 43594 21344
rect 44634 21332 44640 21344
rect 44595 21304 44640 21332
rect 44634 21292 44640 21304
rect 44692 21292 44698 21344
rect 45462 21332 45468 21344
rect 45423 21304 45468 21332
rect 45462 21292 45468 21304
rect 45520 21292 45526 21344
rect 45741 21335 45799 21341
rect 45741 21301 45753 21335
rect 45787 21332 45799 21335
rect 45830 21332 45836 21344
rect 45787 21304 45836 21332
rect 45787 21301 45799 21304
rect 45741 21295 45799 21301
rect 45830 21292 45836 21304
rect 45888 21292 45894 21344
rect 47688 21341 47716 21372
rect 47673 21335 47731 21341
rect 47673 21301 47685 21335
rect 47719 21301 47731 21335
rect 47673 21295 47731 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 16574 21128 16580 21140
rect 16535 21100 16580 21128
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 23014 21088 23020 21140
rect 23072 21128 23078 21140
rect 23845 21131 23903 21137
rect 23845 21128 23857 21131
rect 23072 21100 23857 21128
rect 23072 21088 23078 21100
rect 23845 21097 23857 21100
rect 23891 21097 23903 21131
rect 23845 21091 23903 21097
rect 26605 21131 26663 21137
rect 26605 21097 26617 21131
rect 26651 21128 26663 21131
rect 27430 21128 27436 21140
rect 26651 21100 27436 21128
rect 26651 21097 26663 21100
rect 26605 21091 26663 21097
rect 27430 21088 27436 21100
rect 27488 21088 27494 21140
rect 27617 21131 27675 21137
rect 27617 21097 27629 21131
rect 27663 21128 27675 21131
rect 28166 21128 28172 21140
rect 27663 21100 28172 21128
rect 27663 21097 27675 21100
rect 27617 21091 27675 21097
rect 28166 21088 28172 21100
rect 28224 21088 28230 21140
rect 9950 21060 9956 21072
rect 8956 21032 9956 21060
rect 8956 21001 8984 21032
rect 9950 21020 9956 21032
rect 10008 21020 10014 21072
rect 14277 21063 14335 21069
rect 14277 21029 14289 21063
rect 14323 21060 14335 21063
rect 35802 21060 35808 21072
rect 14323 21032 14872 21060
rect 35763 21032 35808 21060
rect 14323 21029 14335 21032
rect 14277 21023 14335 21029
rect 8941 20995 8999 21001
rect 8941 20961 8953 20995
rect 8987 20961 8999 20995
rect 9122 20992 9128 21004
rect 9083 20964 9128 20992
rect 8941 20955 8999 20961
rect 9122 20952 9128 20964
rect 9180 20952 9186 21004
rect 14844 20936 14872 21032
rect 35802 21020 35808 21032
rect 35860 21020 35866 21072
rect 44266 21060 44272 21072
rect 40696 21032 44272 21060
rect 22370 20992 22376 21004
rect 22331 20964 22376 20992
rect 22370 20952 22376 20964
rect 22428 20952 22434 21004
rect 26786 20952 26792 21004
rect 26844 20992 26850 21004
rect 31665 20995 31723 21001
rect 26844 20964 30604 20992
rect 26844 20952 26850 20964
rect 30576 20936 30604 20964
rect 31665 20961 31677 20995
rect 31711 20992 31723 20995
rect 40696 20992 40724 21032
rect 44266 21020 44272 21032
rect 44324 21020 44330 21072
rect 43438 20992 43444 21004
rect 31711 20964 40724 20992
rect 43399 20964 43444 20992
rect 31711 20961 31723 20964
rect 31665 20955 31723 20961
rect 43438 20952 43444 20964
rect 43496 20952 43502 21004
rect 44082 20992 44088 21004
rect 44043 20964 44088 20992
rect 44082 20952 44088 20964
rect 44140 20952 44146 21004
rect 45189 20995 45247 21001
rect 45189 20961 45201 20995
rect 45235 20992 45247 20995
rect 46293 20995 46351 21001
rect 46293 20992 46305 20995
rect 45235 20964 46305 20992
rect 45235 20961 45247 20964
rect 45189 20955 45247 20961
rect 46293 20961 46305 20964
rect 46339 20961 46351 20995
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 46293 20955 46351 20961
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20893 14151 20927
rect 14826 20924 14832 20936
rect 14787 20896 14832 20924
rect 14093 20887 14151 20893
rect 10778 20856 10784 20868
rect 10739 20828 10784 20856
rect 10778 20816 10784 20828
rect 10836 20816 10842 20868
rect 14108 20856 14136 20887
rect 14826 20884 14832 20896
rect 14884 20884 14890 20936
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20924 16635 20927
rect 16666 20924 16672 20936
rect 16623 20896 16672 20924
rect 16623 20893 16635 20896
rect 16577 20887 16635 20893
rect 16666 20884 16672 20896
rect 16724 20924 16730 20936
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 16724 20896 17417 20924
rect 16724 20884 16730 20896
rect 17405 20893 17417 20896
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 19150 20884 19156 20936
rect 19208 20924 19214 20936
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19208 20896 19257 20924
rect 19208 20884 19214 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 21361 20927 21419 20933
rect 21361 20924 21373 20927
rect 21048 20896 21373 20924
rect 21048 20884 21054 20896
rect 21361 20893 21373 20896
rect 21407 20893 21419 20927
rect 21361 20887 21419 20893
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20924 21695 20927
rect 22097 20927 22155 20933
rect 22097 20924 22109 20927
rect 21683 20896 22109 20924
rect 21683 20893 21695 20896
rect 21637 20887 21695 20893
rect 22097 20893 22109 20896
rect 22143 20893 22155 20927
rect 22097 20887 22155 20893
rect 23474 20884 23480 20936
rect 23532 20884 23538 20936
rect 25958 20884 25964 20936
rect 26016 20924 26022 20936
rect 26421 20927 26479 20933
rect 26421 20924 26433 20927
rect 26016 20896 26433 20924
rect 26016 20884 26022 20896
rect 26421 20893 26433 20896
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 27430 20884 27436 20936
rect 27488 20924 27494 20936
rect 27525 20927 27583 20933
rect 27525 20924 27537 20927
rect 27488 20896 27537 20924
rect 27488 20884 27494 20896
rect 27525 20893 27537 20896
rect 27571 20893 27583 20927
rect 30558 20924 30564 20936
rect 30471 20896 30564 20924
rect 27525 20887 27583 20893
rect 30558 20884 30564 20896
rect 30616 20884 30622 20936
rect 43530 20924 43536 20936
rect 43491 20896 43536 20924
rect 43530 20884 43536 20896
rect 43588 20884 43594 20936
rect 45830 20924 45836 20936
rect 45791 20896 45836 20924
rect 45830 20884 45836 20896
rect 45888 20884 45894 20936
rect 15102 20856 15108 20868
rect 14108 20828 15108 20856
rect 15102 20816 15108 20828
rect 15160 20816 15166 20868
rect 31754 20816 31760 20868
rect 31812 20856 31818 20868
rect 31812 20828 31857 20856
rect 31812 20816 31818 20828
rect 32582 20816 32588 20868
rect 32640 20856 32646 20868
rect 32677 20859 32735 20865
rect 32677 20856 32689 20859
rect 32640 20828 32689 20856
rect 32640 20816 32646 20828
rect 32677 20825 32689 20828
rect 32723 20825 32735 20859
rect 32677 20819 32735 20825
rect 32858 20816 32864 20868
rect 32916 20856 32922 20868
rect 35253 20859 35311 20865
rect 35253 20856 35265 20859
rect 32916 20828 35265 20856
rect 32916 20816 32922 20828
rect 35253 20825 35265 20828
rect 35299 20825 35311 20859
rect 35253 20819 35311 20825
rect 35345 20859 35403 20865
rect 35345 20825 35357 20859
rect 35391 20856 35403 20859
rect 35894 20856 35900 20868
rect 35391 20828 35900 20856
rect 35391 20825 35403 20828
rect 35345 20819 35403 20825
rect 35894 20816 35900 20828
rect 35952 20856 35958 20868
rect 36354 20856 36360 20868
rect 35952 20828 36360 20856
rect 35952 20816 35958 20828
rect 36354 20816 36360 20828
rect 36412 20816 36418 20868
rect 46477 20859 46535 20865
rect 46477 20825 46489 20859
rect 46523 20856 46535 20859
rect 47670 20856 47676 20868
rect 46523 20828 47676 20856
rect 46523 20825 46535 20828
rect 46477 20819 46535 20825
rect 47670 20816 47676 20828
rect 47728 20816 47734 20868
rect 14090 20748 14096 20800
rect 14148 20788 14154 20800
rect 14550 20788 14556 20800
rect 14148 20760 14556 20788
rect 14148 20748 14154 20760
rect 14550 20748 14556 20760
rect 14608 20748 14614 20800
rect 14918 20788 14924 20800
rect 14879 20760 14924 20788
rect 14918 20748 14924 20760
rect 14976 20748 14982 20800
rect 17497 20791 17555 20797
rect 17497 20757 17509 20791
rect 17543 20788 17555 20791
rect 17954 20788 17960 20800
rect 17543 20760 17960 20788
rect 17543 20757 17555 20760
rect 17497 20751 17555 20757
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 19334 20788 19340 20800
rect 19295 20760 19340 20788
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 30650 20788 30656 20800
rect 30611 20760 30656 20788
rect 30650 20748 30656 20760
rect 30708 20748 30714 20800
rect 45649 20791 45707 20797
rect 45649 20757 45661 20791
rect 45695 20788 45707 20791
rect 45922 20788 45928 20800
rect 45695 20760 45928 20788
rect 45695 20757 45707 20760
rect 45649 20751 45707 20757
rect 45922 20748 45928 20760
rect 45980 20748 45986 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 14182 20584 14188 20596
rect 4028 20556 14188 20584
rect 4028 20544 4034 20556
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 19242 20544 19248 20596
rect 19300 20584 19306 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 19300 20556 19717 20584
rect 19300 20544 19306 20556
rect 19705 20553 19717 20556
rect 19751 20553 19763 20587
rect 19705 20547 19763 20553
rect 22002 20544 22008 20596
rect 22060 20584 22066 20596
rect 22097 20587 22155 20593
rect 22097 20584 22109 20587
rect 22060 20556 22109 20584
rect 22060 20544 22066 20556
rect 22097 20553 22109 20556
rect 22143 20553 22155 20587
rect 22097 20547 22155 20553
rect 22278 20544 22284 20596
rect 22336 20584 22342 20596
rect 22373 20587 22431 20593
rect 22373 20584 22385 20587
rect 22336 20556 22385 20584
rect 22336 20544 22342 20556
rect 22373 20553 22385 20556
rect 22419 20553 22431 20587
rect 22373 20547 22431 20553
rect 22925 20587 22983 20593
rect 22925 20553 22937 20587
rect 22971 20584 22983 20587
rect 23474 20584 23480 20596
rect 22971 20556 23480 20584
rect 22971 20553 22983 20556
rect 22925 20547 22983 20553
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 32858 20584 32864 20596
rect 32232 20556 32864 20584
rect 32232 20528 32260 20556
rect 32858 20544 32864 20556
rect 32916 20584 32922 20596
rect 33505 20587 33563 20593
rect 33505 20584 33517 20587
rect 32916 20556 33517 20584
rect 32916 20544 32922 20556
rect 33505 20553 33517 20556
rect 33551 20553 33563 20587
rect 33505 20547 33563 20553
rect 44361 20587 44419 20593
rect 44361 20553 44373 20587
rect 44407 20584 44419 20587
rect 45738 20584 45744 20596
rect 44407 20556 45744 20584
rect 44407 20553 44419 20556
rect 44361 20547 44419 20553
rect 45738 20544 45744 20556
rect 45796 20544 45802 20596
rect 47670 20584 47676 20596
rect 47631 20556 47676 20584
rect 47670 20544 47676 20556
rect 47728 20544 47734 20596
rect 10962 20476 10968 20528
rect 11020 20516 11026 20528
rect 18233 20519 18291 20525
rect 11020 20488 12204 20516
rect 11020 20476 11026 20488
rect 11146 20408 11152 20460
rect 11204 20448 11210 20460
rect 12176 20457 12204 20488
rect 18233 20485 18245 20519
rect 18279 20516 18291 20519
rect 18506 20516 18512 20528
rect 18279 20488 18512 20516
rect 18279 20485 18291 20488
rect 18233 20479 18291 20485
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 21821 20519 21879 20525
rect 21821 20485 21833 20519
rect 21867 20516 21879 20519
rect 24118 20516 24124 20528
rect 21867 20488 24124 20516
rect 21867 20485 21879 20488
rect 21821 20479 21879 20485
rect 24118 20476 24124 20488
rect 24176 20476 24182 20528
rect 32214 20516 32220 20528
rect 32127 20488 32220 20516
rect 32214 20476 32220 20488
rect 32272 20476 32278 20528
rect 32306 20476 32312 20528
rect 32364 20516 32370 20528
rect 44082 20516 44088 20528
rect 32364 20488 32409 20516
rect 40052 20488 44088 20516
rect 32364 20476 32370 20488
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 11204 20420 11713 20448
rect 11204 20408 11210 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11977 20451 12035 20457
rect 11977 20417 11989 20451
rect 12023 20417 12035 20451
rect 11977 20411 12035 20417
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20448 12219 20451
rect 12710 20448 12716 20460
rect 12207 20420 12716 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 11992 20380 12020 20411
rect 12710 20408 12716 20420
rect 12768 20408 12774 20460
rect 12802 20408 12808 20460
rect 12860 20448 12866 20460
rect 12860 20420 12905 20448
rect 12860 20408 12866 20420
rect 14918 20408 14924 20460
rect 14976 20408 14982 20460
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 17221 20451 17279 20457
rect 17221 20448 17233 20451
rect 15160 20420 17233 20448
rect 15160 20408 15166 20420
rect 17221 20417 17233 20420
rect 17267 20417 17279 20451
rect 17954 20448 17960 20460
rect 17915 20420 17960 20448
rect 17221 20411 17279 20417
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 19334 20408 19340 20460
rect 19392 20408 19398 20460
rect 20990 20448 20996 20460
rect 20951 20420 20996 20448
rect 20990 20408 20996 20420
rect 21048 20408 21054 20460
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21968 20420 22017 20448
rect 21968 20408 21974 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22189 20451 22247 20457
rect 22189 20448 22201 20451
rect 22005 20411 22063 20417
rect 22112 20420 22201 20448
rect 12986 20380 12992 20392
rect 11992 20352 12992 20380
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 13081 20383 13139 20389
rect 13081 20349 13093 20383
rect 13127 20380 13139 20383
rect 13541 20383 13599 20389
rect 13541 20380 13553 20383
rect 13127 20352 13553 20380
rect 13127 20349 13139 20352
rect 13081 20343 13139 20349
rect 13541 20349 13553 20352
rect 13587 20349 13599 20383
rect 13541 20343 13599 20349
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20380 13875 20383
rect 15654 20380 15660 20392
rect 13863 20352 15660 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 22112 20380 22140 20420
rect 22189 20417 22201 20420
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 22833 20451 22891 20457
rect 22833 20417 22845 20451
rect 22879 20417 22891 20451
rect 24673 20451 24731 20457
rect 24673 20448 24685 20451
rect 22833 20411 22891 20417
rect 22940 20420 24685 20448
rect 22848 20380 22876 20411
rect 20220 20352 22140 20380
rect 22204 20352 22876 20380
rect 20220 20340 20226 20352
rect 22204 20324 22232 20352
rect 19242 20272 19248 20324
rect 19300 20312 19306 20324
rect 22186 20312 22192 20324
rect 19300 20284 22192 20312
rect 19300 20272 19306 20284
rect 22186 20272 22192 20284
rect 22244 20272 22250 20324
rect 22738 20272 22744 20324
rect 22796 20312 22802 20324
rect 22940 20312 22968 20420
rect 24673 20417 24685 20420
rect 24719 20448 24731 20451
rect 25406 20448 25412 20460
rect 24719 20420 25412 20448
rect 24719 20417 24731 20420
rect 24673 20411 24731 20417
rect 25406 20408 25412 20420
rect 25464 20408 25470 20460
rect 26237 20451 26295 20457
rect 26237 20417 26249 20451
rect 26283 20448 26295 20451
rect 26973 20451 27031 20457
rect 26973 20448 26985 20451
rect 26283 20420 26985 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 26973 20417 26985 20420
rect 27019 20448 27031 20451
rect 27430 20448 27436 20460
rect 27019 20420 27436 20448
rect 27019 20417 27031 20420
rect 26973 20411 27031 20417
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 30006 20408 30012 20460
rect 30064 20448 30070 20460
rect 40052 20457 40080 20488
rect 44082 20476 44088 20488
rect 44140 20476 44146 20528
rect 44634 20476 44640 20528
rect 44692 20516 44698 20528
rect 45373 20519 45431 20525
rect 45373 20516 45385 20519
rect 44692 20488 45385 20516
rect 44692 20476 44698 20488
rect 45373 20485 45385 20488
rect 45419 20485 45431 20519
rect 45373 20479 45431 20485
rect 31113 20451 31171 20457
rect 31113 20448 31125 20451
rect 30064 20420 31125 20448
rect 30064 20408 30070 20420
rect 31113 20417 31125 20420
rect 31159 20417 31171 20451
rect 31113 20411 31171 20417
rect 40037 20451 40095 20457
rect 40037 20417 40049 20451
rect 40083 20417 40095 20451
rect 40037 20411 40095 20417
rect 42613 20451 42671 20457
rect 42613 20417 42625 20451
rect 42659 20417 42671 20451
rect 42794 20448 42800 20460
rect 42755 20420 42800 20448
rect 42613 20411 42671 20417
rect 28353 20383 28411 20389
rect 28353 20349 28365 20383
rect 28399 20349 28411 20383
rect 28534 20380 28540 20392
rect 28495 20352 28540 20380
rect 28353 20343 28411 20349
rect 22796 20284 22968 20312
rect 28368 20312 28396 20343
rect 28534 20340 28540 20352
rect 28592 20340 28598 20392
rect 28810 20380 28816 20392
rect 28771 20352 28816 20380
rect 28810 20340 28816 20352
rect 28868 20340 28874 20392
rect 31128 20380 31156 20411
rect 32306 20380 32312 20392
rect 31128 20352 32312 20380
rect 32306 20340 32312 20352
rect 32364 20340 32370 20392
rect 32582 20380 32588 20392
rect 32543 20352 32588 20380
rect 32582 20340 32588 20352
rect 32640 20340 32646 20392
rect 40221 20383 40279 20389
rect 40221 20349 40233 20383
rect 40267 20380 40279 20383
rect 40402 20380 40408 20392
rect 40267 20352 40408 20380
rect 40267 20349 40279 20352
rect 40221 20343 40279 20349
rect 40402 20340 40408 20352
rect 40460 20340 40466 20392
rect 41874 20380 41880 20392
rect 41835 20352 41880 20380
rect 41874 20340 41880 20352
rect 41932 20340 41938 20392
rect 42628 20380 42656 20411
rect 42794 20408 42800 20420
rect 42852 20408 42858 20460
rect 43714 20448 43720 20460
rect 43675 20420 43720 20448
rect 43714 20408 43720 20420
rect 43772 20408 43778 20460
rect 44100 20448 44128 20476
rect 45189 20451 45247 20457
rect 45189 20448 45201 20451
rect 44100 20420 45201 20448
rect 45189 20417 45201 20420
rect 45235 20417 45247 20451
rect 45189 20411 45247 20417
rect 46750 20408 46756 20460
rect 46808 20448 46814 20460
rect 47581 20451 47639 20457
rect 47581 20448 47593 20451
rect 46808 20420 47593 20448
rect 46808 20408 46814 20420
rect 47581 20417 47593 20420
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 43070 20380 43076 20392
rect 42628 20352 43076 20380
rect 43070 20340 43076 20352
rect 43128 20340 43134 20392
rect 43806 20380 43812 20392
rect 43767 20352 43812 20380
rect 43806 20340 43812 20352
rect 43864 20340 43870 20392
rect 45830 20380 45836 20392
rect 45791 20352 45836 20380
rect 45830 20340 45836 20352
rect 45888 20380 45894 20392
rect 46934 20380 46940 20392
rect 45888 20352 46940 20380
rect 45888 20340 45894 20352
rect 46934 20340 46940 20352
rect 46992 20340 46998 20392
rect 28718 20312 28724 20324
rect 28368 20284 28724 20312
rect 22796 20272 22802 20284
rect 28718 20272 28724 20284
rect 28776 20272 28782 20324
rect 32600 20312 32628 20340
rect 28828 20284 32628 20312
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11480 20216 11529 20244
rect 11480 20204 11486 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 15102 20204 15108 20256
rect 15160 20244 15166 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 15160 20216 15301 20244
rect 15160 20204 15166 20216
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 15289 20207 15347 20213
rect 17405 20247 17463 20253
rect 17405 20213 17417 20247
rect 17451 20244 17463 20247
rect 18230 20244 18236 20256
rect 17451 20216 18236 20244
rect 17451 20213 17463 20216
rect 17405 20207 17463 20213
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 21082 20244 21088 20256
rect 21043 20216 21088 20244
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 23014 20244 23020 20256
rect 21968 20216 23020 20244
rect 21968 20204 21974 20216
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 24857 20247 24915 20253
rect 24857 20213 24869 20247
rect 24903 20244 24915 20247
rect 25038 20244 25044 20256
rect 24903 20216 25044 20244
rect 24903 20213 24915 20216
rect 24857 20207 24915 20213
rect 25038 20204 25044 20216
rect 25096 20204 25102 20256
rect 26326 20244 26332 20256
rect 26287 20216 26332 20244
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 27062 20244 27068 20256
rect 27023 20216 27068 20244
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 28166 20204 28172 20256
rect 28224 20244 28230 20256
rect 28828 20244 28856 20284
rect 40678 20272 40684 20324
rect 40736 20312 40742 20324
rect 46290 20312 46296 20324
rect 40736 20284 46296 20312
rect 40736 20272 40742 20284
rect 46290 20272 46296 20284
rect 46348 20272 46354 20324
rect 31294 20244 31300 20256
rect 28224 20216 28856 20244
rect 31255 20216 31300 20244
rect 28224 20204 28230 20216
rect 31294 20204 31300 20216
rect 31352 20204 31358 20256
rect 31573 20247 31631 20253
rect 31573 20213 31585 20247
rect 31619 20244 31631 20247
rect 32306 20244 32312 20256
rect 31619 20216 32312 20244
rect 31619 20213 31631 20216
rect 31573 20207 31631 20213
rect 32306 20204 32312 20216
rect 32364 20204 32370 20256
rect 42610 20244 42616 20256
rect 42571 20216 42616 20244
rect 42610 20204 42616 20216
rect 42668 20204 42674 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 3418 20000 3424 20052
rect 3476 20040 3482 20052
rect 28810 20040 28816 20052
rect 3476 20012 28816 20040
rect 3476 20000 3482 20012
rect 28810 20000 28816 20012
rect 28868 20000 28874 20052
rect 40402 20040 40408 20052
rect 40363 20012 40408 20040
rect 40402 20000 40408 20012
rect 40460 20000 40466 20052
rect 42150 20000 42156 20052
rect 42208 20040 42214 20052
rect 42208 20012 43668 20040
rect 42208 20000 42214 20012
rect 12710 19932 12716 19984
rect 12768 19972 12774 19984
rect 12897 19975 12955 19981
rect 12897 19972 12909 19975
rect 12768 19944 12909 19972
rect 12768 19932 12774 19944
rect 12897 19941 12909 19944
rect 12943 19972 12955 19975
rect 14093 19975 14151 19981
rect 14093 19972 14105 19975
rect 12943 19944 14105 19972
rect 12943 19941 12955 19944
rect 12897 19935 12955 19941
rect 14093 19941 14105 19944
rect 14139 19941 14151 19975
rect 14093 19935 14151 19941
rect 14366 19932 14372 19984
rect 14424 19972 14430 19984
rect 14645 19975 14703 19981
rect 14645 19972 14657 19975
rect 14424 19944 14657 19972
rect 14424 19932 14430 19944
rect 14645 19941 14657 19944
rect 14691 19941 14703 19975
rect 15654 19972 15660 19984
rect 15615 19944 15660 19972
rect 14645 19935 14703 19941
rect 15654 19932 15660 19944
rect 15712 19932 15718 19984
rect 20625 19975 20683 19981
rect 20625 19941 20637 19975
rect 20671 19972 20683 19975
rect 22833 19975 22891 19981
rect 20671 19944 21220 19972
rect 20671 19941 20683 19944
rect 20625 19935 20683 19941
rect 11422 19904 11428 19916
rect 11383 19876 11428 19904
rect 11422 19864 11428 19876
rect 11480 19864 11486 19916
rect 14826 19904 14832 19916
rect 13372 19876 14832 19904
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 13372 19845 13400 19876
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15197 19907 15255 19913
rect 15197 19904 15209 19907
rect 15068 19876 15209 19904
rect 15068 19864 15074 19876
rect 15197 19873 15209 19876
rect 15243 19873 15255 19907
rect 15197 19867 15255 19873
rect 20349 19907 20407 19913
rect 20349 19873 20361 19907
rect 20395 19873 20407 19907
rect 21082 19904 21088 19916
rect 21043 19876 21088 19904
rect 20349 19867 20407 19873
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19836 10747 19839
rect 11149 19839 11207 19845
rect 11149 19836 11161 19839
rect 10735 19808 11161 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 11149 19805 11161 19808
rect 11195 19805 11207 19839
rect 11149 19799 11207 19805
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19805 13415 19839
rect 14274 19836 14280 19848
rect 14235 19808 14280 19836
rect 13357 19799 13415 19805
rect 10612 19700 10640 19799
rect 14274 19796 14280 19808
rect 14332 19836 14338 19848
rect 15102 19836 15108 19848
rect 14332 19808 15108 19836
rect 14332 19796 14338 19808
rect 15102 19796 15108 19808
rect 15160 19836 15166 19848
rect 15289 19839 15347 19845
rect 15289 19836 15301 19839
rect 15160 19808 15301 19836
rect 15160 19796 15166 19808
rect 15289 19805 15301 19808
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 16666 19796 16672 19848
rect 16724 19836 16730 19848
rect 16945 19839 17003 19845
rect 16945 19836 16957 19839
rect 16724 19808 16957 19836
rect 16724 19796 16730 19808
rect 16945 19805 16957 19808
rect 16991 19805 17003 19839
rect 18230 19836 18236 19848
rect 18143 19808 18236 19836
rect 16945 19799 17003 19805
rect 18230 19796 18236 19808
rect 18288 19836 18294 19848
rect 19150 19836 19156 19848
rect 18288 19808 19156 19836
rect 18288 19796 18294 19808
rect 19150 19796 19156 19808
rect 19208 19796 19214 19848
rect 20257 19839 20315 19845
rect 20257 19805 20269 19839
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 13449 19771 13507 19777
rect 13449 19768 13461 19771
rect 12650 19740 13461 19768
rect 13449 19737 13461 19740
rect 13495 19737 13507 19771
rect 13449 19731 13507 19737
rect 14182 19728 14188 19780
rect 14240 19768 14246 19780
rect 14240 19740 14504 19768
rect 14240 19728 14246 19740
rect 12802 19700 12808 19712
rect 10612 19672 12808 19700
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 14366 19700 14372 19712
rect 14327 19672 14372 19700
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 14476 19709 14504 19740
rect 14461 19703 14519 19709
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 14642 19700 14648 19712
rect 14507 19672 14648 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 17037 19703 17095 19709
rect 17037 19669 17049 19703
rect 17083 19700 17095 19703
rect 17218 19700 17224 19712
rect 17083 19672 17224 19700
rect 17083 19669 17095 19672
rect 17037 19663 17095 19669
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 18230 19660 18236 19712
rect 18288 19700 18294 19712
rect 18325 19703 18383 19709
rect 18325 19700 18337 19703
rect 18288 19672 18337 19700
rect 18288 19660 18294 19672
rect 18325 19669 18337 19672
rect 18371 19669 18383 19703
rect 20272 19700 20300 19799
rect 20364 19768 20392 19867
rect 21082 19864 21088 19876
rect 21140 19864 21146 19916
rect 21192 19904 21220 19944
rect 22833 19941 22845 19975
rect 22879 19972 22891 19975
rect 24118 19972 24124 19984
rect 22879 19944 24124 19972
rect 22879 19941 22891 19944
rect 22833 19935 22891 19941
rect 21361 19907 21419 19913
rect 21361 19904 21373 19907
rect 21192 19876 21373 19904
rect 21361 19873 21373 19876
rect 21407 19873 21419 19907
rect 21361 19867 21419 19873
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 22738 19904 22744 19916
rect 21508 19876 22744 19904
rect 21508 19864 21514 19876
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 21082 19768 21088 19780
rect 20364 19740 21088 19768
rect 21082 19728 21088 19740
rect 21140 19728 21146 19780
rect 22370 19728 22376 19780
rect 22428 19728 22434 19780
rect 22848 19700 22876 19935
rect 24118 19932 24124 19944
rect 24176 19932 24182 19984
rect 43438 19972 43444 19984
rect 28828 19944 35894 19972
rect 43399 19944 43444 19972
rect 28828 19916 28856 19944
rect 25038 19904 25044 19916
rect 24999 19876 25044 19904
rect 25038 19864 25044 19876
rect 25096 19864 25102 19916
rect 26878 19864 26884 19916
rect 26936 19904 26942 19916
rect 27065 19907 27123 19913
rect 27065 19904 27077 19907
rect 26936 19876 27077 19904
rect 26936 19864 26942 19876
rect 27065 19873 27077 19876
rect 27111 19904 27123 19907
rect 27154 19904 27160 19916
rect 27111 19876 27160 19904
rect 27111 19873 27123 19876
rect 27065 19867 27123 19873
rect 27154 19864 27160 19876
rect 27212 19864 27218 19916
rect 28169 19907 28227 19913
rect 28169 19873 28181 19907
rect 28215 19904 28227 19907
rect 28258 19904 28264 19916
rect 28215 19876 28264 19904
rect 28215 19873 28227 19876
rect 28169 19867 28227 19873
rect 28258 19864 28264 19876
rect 28316 19864 28322 19916
rect 28810 19864 28816 19916
rect 28868 19864 28874 19916
rect 30650 19904 30656 19916
rect 30611 19876 30656 19904
rect 30650 19864 30656 19876
rect 30708 19864 30714 19916
rect 32309 19907 32367 19913
rect 32309 19873 32321 19907
rect 32355 19904 32367 19907
rect 33042 19904 33048 19916
rect 32355 19876 33048 19904
rect 32355 19873 32367 19876
rect 32309 19867 32367 19873
rect 33042 19864 33048 19876
rect 33100 19864 33106 19916
rect 35866 19904 35894 19944
rect 43438 19932 43444 19944
rect 43496 19932 43502 19984
rect 43640 19972 43668 20012
rect 43714 20000 43720 20052
rect 43772 20040 43778 20052
rect 43993 20043 44051 20049
rect 43993 20040 44005 20043
rect 43772 20012 44005 20040
rect 43772 20000 43778 20012
rect 43993 20009 44005 20012
rect 44039 20009 44051 20043
rect 43993 20003 44051 20009
rect 45830 19972 45836 19984
rect 43640 19944 45836 19972
rect 45830 19932 45836 19944
rect 45888 19972 45894 19984
rect 45888 19944 46244 19972
rect 45888 19932 45894 19944
rect 40678 19904 40684 19916
rect 35866 19876 40684 19904
rect 40678 19864 40684 19876
rect 40736 19864 40742 19916
rect 42610 19864 42616 19916
rect 42668 19904 42674 19916
rect 45738 19904 45744 19916
rect 42668 19876 44220 19904
rect 45699 19876 45744 19904
rect 42668 19864 42674 19876
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19836 24639 19839
rect 24854 19836 24860 19848
rect 24627 19808 24860 19836
rect 24627 19805 24639 19808
rect 24581 19799 24639 19805
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 28350 19836 28356 19848
rect 28311 19808 28356 19836
rect 28350 19796 28356 19808
rect 28408 19796 28414 19848
rect 30469 19839 30527 19845
rect 30469 19805 30481 19839
rect 30515 19805 30527 19839
rect 30469 19799 30527 19805
rect 40313 19839 40371 19845
rect 40313 19805 40325 19839
rect 40359 19805 40371 19839
rect 40313 19799 40371 19805
rect 25317 19771 25375 19777
rect 25317 19737 25329 19771
rect 25363 19737 25375 19771
rect 25317 19731 25375 19737
rect 20272 19672 22876 19700
rect 24397 19703 24455 19709
rect 18325 19663 18383 19669
rect 24397 19669 24409 19703
rect 24443 19700 24455 19703
rect 25332 19700 25360 19731
rect 26326 19728 26332 19780
rect 26384 19728 26390 19780
rect 27154 19728 27160 19780
rect 27212 19768 27218 19780
rect 30484 19768 30512 19799
rect 27212 19740 30512 19768
rect 27212 19728 27218 19740
rect 24443 19672 25360 19700
rect 28537 19703 28595 19709
rect 24443 19669 24455 19672
rect 24397 19663 24455 19669
rect 28537 19669 28549 19703
rect 28583 19700 28595 19703
rect 28902 19700 28908 19712
rect 28583 19672 28908 19700
rect 28583 19669 28595 19672
rect 28537 19663 28595 19669
rect 28902 19660 28908 19672
rect 28960 19660 28966 19712
rect 40328 19700 40356 19799
rect 42242 19796 42248 19848
rect 42300 19836 42306 19848
rect 42797 19839 42855 19845
rect 42797 19836 42809 19839
rect 42300 19808 42809 19836
rect 42300 19796 42306 19808
rect 42797 19805 42809 19808
rect 42843 19805 42855 19839
rect 42797 19799 42855 19805
rect 42981 19839 43039 19845
rect 42981 19805 42993 19839
rect 43027 19805 43039 19839
rect 43254 19836 43260 19848
rect 43215 19808 43260 19836
rect 42981 19799 43039 19805
rect 42996 19768 43024 19799
rect 43254 19796 43260 19808
rect 43312 19796 43318 19848
rect 43438 19836 43444 19848
rect 43399 19808 43444 19836
rect 43438 19796 43444 19808
rect 43496 19836 43502 19848
rect 44192 19845 44220 19876
rect 45738 19864 45744 19876
rect 45796 19864 45802 19916
rect 45922 19904 45928 19916
rect 45883 19876 45928 19904
rect 45922 19864 45928 19876
rect 45980 19864 45986 19916
rect 46216 19913 46244 19944
rect 46201 19907 46259 19913
rect 46201 19873 46213 19907
rect 46247 19873 46259 19907
rect 46201 19867 46259 19873
rect 43993 19839 44051 19845
rect 43993 19836 44005 19839
rect 43496 19808 44005 19836
rect 43496 19796 43502 19808
rect 43993 19805 44005 19808
rect 44039 19805 44051 19839
rect 43993 19799 44051 19805
rect 44177 19839 44235 19845
rect 44177 19805 44189 19839
rect 44223 19805 44235 19839
rect 44177 19799 44235 19805
rect 45281 19839 45339 19845
rect 45281 19805 45293 19839
rect 45327 19836 45339 19839
rect 45554 19836 45560 19848
rect 45327 19808 45560 19836
rect 45327 19805 45339 19808
rect 45281 19799 45339 19805
rect 45554 19796 45560 19808
rect 45612 19796 45618 19848
rect 43714 19768 43720 19780
rect 42996 19740 43720 19768
rect 43714 19728 43720 19740
rect 43772 19728 43778 19780
rect 46474 19768 46480 19780
rect 43916 19740 46480 19768
rect 41138 19700 41144 19712
rect 40328 19672 41144 19700
rect 41138 19660 41144 19672
rect 41196 19700 41202 19712
rect 43916 19700 43944 19740
rect 46474 19728 46480 19740
rect 46532 19728 46538 19780
rect 41196 19672 43944 19700
rect 41196 19660 41202 19672
rect 45002 19660 45008 19712
rect 45060 19700 45066 19712
rect 45097 19703 45155 19709
rect 45097 19700 45109 19703
rect 45060 19672 45109 19700
rect 45060 19660 45066 19672
rect 45097 19669 45109 19672
rect 45143 19669 45155 19703
rect 45097 19663 45155 19669
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 13906 19456 13912 19508
rect 13964 19496 13970 19508
rect 15010 19496 15016 19508
rect 13964 19468 15016 19496
rect 13964 19456 13970 19468
rect 15010 19456 15016 19468
rect 15068 19496 15074 19508
rect 15289 19499 15347 19505
rect 15289 19496 15301 19499
rect 15068 19468 15301 19496
rect 15068 19456 15074 19468
rect 15289 19465 15301 19468
rect 15335 19465 15347 19499
rect 15289 19459 15347 19465
rect 20162 19456 20168 19508
rect 20220 19496 20226 19508
rect 20993 19499 21051 19505
rect 20220 19468 20852 19496
rect 20220 19456 20226 19468
rect 14093 19431 14151 19437
rect 14093 19397 14105 19431
rect 14139 19428 14151 19431
rect 14366 19428 14372 19440
rect 14139 19400 14372 19428
rect 14139 19397 14151 19400
rect 14093 19391 14151 19397
rect 14366 19388 14372 19400
rect 14424 19428 14430 19440
rect 14734 19428 14740 19440
rect 14424 19400 14740 19428
rect 14424 19388 14430 19400
rect 14734 19388 14740 19400
rect 14792 19428 14798 19440
rect 14921 19431 14979 19437
rect 14921 19428 14933 19431
rect 14792 19400 14933 19428
rect 14792 19388 14798 19400
rect 14921 19397 14933 19400
rect 14967 19397 14979 19431
rect 15121 19431 15179 19437
rect 15121 19428 15133 19431
rect 14921 19391 14979 19397
rect 15028 19400 15133 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 12802 19320 12808 19372
rect 12860 19360 12866 19372
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 12860 19332 13093 19360
rect 12860 19320 12866 19332
rect 13081 19329 13093 19332
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19360 13231 19363
rect 13998 19360 14004 19372
rect 13219 19332 14004 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 14182 19360 14188 19372
rect 14143 19332 14188 19360
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 14550 19360 14556 19372
rect 14323 19332 14556 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 14550 19320 14556 19332
rect 14608 19360 14614 19372
rect 15028 19360 15056 19400
rect 15121 19397 15133 19400
rect 15167 19397 15179 19431
rect 15121 19391 15179 19397
rect 18230 19388 18236 19440
rect 18288 19388 18294 19440
rect 20824 19437 20852 19468
rect 20993 19465 21005 19499
rect 21039 19496 21051 19499
rect 21082 19496 21088 19508
rect 21039 19468 21088 19496
rect 21039 19465 21051 19468
rect 20993 19459 21051 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 22281 19499 22339 19505
rect 22281 19465 22293 19499
rect 22327 19496 22339 19499
rect 22370 19496 22376 19508
rect 22327 19468 22376 19496
rect 22327 19465 22339 19468
rect 22281 19459 22339 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 28350 19496 28356 19508
rect 23124 19468 28212 19496
rect 28311 19468 28356 19496
rect 19889 19431 19947 19437
rect 19889 19397 19901 19431
rect 19935 19428 19947 19431
rect 20625 19431 20683 19437
rect 20625 19428 20637 19431
rect 19935 19400 20637 19428
rect 19935 19397 19947 19400
rect 19889 19391 19947 19397
rect 20625 19397 20637 19400
rect 20671 19397 20683 19431
rect 20824 19431 20883 19437
rect 20824 19400 20837 19431
rect 20625 19391 20683 19397
rect 20825 19397 20837 19400
rect 20871 19397 20883 19431
rect 23014 19428 23020 19440
rect 20825 19391 20883 19397
rect 22066 19400 23020 19428
rect 17218 19360 17224 19372
rect 14608 19332 15056 19360
rect 17179 19332 17224 19360
rect 14608 19320 14614 19332
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 20073 19363 20131 19369
rect 20073 19360 20085 19363
rect 18984 19332 20085 19360
rect 18984 19304 19012 19332
rect 20073 19329 20085 19332
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 17497 19295 17555 19301
rect 2746 19264 17264 19292
rect 1578 19184 1584 19236
rect 1636 19224 1642 19236
rect 2746 19224 2774 19264
rect 1636 19196 2774 19224
rect 13909 19227 13967 19233
rect 1636 19184 1642 19196
rect 13909 19193 13921 19227
rect 13955 19224 13967 19227
rect 14274 19224 14280 19236
rect 13955 19196 14280 19224
rect 13955 19193 13967 19196
rect 13909 19187 13967 19193
rect 14274 19184 14280 19196
rect 14332 19184 14338 19236
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 14461 19159 14519 19165
rect 14461 19156 14473 19159
rect 13044 19128 14473 19156
rect 13044 19116 13050 19128
rect 14461 19125 14473 19128
rect 14507 19125 14519 19159
rect 14461 19119 14519 19125
rect 14642 19116 14648 19168
rect 14700 19156 14706 19168
rect 15105 19159 15163 19165
rect 15105 19156 15117 19159
rect 14700 19128 15117 19156
rect 14700 19116 14706 19128
rect 15105 19125 15117 19128
rect 15151 19125 15163 19159
rect 17236 19156 17264 19264
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 18506 19292 18512 19304
rect 17543 19264 18512 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 18966 19292 18972 19304
rect 18879 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 20088 19292 20116 19323
rect 20162 19320 20168 19372
rect 20220 19360 20226 19372
rect 20640 19360 20668 19391
rect 22066 19360 22094 19400
rect 23014 19388 23020 19400
rect 23072 19388 23078 19440
rect 22186 19360 22192 19372
rect 20220 19332 20265 19360
rect 20640 19332 22094 19360
rect 22147 19332 22192 19360
rect 20220 19320 20226 19332
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 23124 19360 23152 19468
rect 26234 19428 26240 19440
rect 24596 19400 26240 19428
rect 24596 19369 24624 19400
rect 26234 19388 26240 19400
rect 26292 19428 26298 19440
rect 27154 19428 27160 19440
rect 26292 19400 27160 19428
rect 26292 19388 26298 19400
rect 27154 19388 27160 19400
rect 27212 19388 27218 19440
rect 27982 19428 27988 19440
rect 27943 19400 27988 19428
rect 27982 19388 27988 19400
rect 28040 19388 28046 19440
rect 28184 19428 28212 19468
rect 28350 19456 28356 19468
rect 28408 19456 28414 19508
rect 28534 19456 28540 19508
rect 28592 19496 28598 19508
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 28592 19468 28917 19496
rect 28592 19456 28598 19468
rect 28905 19465 28917 19468
rect 28951 19465 28963 19499
rect 28905 19459 28963 19465
rect 31754 19456 31760 19508
rect 31812 19496 31818 19508
rect 32125 19499 32183 19505
rect 32125 19496 32137 19499
rect 31812 19468 32137 19496
rect 31812 19456 31818 19468
rect 32125 19465 32137 19468
rect 32171 19465 32183 19499
rect 32125 19459 32183 19465
rect 43257 19499 43315 19505
rect 43257 19465 43269 19499
rect 43303 19496 43315 19499
rect 43438 19496 43444 19508
rect 43303 19468 43444 19496
rect 43303 19465 43315 19468
rect 43257 19459 43315 19465
rect 43438 19456 43444 19468
rect 43496 19456 43502 19508
rect 43806 19496 43812 19508
rect 43767 19468 43812 19496
rect 43806 19456 43812 19468
rect 43864 19456 43870 19508
rect 28184 19400 28672 19428
rect 22296 19332 23152 19360
rect 24581 19363 24639 19369
rect 20806 19292 20812 19304
rect 20088 19264 20812 19292
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 22296 19292 22324 19332
rect 24581 19329 24593 19363
rect 24627 19329 24639 19363
rect 25406 19360 25412 19372
rect 25367 19332 25412 19360
rect 24581 19323 24639 19329
rect 25406 19320 25412 19332
rect 25464 19320 25470 19372
rect 28166 19360 28172 19372
rect 28127 19332 28172 19360
rect 28166 19320 28172 19332
rect 28224 19320 28230 19372
rect 24670 19292 24676 19304
rect 20956 19264 22324 19292
rect 24631 19264 24676 19292
rect 20956 19252 20962 19264
rect 24670 19252 24676 19264
rect 24728 19252 24734 19304
rect 28644 19292 28672 19400
rect 28718 19388 28724 19440
rect 28776 19428 28782 19440
rect 29733 19431 29791 19437
rect 28776 19400 29592 19428
rect 28776 19388 28782 19400
rect 28810 19360 28816 19372
rect 28771 19332 28816 19360
rect 28810 19320 28816 19332
rect 28868 19320 28874 19372
rect 29564 19369 29592 19400
rect 29733 19397 29745 19431
rect 29779 19428 29791 19431
rect 30374 19428 30380 19440
rect 29779 19400 30380 19428
rect 29779 19397 29791 19400
rect 29733 19391 29791 19397
rect 30374 19388 30380 19400
rect 30432 19388 30438 19440
rect 41414 19428 41420 19440
rect 31220 19400 41420 19428
rect 29549 19363 29607 19369
rect 28920 19332 29500 19360
rect 28920 19292 28948 19332
rect 24780 19264 26234 19292
rect 28644 19264 28948 19292
rect 29472 19292 29500 19332
rect 29549 19329 29561 19363
rect 29595 19329 29607 19363
rect 29549 19323 29607 19329
rect 30009 19295 30067 19301
rect 30009 19292 30021 19295
rect 29472 19264 30021 19292
rect 24780 19224 24808 19264
rect 18524 19196 24808 19224
rect 24949 19227 25007 19233
rect 18524 19156 18552 19196
rect 24949 19193 24961 19227
rect 24995 19224 25007 19227
rect 25498 19224 25504 19236
rect 24995 19196 25504 19224
rect 24995 19193 25007 19196
rect 24949 19187 25007 19193
rect 25498 19184 25504 19196
rect 25556 19184 25562 19236
rect 26206 19224 26234 19264
rect 30009 19261 30021 19264
rect 30055 19292 30067 19295
rect 30466 19292 30472 19304
rect 30055 19264 30472 19292
rect 30055 19261 30067 19264
rect 30009 19255 30067 19261
rect 30466 19252 30472 19264
rect 30524 19292 30530 19304
rect 31220 19292 31248 19400
rect 41414 19388 41420 19400
rect 41472 19428 41478 19440
rect 42150 19428 42156 19440
rect 41472 19400 42156 19428
rect 41472 19388 41478 19400
rect 42150 19388 42156 19400
rect 42208 19388 42214 19440
rect 42242 19388 42248 19440
rect 42300 19428 42306 19440
rect 42300 19400 43760 19428
rect 42300 19388 42306 19400
rect 32306 19360 32312 19372
rect 32267 19332 32312 19360
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 42794 19320 42800 19372
rect 42852 19360 42858 19372
rect 42889 19363 42947 19369
rect 42889 19360 42901 19363
rect 42852 19332 42901 19360
rect 42852 19320 42858 19332
rect 42889 19329 42901 19332
rect 42935 19329 42947 19363
rect 43070 19360 43076 19372
rect 43031 19332 43076 19360
rect 42889 19323 42947 19329
rect 43070 19320 43076 19332
rect 43128 19320 43134 19372
rect 43732 19369 43760 19400
rect 44174 19388 44180 19440
rect 44232 19428 44238 19440
rect 47765 19431 47823 19437
rect 47765 19428 47777 19431
rect 44232 19400 47777 19428
rect 44232 19388 44238 19400
rect 47765 19397 47777 19400
rect 47811 19397 47823 19431
rect 47765 19391 47823 19397
rect 43717 19363 43775 19369
rect 43717 19329 43729 19363
rect 43763 19329 43775 19363
rect 43898 19360 43904 19372
rect 43859 19332 43904 19360
rect 43717 19323 43775 19329
rect 43898 19320 43904 19332
rect 43956 19320 43962 19372
rect 44082 19320 44088 19372
rect 44140 19360 44146 19372
rect 45189 19363 45247 19369
rect 45189 19360 45201 19363
rect 44140 19332 45201 19360
rect 44140 19320 44146 19332
rect 45189 19329 45201 19332
rect 45235 19329 45247 19363
rect 45189 19323 45247 19329
rect 47857 19363 47915 19369
rect 47857 19329 47869 19363
rect 47903 19329 47915 19363
rect 47857 19323 47915 19329
rect 43162 19292 43168 19304
rect 30524 19264 31248 19292
rect 31496 19264 43168 19292
rect 30524 19252 30530 19264
rect 31496 19224 31524 19264
rect 43162 19252 43168 19264
rect 43220 19252 43226 19304
rect 43254 19252 43260 19304
rect 43312 19292 43318 19304
rect 43916 19292 43944 19320
rect 45370 19292 45376 19304
rect 43312 19264 43944 19292
rect 45331 19264 45376 19292
rect 43312 19252 43318 19264
rect 45370 19252 45376 19264
rect 45428 19252 45434 19304
rect 45830 19292 45836 19304
rect 45791 19264 45836 19292
rect 45830 19252 45836 19264
rect 45888 19252 45894 19304
rect 46842 19224 46848 19236
rect 26206 19196 31524 19224
rect 35866 19196 46848 19224
rect 17236 19128 18552 19156
rect 19889 19159 19947 19165
rect 15105 19119 15163 19125
rect 19889 19125 19901 19159
rect 19935 19156 19947 19159
rect 20530 19156 20536 19168
rect 19935 19128 20536 19156
rect 19935 19125 19947 19128
rect 19889 19119 19947 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 20806 19156 20812 19168
rect 20719 19128 20812 19156
rect 20806 19116 20812 19128
rect 20864 19156 20870 19168
rect 22002 19156 22008 19168
rect 20864 19128 22008 19156
rect 20864 19116 20870 19128
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 25222 19116 25228 19168
rect 25280 19156 25286 19168
rect 25409 19159 25467 19165
rect 25409 19156 25421 19159
rect 25280 19128 25421 19156
rect 25280 19116 25286 19128
rect 25409 19125 25421 19128
rect 25455 19125 25467 19159
rect 25409 19119 25467 19125
rect 25682 19116 25688 19168
rect 25740 19156 25746 19168
rect 35866 19156 35894 19196
rect 46842 19184 46848 19196
rect 46900 19184 46906 19236
rect 47578 19224 47584 19236
rect 47539 19196 47584 19224
rect 47578 19184 47584 19196
rect 47636 19184 47642 19236
rect 25740 19128 35894 19156
rect 25740 19116 25746 19128
rect 43162 19116 43168 19168
rect 43220 19156 43226 19168
rect 43990 19156 43996 19168
rect 43220 19128 43996 19156
rect 43220 19116 43226 19128
rect 43990 19116 43996 19128
rect 44048 19156 44054 19168
rect 47872 19156 47900 19323
rect 47946 19320 47952 19372
rect 48004 19360 48010 19372
rect 48004 19332 48049 19360
rect 48004 19320 48010 19332
rect 48038 19252 48044 19304
rect 48096 19292 48102 19304
rect 48133 19295 48191 19301
rect 48133 19292 48145 19295
rect 48096 19264 48145 19292
rect 48096 19252 48102 19264
rect 48133 19261 48145 19264
rect 48179 19261 48191 19295
rect 48133 19255 48191 19261
rect 44048 19128 47900 19156
rect 44048 19116 44054 19128
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 43901 18955 43959 18961
rect 3292 18924 35894 18952
rect 3292 18912 3298 18924
rect 18506 18884 18512 18896
rect 18467 18856 18512 18884
rect 18506 18844 18512 18856
rect 18564 18844 18570 18896
rect 20898 18844 20904 18896
rect 20956 18884 20962 18896
rect 21174 18884 21180 18896
rect 20956 18856 21180 18884
rect 20956 18844 20962 18856
rect 21174 18844 21180 18856
rect 21232 18844 21238 18896
rect 26973 18887 27031 18893
rect 26973 18853 26985 18887
rect 27019 18884 27031 18887
rect 27154 18884 27160 18896
rect 27019 18856 27160 18884
rect 27019 18853 27031 18856
rect 26973 18847 27031 18853
rect 27154 18844 27160 18856
rect 27212 18844 27218 18896
rect 28718 18884 28724 18896
rect 28679 18856 28724 18884
rect 28718 18844 28724 18856
rect 28776 18844 28782 18896
rect 13998 18776 14004 18828
rect 14056 18816 14062 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 14056 18788 14105 18816
rect 14056 18776 14062 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 18233 18819 18291 18825
rect 14976 18788 16712 18816
rect 14976 18776 14982 18788
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 2314 18748 2320 18760
rect 2179 18720 2320 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 2314 18708 2320 18720
rect 2372 18748 2378 18760
rect 13354 18748 13360 18760
rect 2372 18720 2774 18748
rect 13315 18720 13360 18748
rect 2372 18708 2378 18720
rect 2746 18612 2774 18720
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 13906 18748 13912 18760
rect 13587 18720 13912 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 13906 18708 13912 18720
rect 13964 18708 13970 18760
rect 16684 18757 16712 18788
rect 18233 18785 18245 18819
rect 18279 18816 18291 18819
rect 20162 18816 20168 18828
rect 18279 18788 20168 18816
rect 18279 18785 18291 18788
rect 18233 18779 18291 18785
rect 20162 18776 20168 18788
rect 20220 18776 20226 18828
rect 21082 18816 21088 18828
rect 20732 18788 21088 18816
rect 16669 18751 16727 18757
rect 16669 18717 16681 18751
rect 16715 18748 16727 18751
rect 16758 18748 16764 18760
rect 16715 18720 16764 18748
rect 16715 18717 16727 18720
rect 16669 18711 16727 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18748 18199 18751
rect 18966 18748 18972 18760
rect 18187 18720 18972 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 18966 18708 18972 18720
rect 19024 18708 19030 18760
rect 20530 18748 20536 18760
rect 20491 18720 20536 18748
rect 20530 18708 20536 18720
rect 20588 18708 20594 18760
rect 20732 18757 20760 18788
rect 21082 18776 21088 18788
rect 21140 18776 21146 18828
rect 25222 18816 25228 18828
rect 25183 18788 25228 18816
rect 25222 18776 25228 18788
rect 25280 18776 25286 18828
rect 25498 18816 25504 18828
rect 25459 18788 25504 18816
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 30466 18816 30472 18828
rect 30427 18788 30472 18816
rect 30466 18776 30472 18788
rect 30524 18776 30530 18828
rect 35866 18816 35894 18924
rect 43901 18921 43913 18955
rect 43947 18952 43959 18955
rect 45370 18952 45376 18964
rect 43947 18924 45376 18952
rect 43947 18921 43959 18924
rect 43901 18915 43959 18921
rect 45370 18912 45376 18924
rect 45428 18912 45434 18964
rect 47578 18912 47584 18964
rect 47636 18952 47642 18964
rect 48038 18952 48044 18964
rect 47636 18924 48044 18952
rect 47636 18912 47642 18924
rect 48038 18912 48044 18924
rect 48096 18912 48102 18964
rect 45097 18819 45155 18825
rect 45097 18816 45109 18819
rect 35866 18788 40724 18816
rect 40696 18760 40724 18788
rect 42444 18788 45109 18816
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18717 20775 18751
rect 21174 18748 21180 18760
rect 21135 18720 21180 18748
rect 20717 18711 20775 18717
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 23658 18748 23664 18760
rect 23619 18720 23664 18748
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18748 23903 18751
rect 24302 18748 24308 18760
rect 23891 18720 24308 18748
rect 23891 18717 23903 18720
rect 23845 18711 23903 18717
rect 24302 18708 24308 18720
rect 24360 18748 24366 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24360 18720 24593 18748
rect 24360 18708 24366 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 27982 18748 27988 18760
rect 27943 18720 27988 18748
rect 24581 18711 24639 18717
rect 27982 18708 27988 18720
rect 28040 18708 28046 18760
rect 28166 18748 28172 18760
rect 28127 18720 28172 18748
rect 28166 18708 28172 18720
rect 28224 18708 28230 18760
rect 28902 18748 28908 18760
rect 28863 18720 28908 18748
rect 28902 18708 28908 18720
rect 28960 18708 28966 18760
rect 29638 18748 29644 18760
rect 29599 18720 29644 18748
rect 29638 18708 29644 18720
rect 29696 18708 29702 18760
rect 40494 18748 40500 18760
rect 40455 18720 40500 18748
rect 40494 18708 40500 18720
rect 40552 18708 40558 18760
rect 40678 18708 40684 18760
rect 40736 18748 40742 18760
rect 40736 18720 40829 18748
rect 40736 18708 40742 18720
rect 41690 18708 41696 18760
rect 41748 18748 41754 18760
rect 42444 18757 42472 18788
rect 45097 18785 45109 18788
rect 45143 18785 45155 18819
rect 47596 18816 47624 18912
rect 48130 18816 48136 18828
rect 45097 18779 45155 18785
rect 45388 18788 47624 18816
rect 48091 18788 48136 18816
rect 42429 18751 42487 18757
rect 42429 18748 42441 18751
rect 41748 18720 42441 18748
rect 41748 18708 41754 18720
rect 42429 18717 42441 18720
rect 42475 18717 42487 18751
rect 42429 18711 42487 18717
rect 42613 18751 42671 18757
rect 42613 18717 42625 18751
rect 42659 18748 42671 18751
rect 43254 18748 43260 18760
rect 42659 18720 43260 18748
rect 42659 18717 42671 18720
rect 42613 18711 42671 18717
rect 43254 18708 43260 18720
rect 43312 18708 43318 18760
rect 43441 18751 43499 18757
rect 43441 18717 43453 18751
rect 43487 18717 43499 18751
rect 43441 18711 43499 18717
rect 13449 18683 13507 18689
rect 13449 18649 13461 18683
rect 13495 18680 13507 18683
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 13495 18652 14381 18680
rect 13495 18649 13507 18652
rect 13449 18643 13507 18649
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 15102 18640 15108 18692
rect 15160 18640 15166 18692
rect 16022 18640 16028 18692
rect 16080 18680 16086 18692
rect 16945 18683 17003 18689
rect 16945 18680 16957 18683
rect 16080 18652 16957 18680
rect 16080 18640 16086 18652
rect 16945 18649 16957 18652
rect 16991 18649 17003 18683
rect 16945 18643 17003 18649
rect 20625 18683 20683 18689
rect 20625 18649 20637 18683
rect 20671 18680 20683 18683
rect 21453 18683 21511 18689
rect 21453 18680 21465 18683
rect 20671 18652 21465 18680
rect 20671 18649 20683 18652
rect 20625 18643 20683 18649
rect 21453 18649 21465 18652
rect 21499 18649 21511 18683
rect 21453 18643 21511 18649
rect 22094 18640 22100 18692
rect 22152 18640 22158 18692
rect 23676 18680 23704 18708
rect 24394 18680 24400 18692
rect 23676 18652 24400 18680
rect 24394 18640 24400 18652
rect 24452 18640 24458 18692
rect 27062 18680 27068 18692
rect 26726 18652 27068 18680
rect 27062 18640 27068 18652
rect 27120 18640 27126 18692
rect 28258 18680 28264 18692
rect 28219 18652 28264 18680
rect 28258 18640 28264 18652
rect 28316 18640 28322 18692
rect 29822 18680 29828 18692
rect 29783 18652 29828 18680
rect 29822 18640 29828 18652
rect 29880 18640 29886 18692
rect 13722 18612 13728 18624
rect 2746 18584 13728 18612
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 14274 18572 14280 18624
rect 14332 18612 14338 18624
rect 14734 18612 14740 18624
rect 14332 18584 14740 18612
rect 14332 18572 14338 18584
rect 14734 18572 14740 18584
rect 14792 18612 14798 18624
rect 15841 18615 15899 18621
rect 15841 18612 15853 18615
rect 14792 18584 15853 18612
rect 14792 18572 14798 18584
rect 15841 18581 15853 18584
rect 15887 18612 15899 18615
rect 16390 18612 16396 18624
rect 15887 18584 16396 18612
rect 15887 18581 15899 18584
rect 15841 18575 15899 18581
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 22925 18615 22983 18621
rect 22925 18581 22937 18615
rect 22971 18612 22983 18615
rect 23014 18612 23020 18624
rect 22971 18584 23020 18612
rect 22971 18581 22983 18584
rect 22925 18575 22983 18581
rect 23014 18572 23020 18584
rect 23072 18572 23078 18624
rect 23845 18615 23903 18621
rect 23845 18581 23857 18615
rect 23891 18612 23903 18615
rect 24670 18612 24676 18624
rect 23891 18584 24676 18612
rect 23891 18581 23903 18584
rect 23845 18575 23903 18581
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 24946 18612 24952 18624
rect 24811 18584 24952 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 40681 18615 40739 18621
rect 40681 18581 40693 18615
rect 40727 18612 40739 18615
rect 41046 18612 41052 18624
rect 40727 18584 41052 18612
rect 40727 18581 40739 18584
rect 40681 18575 40739 18581
rect 41046 18572 41052 18584
rect 41104 18572 41110 18624
rect 42613 18615 42671 18621
rect 42613 18581 42625 18615
rect 42659 18612 42671 18615
rect 42702 18612 42708 18624
rect 42659 18584 42708 18612
rect 42659 18581 42671 18584
rect 42613 18575 42671 18581
rect 42702 18572 42708 18584
rect 42760 18572 42766 18624
rect 43456 18612 43484 18711
rect 43806 18708 43812 18760
rect 43864 18748 43870 18760
rect 43990 18748 43996 18760
rect 43864 18720 43996 18748
rect 43864 18708 43870 18720
rect 43990 18708 43996 18720
rect 44048 18708 44054 18760
rect 44174 18748 44180 18760
rect 44135 18720 44180 18748
rect 44174 18708 44180 18720
rect 44232 18708 44238 18760
rect 44453 18751 44511 18757
rect 44453 18717 44465 18751
rect 44499 18717 44511 18751
rect 45002 18748 45008 18760
rect 44963 18720 45008 18748
rect 44453 18711 44511 18717
rect 43714 18640 43720 18692
rect 43772 18680 43778 18692
rect 44468 18680 44496 18711
rect 45002 18708 45008 18720
rect 45060 18708 45066 18760
rect 45189 18751 45247 18757
rect 45189 18717 45201 18751
rect 45235 18748 45247 18751
rect 45278 18748 45284 18760
rect 45235 18720 45284 18748
rect 45235 18717 45247 18720
rect 45189 18711 45247 18717
rect 45278 18708 45284 18720
rect 45336 18708 45342 18760
rect 45388 18680 45416 18788
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 45833 18751 45891 18757
rect 45833 18717 45845 18751
rect 45879 18748 45891 18751
rect 46293 18751 46351 18757
rect 46293 18748 46305 18751
rect 45879 18720 46305 18748
rect 45879 18717 45891 18720
rect 45833 18711 45891 18717
rect 46293 18717 46305 18720
rect 46339 18717 46351 18751
rect 46293 18711 46351 18717
rect 43772 18652 45416 18680
rect 46477 18683 46535 18689
rect 43772 18640 43778 18652
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 47670 18680 47676 18692
rect 46523 18652 47676 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 47670 18640 47676 18652
rect 47728 18640 47734 18692
rect 47210 18612 47216 18624
rect 43456 18584 47216 18612
rect 47210 18572 47216 18584
rect 47268 18612 47274 18624
rect 47946 18612 47952 18624
rect 47268 18584 47952 18612
rect 47268 18572 47274 18584
rect 47946 18572 47952 18584
rect 48004 18572 48010 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 29454 18408 29460 18420
rect 1627 18380 29460 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 29454 18368 29460 18380
rect 29512 18368 29518 18420
rect 29822 18368 29828 18420
rect 29880 18408 29886 18420
rect 32125 18411 32183 18417
rect 32125 18408 32137 18411
rect 29880 18380 32137 18408
rect 29880 18368 29886 18380
rect 32125 18377 32137 18380
rect 32171 18377 32183 18411
rect 44174 18408 44180 18420
rect 32125 18371 32183 18377
rect 32324 18380 44180 18408
rect 14274 18340 14280 18352
rect 14235 18312 14280 18340
rect 14274 18300 14280 18312
rect 14332 18300 14338 18352
rect 15102 18340 15108 18352
rect 15063 18312 15108 18340
rect 15102 18300 15108 18312
rect 15160 18300 15166 18352
rect 18049 18343 18107 18349
rect 18049 18309 18061 18343
rect 18095 18340 18107 18343
rect 18785 18343 18843 18349
rect 18785 18340 18797 18343
rect 18095 18312 18797 18340
rect 18095 18309 18107 18312
rect 18049 18303 18107 18309
rect 18785 18309 18797 18312
rect 18831 18309 18843 18343
rect 18785 18303 18843 18309
rect 21174 18300 21180 18352
rect 21232 18340 21238 18352
rect 21269 18343 21327 18349
rect 21269 18340 21281 18343
rect 21232 18312 21281 18340
rect 21232 18300 21238 18312
rect 21269 18309 21281 18312
rect 21315 18309 21327 18343
rect 21269 18303 21327 18309
rect 22094 18300 22100 18352
rect 22152 18340 22158 18352
rect 22281 18343 22339 18349
rect 22281 18340 22293 18343
rect 22152 18312 22293 18340
rect 22152 18300 22158 18312
rect 22281 18309 22293 18312
rect 22327 18309 22339 18343
rect 22281 18303 22339 18309
rect 24854 18300 24860 18352
rect 24912 18340 24918 18352
rect 25133 18343 25191 18349
rect 25133 18340 25145 18343
rect 24912 18312 25145 18340
rect 24912 18300 24918 18312
rect 25133 18309 25145 18312
rect 25179 18309 25191 18343
rect 25133 18303 25191 18309
rect 26206 18312 30236 18340
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 14458 18272 14464 18284
rect 14419 18244 14464 18272
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 14918 18272 14924 18284
rect 14608 18244 14924 18272
rect 14608 18232 14614 18244
rect 14918 18232 14924 18244
rect 14976 18232 14982 18284
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18272 15071 18275
rect 16758 18272 16764 18284
rect 15059 18244 15148 18272
rect 16719 18244 16764 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 15120 18216 15148 18244
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 17957 18275 18015 18281
rect 17957 18241 17969 18275
rect 18003 18241 18015 18275
rect 17957 18235 18015 18241
rect 2501 18207 2559 18213
rect 2501 18173 2513 18207
rect 2547 18173 2559 18207
rect 2501 18167 2559 18173
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18204 2743 18207
rect 2866 18204 2872 18216
rect 2731 18176 2872 18204
rect 2731 18173 2743 18176
rect 2685 18167 2743 18173
rect 2516 18136 2544 18167
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 2958 18164 2964 18216
rect 3016 18204 3022 18216
rect 3016 18176 3061 18204
rect 3016 18164 3022 18176
rect 14826 18164 14832 18216
rect 14884 18204 14890 18216
rect 15102 18204 15108 18216
rect 14884 18176 15108 18204
rect 14884 18164 14890 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 17972 18204 18000 18235
rect 18414 18232 18420 18284
rect 18472 18272 18478 18284
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 18472 18244 18613 18272
rect 18472 18232 18478 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 20898 18272 20904 18284
rect 18601 18235 18659 18241
rect 20272 18244 20904 18272
rect 20272 18204 20300 18244
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 21085 18275 21143 18281
rect 21085 18272 21097 18275
rect 21048 18244 21097 18272
rect 21048 18232 21054 18244
rect 21085 18241 21097 18244
rect 21131 18272 21143 18275
rect 22186 18272 22192 18284
rect 21131 18244 21220 18272
rect 22147 18244 22192 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 21192 18216 21220 18244
rect 22186 18232 22192 18244
rect 22244 18232 22250 18284
rect 24670 18232 24676 18284
rect 24728 18272 24734 18284
rect 24765 18275 24823 18281
rect 24765 18272 24777 18275
rect 24728 18244 24777 18272
rect 24728 18232 24734 18244
rect 24765 18241 24777 18244
rect 24811 18241 24823 18275
rect 24946 18272 24952 18284
rect 24907 18244 24952 18272
rect 24765 18235 24823 18241
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 20438 18204 20444 18216
rect 16080 18176 20300 18204
rect 20399 18176 20444 18204
rect 16080 18164 16086 18176
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 21174 18164 21180 18216
rect 21232 18164 21238 18216
rect 23198 18164 23204 18216
rect 23256 18204 23262 18216
rect 26206 18204 26234 18312
rect 27614 18272 27620 18284
rect 27575 18244 27620 18272
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 28258 18272 28264 18284
rect 28219 18244 28264 18272
rect 28258 18232 28264 18244
rect 28316 18232 28322 18284
rect 30208 18281 30236 18312
rect 30374 18300 30380 18352
rect 30432 18340 30438 18352
rect 32324 18340 32352 18380
rect 44174 18368 44180 18380
rect 44232 18368 44238 18420
rect 47670 18408 47676 18420
rect 47631 18380 47676 18408
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 45646 18340 45652 18352
rect 30432 18312 32352 18340
rect 35866 18312 45652 18340
rect 30432 18300 30438 18312
rect 30852 18281 30880 18312
rect 30193 18275 30251 18281
rect 30193 18241 30205 18275
rect 30239 18241 30251 18275
rect 30193 18235 30251 18241
rect 30837 18275 30895 18281
rect 30837 18241 30849 18275
rect 30883 18241 30895 18275
rect 30837 18235 30895 18241
rect 32309 18275 32367 18281
rect 32309 18241 32321 18275
rect 32355 18272 32367 18275
rect 32398 18272 32404 18284
rect 32355 18244 32404 18272
rect 32355 18241 32367 18244
rect 32309 18235 32367 18241
rect 23256 18176 26234 18204
rect 30208 18204 30236 18235
rect 32398 18232 32404 18244
rect 32456 18232 32462 18284
rect 35866 18204 35894 18312
rect 45646 18300 45652 18312
rect 45704 18300 45710 18352
rect 45830 18340 45836 18352
rect 45791 18312 45836 18340
rect 45830 18300 45836 18312
rect 45888 18300 45894 18352
rect 40405 18275 40463 18281
rect 40405 18241 40417 18275
rect 40451 18272 40463 18275
rect 40494 18272 40500 18284
rect 40451 18244 40500 18272
rect 40451 18241 40463 18244
rect 40405 18235 40463 18241
rect 40494 18232 40500 18244
rect 40552 18232 40558 18284
rect 40589 18275 40647 18281
rect 40589 18241 40601 18275
rect 40635 18272 40647 18275
rect 40678 18272 40684 18284
rect 40635 18244 40684 18272
rect 40635 18241 40647 18244
rect 40589 18235 40647 18241
rect 40678 18232 40684 18244
rect 40736 18232 40742 18284
rect 40954 18232 40960 18284
rect 41012 18272 41018 18284
rect 41325 18275 41383 18281
rect 41325 18272 41337 18275
rect 41012 18244 41337 18272
rect 41012 18232 41018 18244
rect 41325 18241 41337 18244
rect 41371 18241 41383 18275
rect 42702 18272 42708 18284
rect 42663 18244 42708 18272
rect 41325 18235 41383 18241
rect 42702 18232 42708 18244
rect 42760 18232 42766 18284
rect 43714 18272 43720 18284
rect 42812 18244 43720 18272
rect 30208 18176 35894 18204
rect 23256 18164 23262 18176
rect 41046 18164 41052 18216
rect 41104 18204 41110 18216
rect 41601 18207 41659 18213
rect 41601 18204 41613 18207
rect 41104 18176 41613 18204
rect 41104 18164 41110 18176
rect 41601 18173 41613 18176
rect 41647 18173 41659 18207
rect 42812 18204 42840 18244
rect 43714 18232 43720 18244
rect 43772 18232 43778 18284
rect 46842 18272 46848 18284
rect 46803 18244 46848 18272
rect 46842 18232 46848 18244
rect 46900 18232 46906 18284
rect 47210 18232 47216 18284
rect 47268 18272 47274 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47268 18244 47593 18272
rect 47268 18232 47274 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 42720 18196 42840 18204
rect 41601 18167 41659 18173
rect 42536 18176 42840 18196
rect 42889 18207 42947 18213
rect 42536 18168 42748 18176
rect 42889 18173 42901 18207
rect 42935 18173 42947 18207
rect 43438 18204 43444 18216
rect 43399 18176 43444 18204
rect 28997 18139 29055 18145
rect 28997 18136 29009 18139
rect 2516 18108 29009 18136
rect 28997 18105 29009 18108
rect 29043 18136 29055 18139
rect 29638 18136 29644 18148
rect 29043 18108 29644 18136
rect 29043 18105 29055 18108
rect 28997 18099 29055 18105
rect 29638 18096 29644 18108
rect 29696 18096 29702 18148
rect 42536 18136 42564 18168
rect 42889 18167 42947 18173
rect 42904 18136 42932 18167
rect 43438 18164 43444 18176
rect 43496 18164 43502 18216
rect 43990 18204 43996 18216
rect 43951 18176 43996 18204
rect 43990 18164 43996 18176
rect 44048 18164 44054 18216
rect 44174 18204 44180 18216
rect 44135 18176 44180 18204
rect 44174 18164 44180 18176
rect 44232 18164 44238 18216
rect 31128 18108 42564 18136
rect 42720 18108 42932 18136
rect 43456 18136 43484 18164
rect 44082 18136 44088 18148
rect 43456 18108 44088 18136
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 14277 18071 14335 18077
rect 14277 18068 14289 18071
rect 13412 18040 14289 18068
rect 13412 18028 13418 18040
rect 14277 18037 14289 18040
rect 14323 18037 14335 18071
rect 14277 18031 14335 18037
rect 16666 18028 16672 18080
rect 16724 18068 16730 18080
rect 16945 18071 17003 18077
rect 16945 18068 16957 18071
rect 16724 18040 16957 18068
rect 16724 18028 16730 18040
rect 16945 18037 16957 18040
rect 16991 18037 17003 18071
rect 16945 18031 17003 18037
rect 30285 18071 30343 18077
rect 30285 18037 30297 18071
rect 30331 18068 30343 18071
rect 30742 18068 30748 18080
rect 30331 18040 30748 18068
rect 30331 18037 30343 18040
rect 30285 18031 30343 18037
rect 30742 18028 30748 18040
rect 30800 18028 30806 18080
rect 31128 18077 31156 18108
rect 31113 18071 31171 18077
rect 31113 18037 31125 18071
rect 31159 18037 31171 18071
rect 31113 18031 31171 18037
rect 31297 18071 31355 18077
rect 31297 18037 31309 18071
rect 31343 18068 31355 18071
rect 32398 18068 32404 18080
rect 31343 18040 32404 18068
rect 31343 18037 31355 18040
rect 31297 18031 31355 18037
rect 32398 18028 32404 18040
rect 32456 18028 32462 18080
rect 40405 18071 40463 18077
rect 40405 18037 40417 18071
rect 40451 18068 40463 18071
rect 41322 18068 41328 18080
rect 40451 18040 41328 18068
rect 40451 18037 40463 18040
rect 40405 18031 40463 18037
rect 41322 18028 41328 18040
rect 41380 18068 41386 18080
rect 41417 18071 41475 18077
rect 41417 18068 41429 18071
rect 41380 18040 41429 18068
rect 41380 18028 41386 18040
rect 41417 18037 41429 18040
rect 41463 18037 41475 18071
rect 41417 18031 41475 18037
rect 41509 18071 41567 18077
rect 41509 18037 41521 18071
rect 41555 18068 41567 18071
rect 42720 18068 42748 18108
rect 44082 18096 44088 18108
rect 44140 18096 44146 18148
rect 46934 18068 46940 18080
rect 41555 18040 42748 18068
rect 46895 18040 46940 18068
rect 41555 18037 41567 18040
rect 41509 18031 41567 18037
rect 46934 18028 46940 18040
rect 46992 18028 46998 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 14090 17824 14096 17876
rect 14148 17864 14154 17876
rect 14826 17864 14832 17876
rect 14148 17836 14832 17864
rect 14148 17824 14154 17836
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 21450 17864 21456 17876
rect 21411 17836 21456 17864
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 24302 17824 24308 17876
rect 24360 17864 24366 17876
rect 24397 17867 24455 17873
rect 24397 17864 24409 17867
rect 24360 17836 24409 17864
rect 24360 17824 24366 17836
rect 24397 17833 24409 17836
rect 24443 17833 24455 17867
rect 41322 17864 41328 17876
rect 24397 17827 24455 17833
rect 40880 17836 41328 17864
rect 28810 17728 28816 17740
rect 12406 17700 28816 17728
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17660 2835 17663
rect 2866 17660 2872 17672
rect 2823 17632 2872 17660
rect 2823 17629 2835 17632
rect 2777 17623 2835 17629
rect 2866 17620 2872 17632
rect 2924 17660 2930 17672
rect 12406 17660 12434 17700
rect 28810 17688 28816 17700
rect 28868 17688 28874 17740
rect 30742 17728 30748 17740
rect 30703 17700 30748 17728
rect 30742 17688 30748 17700
rect 30800 17688 30806 17740
rect 40773 17731 40831 17737
rect 40773 17697 40785 17731
rect 40819 17728 40831 17731
rect 40880 17728 40908 17836
rect 41322 17824 41328 17836
rect 41380 17864 41386 17876
rect 41380 17836 42196 17864
rect 41380 17824 41386 17836
rect 41046 17796 41052 17808
rect 41007 17768 41052 17796
rect 41046 17756 41052 17768
rect 41104 17796 41110 17808
rect 41104 17768 41920 17796
rect 41104 17756 41110 17768
rect 41690 17728 41696 17740
rect 40819 17700 40908 17728
rect 41651 17700 41696 17728
rect 40819 17697 40831 17700
rect 40773 17691 40831 17697
rect 41690 17688 41696 17700
rect 41748 17688 41754 17740
rect 2924 17632 12434 17660
rect 14737 17663 14795 17669
rect 2924 17620 2930 17632
rect 14737 17629 14749 17663
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 14752 17592 14780 17623
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 16390 17660 16396 17672
rect 14884 17632 14929 17660
rect 16351 17632 16396 17660
rect 14884 17620 14890 17632
rect 16390 17620 16396 17632
rect 16448 17620 16454 17672
rect 22922 17620 22928 17672
rect 22980 17660 22986 17672
rect 24581 17663 24639 17669
rect 24581 17660 24593 17663
rect 22980 17632 24593 17660
rect 22980 17620 22986 17632
rect 24581 17629 24593 17632
rect 24627 17660 24639 17663
rect 26878 17660 26884 17672
rect 24627 17632 26884 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 26878 17620 26884 17632
rect 26936 17620 26942 17672
rect 27614 17660 27620 17672
rect 27575 17632 27620 17660
rect 27614 17620 27620 17632
rect 27672 17620 27678 17672
rect 27982 17660 27988 17672
rect 27943 17632 27988 17660
rect 27982 17620 27988 17632
rect 28040 17620 28046 17672
rect 28166 17620 28172 17672
rect 28224 17660 28230 17672
rect 28261 17663 28319 17669
rect 28261 17660 28273 17663
rect 28224 17632 28273 17660
rect 28224 17620 28230 17632
rect 28261 17629 28273 17632
rect 28307 17629 28319 17663
rect 28626 17660 28632 17672
rect 28587 17632 28632 17660
rect 28261 17623 28319 17629
rect 28626 17620 28632 17632
rect 28684 17620 28690 17672
rect 41892 17669 41920 17768
rect 42168 17669 42196 17836
rect 43898 17824 43904 17876
rect 43956 17864 43962 17876
rect 45373 17867 45431 17873
rect 45373 17864 45385 17867
rect 43956 17836 45385 17864
rect 43956 17824 43962 17836
rect 45373 17833 45385 17836
rect 45419 17833 45431 17867
rect 45373 17827 45431 17833
rect 42242 17756 42248 17808
rect 42300 17796 42306 17808
rect 44174 17796 44180 17808
rect 42300 17768 42345 17796
rect 44135 17768 44180 17796
rect 42300 17756 42306 17768
rect 44174 17756 44180 17768
rect 44232 17756 44238 17808
rect 43714 17688 43720 17740
rect 43772 17728 43778 17740
rect 46477 17731 46535 17737
rect 43772 17700 43944 17728
rect 43772 17688 43778 17700
rect 30561 17663 30619 17669
rect 30561 17660 30573 17663
rect 28736 17632 30573 17660
rect 15194 17592 15200 17604
rect 14752 17564 15200 17592
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 16577 17595 16635 17601
rect 16577 17561 16589 17595
rect 16623 17592 16635 17595
rect 16758 17592 16764 17604
rect 16623 17564 16764 17592
rect 16623 17561 16635 17564
rect 16577 17555 16635 17561
rect 16758 17552 16764 17564
rect 16816 17552 16822 17604
rect 18230 17592 18236 17604
rect 18191 17564 18236 17592
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 21174 17592 21180 17604
rect 21135 17564 21180 17592
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 28736 17592 28764 17632
rect 30561 17629 30573 17632
rect 30607 17629 30619 17663
rect 30561 17623 30619 17629
rect 41877 17663 41935 17669
rect 41877 17629 41889 17663
rect 41923 17629 41935 17663
rect 41877 17623 41935 17629
rect 42153 17663 42211 17669
rect 42153 17629 42165 17663
rect 42199 17629 42211 17663
rect 43806 17660 43812 17672
rect 43767 17632 43812 17660
rect 42153 17623 42211 17629
rect 43806 17620 43812 17632
rect 43864 17620 43870 17672
rect 43916 17669 43944 17700
rect 46477 17697 46489 17731
rect 46523 17728 46535 17731
rect 46934 17728 46940 17740
rect 46523 17700 46940 17728
rect 46523 17697 46535 17700
rect 46477 17691 46535 17697
rect 46934 17688 46940 17700
rect 46992 17688 46998 17740
rect 43901 17663 43959 17669
rect 43901 17629 43913 17663
rect 43947 17629 43959 17663
rect 44266 17660 44272 17672
rect 44227 17632 44272 17660
rect 43901 17623 43959 17629
rect 44266 17620 44272 17632
rect 44324 17620 44330 17672
rect 45002 17660 45008 17672
rect 44963 17632 45008 17660
rect 45002 17620 45008 17632
rect 45060 17620 45066 17672
rect 46290 17660 46296 17672
rect 46251 17632 46296 17660
rect 46290 17620 46296 17632
rect 46348 17620 46354 17672
rect 23072 17564 28764 17592
rect 28905 17595 28963 17601
rect 23072 17552 23078 17564
rect 28905 17561 28917 17595
rect 28951 17561 28963 17595
rect 32398 17592 32404 17604
rect 32359 17564 32404 17592
rect 28905 17555 28963 17561
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2225 17527 2283 17533
rect 2225 17524 2237 17527
rect 2004 17496 2237 17524
rect 2004 17484 2010 17496
rect 2225 17493 2237 17496
rect 2271 17493 2283 17527
rect 15010 17524 15016 17536
rect 14971 17496 15016 17524
rect 2225 17487 2283 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 28920 17524 28948 17555
rect 32398 17552 32404 17564
rect 32456 17552 32462 17604
rect 42521 17595 42579 17601
rect 40972 17564 41414 17592
rect 40972 17536 41000 17564
rect 40954 17524 40960 17536
rect 28920 17496 40960 17524
rect 40954 17484 40960 17496
rect 41012 17484 41018 17536
rect 41230 17524 41236 17536
rect 41191 17496 41236 17524
rect 41230 17484 41236 17496
rect 41288 17484 41294 17536
rect 41386 17524 41414 17564
rect 42521 17561 42533 17595
rect 42567 17561 42579 17595
rect 42521 17555 42579 17561
rect 45189 17595 45247 17601
rect 45189 17561 45201 17595
rect 45235 17592 45247 17595
rect 45278 17592 45284 17604
rect 45235 17564 45284 17592
rect 45235 17561 45247 17564
rect 45189 17555 45247 17561
rect 42536 17524 42564 17555
rect 45278 17552 45284 17564
rect 45336 17552 45342 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 42610 17524 42616 17536
rect 41386 17496 42616 17524
rect 42610 17484 42616 17496
rect 42668 17484 42674 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 16758 17320 16764 17332
rect 16719 17292 16764 17320
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 24121 17323 24179 17329
rect 24121 17320 24133 17323
rect 22066 17292 24133 17320
rect 1946 17252 1952 17264
rect 1907 17224 1952 17252
rect 1946 17212 1952 17224
rect 2004 17212 2010 17264
rect 15194 17212 15200 17264
rect 15252 17252 15258 17264
rect 22066 17252 22094 17292
rect 24121 17289 24133 17292
rect 24167 17289 24179 17323
rect 24121 17283 24179 17289
rect 24302 17280 24308 17332
rect 24360 17320 24366 17332
rect 24762 17320 24768 17332
rect 24360 17292 24768 17320
rect 24360 17280 24366 17292
rect 24762 17280 24768 17292
rect 24820 17320 24826 17332
rect 25133 17323 25191 17329
rect 25133 17320 25145 17323
rect 24820 17292 25145 17320
rect 24820 17280 24826 17292
rect 25133 17289 25145 17292
rect 25179 17289 25191 17323
rect 25133 17283 25191 17289
rect 27614 17280 27620 17332
rect 27672 17280 27678 17332
rect 32398 17280 32404 17332
rect 32456 17320 32462 17332
rect 41782 17320 41788 17332
rect 32456 17292 41788 17320
rect 32456 17280 32462 17292
rect 41782 17280 41788 17292
rect 41840 17280 41846 17332
rect 15252 17224 22094 17252
rect 15252 17212 15258 17224
rect 22186 17212 22192 17264
rect 22244 17252 22250 17264
rect 23109 17255 23167 17261
rect 23109 17252 23121 17255
rect 22244 17224 23121 17252
rect 22244 17212 22250 17224
rect 23109 17221 23121 17224
rect 23155 17221 23167 17255
rect 24213 17255 24271 17261
rect 24213 17252 24225 17255
rect 23109 17215 23167 17221
rect 23492 17224 24225 17252
rect 14550 17184 14556 17196
rect 14511 17156 14556 17184
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 15102 17184 15108 17196
rect 15063 17156 15108 17184
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 16666 17184 16672 17196
rect 16627 17156 16672 17184
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17184 20223 17187
rect 21174 17184 21180 17196
rect 20211 17156 21180 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 21174 17144 21180 17156
rect 21232 17144 21238 17196
rect 22922 17184 22928 17196
rect 22883 17156 22928 17184
rect 22922 17144 22928 17156
rect 22980 17144 22986 17196
rect 23017 17187 23075 17193
rect 23017 17153 23029 17187
rect 23063 17184 23075 17187
rect 23290 17184 23296 17196
rect 23063 17156 23296 17184
rect 23063 17153 23075 17156
rect 23017 17147 23075 17153
rect 23290 17144 23296 17156
rect 23348 17184 23354 17196
rect 23492 17184 23520 17224
rect 24213 17221 24225 17224
rect 24259 17221 24271 17255
rect 26234 17252 26240 17264
rect 24213 17215 24271 17221
rect 25056 17224 26240 17252
rect 23348 17156 23520 17184
rect 24029 17187 24087 17193
rect 23348 17144 23354 17156
rect 24029 17153 24041 17187
rect 24075 17184 24087 17187
rect 24302 17184 24308 17196
rect 24075 17156 24308 17184
rect 24075 17153 24087 17156
rect 24029 17147 24087 17153
rect 24302 17144 24308 17156
rect 24360 17144 24366 17196
rect 24946 17144 24952 17196
rect 25004 17184 25010 17196
rect 25056 17193 25084 17224
rect 26234 17212 26240 17224
rect 26292 17212 26298 17264
rect 27632 17252 27660 17280
rect 45373 17255 45431 17261
rect 27632 17224 28014 17252
rect 45373 17221 45385 17255
rect 45419 17252 45431 17255
rect 47673 17255 47731 17261
rect 47673 17252 47685 17255
rect 45419 17224 47685 17252
rect 45419 17221 45431 17224
rect 45373 17215 45431 17221
rect 47673 17221 47685 17224
rect 47719 17221 47731 17255
rect 47673 17215 47731 17221
rect 25041 17187 25099 17193
rect 25041 17184 25053 17187
rect 25004 17156 25053 17184
rect 25004 17144 25010 17156
rect 25041 17153 25053 17156
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17153 25283 17187
rect 25225 17147 25283 17153
rect 25869 17187 25927 17193
rect 25869 17153 25881 17187
rect 25915 17184 25927 17187
rect 25958 17184 25964 17196
rect 25915 17156 25964 17184
rect 25915 17153 25927 17156
rect 25869 17147 25927 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 2038 17116 2044 17128
rect 1811 17088 2044 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2774 17076 2780 17128
rect 2832 17116 2838 17128
rect 2832 17088 2877 17116
rect 2832 17076 2838 17088
rect 3510 17076 3516 17128
rect 3568 17116 3574 17128
rect 9030 17116 9036 17128
rect 3568 17088 9036 17116
rect 3568 17076 3574 17088
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 14826 17076 14832 17128
rect 14884 17116 14890 17128
rect 14884 17088 23336 17116
rect 14884 17076 14890 17088
rect 17678 17008 17684 17060
rect 17736 17048 17742 17060
rect 21082 17048 21088 17060
rect 17736 17020 21088 17048
rect 17736 17008 17742 17020
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 22002 17008 22008 17060
rect 22060 17048 22066 17060
rect 23308 17057 23336 17088
rect 24394 17076 24400 17128
rect 24452 17116 24458 17128
rect 24578 17116 24584 17128
rect 24452 17088 24584 17116
rect 24452 17076 24458 17088
rect 24578 17076 24584 17088
rect 24636 17116 24642 17128
rect 25240 17116 25268 17147
rect 25958 17144 25964 17156
rect 26016 17144 26022 17196
rect 26878 17144 26884 17196
rect 26936 17184 26942 17196
rect 27065 17187 27123 17193
rect 27065 17184 27077 17187
rect 26936 17156 27077 17184
rect 26936 17144 26942 17156
rect 27065 17153 27077 17156
rect 27111 17153 27123 17187
rect 27065 17147 27123 17153
rect 27154 17144 27160 17196
rect 27212 17184 27218 17196
rect 27617 17187 27675 17193
rect 27617 17184 27629 17187
rect 27212 17156 27629 17184
rect 27212 17144 27218 17156
rect 27617 17153 27629 17156
rect 27663 17153 27675 17187
rect 42610 17184 42616 17196
rect 42571 17156 42616 17184
rect 27617 17147 27675 17153
rect 42610 17144 42616 17156
rect 42668 17144 42674 17196
rect 47581 17187 47639 17193
rect 47581 17153 47593 17187
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 24636 17088 25268 17116
rect 24636 17076 24642 17088
rect 41230 17076 41236 17128
rect 41288 17116 41294 17128
rect 42521 17119 42579 17125
rect 42521 17116 42533 17119
rect 41288 17088 42533 17116
rect 41288 17076 41294 17088
rect 42521 17085 42533 17088
rect 42567 17085 42579 17119
rect 42521 17079 42579 17085
rect 45189 17119 45247 17125
rect 45189 17085 45201 17119
rect 45235 17116 45247 17119
rect 46382 17116 46388 17128
rect 45235 17088 46388 17116
rect 45235 17085 45247 17088
rect 45189 17079 45247 17085
rect 46382 17076 46388 17088
rect 46440 17076 46446 17128
rect 46842 17116 46848 17128
rect 46803 17088 46848 17116
rect 46842 17076 46848 17088
rect 46900 17076 46906 17128
rect 22741 17051 22799 17057
rect 22741 17048 22753 17051
rect 22060 17020 22753 17048
rect 22060 17008 22066 17020
rect 22741 17017 22753 17020
rect 22787 17017 22799 17051
rect 22741 17011 22799 17017
rect 23293 17051 23351 17057
rect 23293 17017 23305 17051
rect 23339 17017 23351 17051
rect 23293 17011 23351 17017
rect 23845 17051 23903 17057
rect 23845 17017 23857 17051
rect 23891 17048 23903 17051
rect 24857 17051 24915 17057
rect 24857 17048 24869 17051
rect 23891 17020 24869 17048
rect 23891 17017 23903 17020
rect 23845 17011 23903 17017
rect 24857 17017 24869 17020
rect 24903 17048 24915 17051
rect 25038 17048 25044 17060
rect 24903 17020 25044 17048
rect 24903 17017 24915 17020
rect 24857 17011 24915 17017
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 14369 16983 14427 16989
rect 14369 16980 14381 16983
rect 14148 16952 14381 16980
rect 14148 16940 14154 16952
rect 14369 16949 14381 16952
rect 14415 16949 14427 16983
rect 14369 16943 14427 16949
rect 15197 16983 15255 16989
rect 15197 16949 15209 16983
rect 15243 16980 15255 16983
rect 15378 16980 15384 16992
rect 15243 16952 15384 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 22756 16980 22784 17011
rect 23860 16980 23888 17011
rect 25038 17008 25044 17020
rect 25096 17008 25102 17060
rect 42978 17048 42984 17060
rect 42939 17020 42984 17048
rect 42978 17008 42984 17020
rect 43036 17008 43042 17060
rect 44542 17008 44548 17060
rect 44600 17048 44606 17060
rect 45462 17048 45468 17060
rect 44600 17020 45468 17048
rect 44600 17008 44606 17020
rect 45462 17008 45468 17020
rect 45520 17048 45526 17060
rect 47596 17048 47624 17147
rect 45520 17020 47624 17048
rect 45520 17008 45526 17020
rect 24394 16980 24400 16992
rect 22756 16952 23888 16980
rect 24355 16952 24400 16980
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 24670 16940 24676 16992
rect 24728 16980 24734 16992
rect 25409 16983 25467 16989
rect 25409 16980 25421 16983
rect 24728 16952 25421 16980
rect 24728 16940 24734 16952
rect 25409 16949 25421 16952
rect 25455 16949 25467 16983
rect 26050 16980 26056 16992
rect 26011 16952 26056 16980
rect 25409 16943 25467 16949
rect 26050 16940 26056 16952
rect 26108 16940 26114 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 14608 16748 18460 16776
rect 14608 16736 14614 16748
rect 14090 16640 14096 16652
rect 14051 16612 14096 16640
rect 14090 16600 14096 16612
rect 14148 16600 14154 16652
rect 17402 16600 17408 16652
rect 17460 16640 17466 16652
rect 17678 16640 17684 16652
rect 17460 16612 17684 16640
rect 17460 16600 17466 16612
rect 17678 16600 17684 16612
rect 17736 16600 17742 16652
rect 17954 16640 17960 16652
rect 17915 16612 17960 16640
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 18432 16584 18460 16748
rect 21082 16736 21088 16788
rect 21140 16776 21146 16788
rect 24394 16776 24400 16788
rect 21140 16748 24400 16776
rect 21140 16736 21146 16748
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 27249 16779 27307 16785
rect 27249 16745 27261 16779
rect 27295 16776 27307 16779
rect 28626 16776 28632 16788
rect 27295 16748 28632 16776
rect 27295 16745 27307 16748
rect 27249 16739 27307 16745
rect 28626 16736 28632 16748
rect 28684 16736 28690 16788
rect 46290 16736 46296 16788
rect 46348 16776 46354 16788
rect 47673 16779 47731 16785
rect 47673 16776 47685 16779
rect 46348 16748 47685 16776
rect 46348 16736 46354 16748
rect 47673 16745 47685 16748
rect 47719 16745 47731 16779
rect 47673 16739 47731 16745
rect 23753 16711 23811 16717
rect 23753 16677 23765 16711
rect 23799 16708 23811 16711
rect 24581 16711 24639 16717
rect 24581 16708 24593 16711
rect 23799 16680 24593 16708
rect 23799 16677 23811 16680
rect 23753 16671 23811 16677
rect 24581 16677 24593 16680
rect 24627 16677 24639 16711
rect 24581 16671 24639 16677
rect 24670 16668 24676 16720
rect 24728 16668 24734 16720
rect 24762 16668 24768 16720
rect 24820 16668 24826 16720
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 23385 16643 23443 16649
rect 23385 16640 23397 16643
rect 22152 16612 23397 16640
rect 22152 16600 22158 16612
rect 23385 16609 23397 16612
rect 23431 16640 23443 16643
rect 24688 16640 24716 16668
rect 23431 16612 24716 16640
rect 24780 16640 24808 16668
rect 24857 16643 24915 16649
rect 24857 16640 24869 16643
rect 24780 16612 24869 16640
rect 23431 16609 23443 16612
rect 23385 16603 23443 16609
rect 24857 16609 24869 16612
rect 24903 16609 24915 16643
rect 25038 16640 25044 16652
rect 24999 16612 25044 16640
rect 24857 16603 24915 16609
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 26878 16640 26884 16652
rect 26839 16612 26884 16640
rect 26878 16600 26884 16612
rect 26936 16640 26942 16652
rect 27154 16640 27160 16652
rect 26936 16612 27160 16640
rect 26936 16600 26942 16612
rect 27154 16600 27160 16612
rect 27212 16600 27218 16652
rect 42978 16600 42984 16652
rect 43036 16640 43042 16652
rect 43990 16640 43996 16652
rect 43036 16612 43996 16640
rect 43036 16600 43042 16612
rect 43990 16600 43996 16612
rect 44048 16640 44054 16652
rect 45005 16643 45063 16649
rect 45005 16640 45017 16643
rect 44048 16612 45017 16640
rect 44048 16600 44054 16612
rect 45005 16609 45017 16612
rect 45051 16609 45063 16643
rect 45462 16640 45468 16652
rect 45423 16612 45468 16640
rect 45005 16603 45063 16609
rect 45462 16600 45468 16612
rect 45520 16600 45526 16652
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16572 17647 16575
rect 17862 16572 17868 16584
rect 17635 16544 17868 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 18414 16572 18420 16584
rect 18327 16544 18420 16572
rect 18414 16532 18420 16544
rect 18472 16532 18478 16584
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16572 19303 16575
rect 19426 16572 19432 16584
rect 19291 16544 19432 16572
rect 19291 16541 19303 16544
rect 19245 16535 19303 16541
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 21637 16575 21695 16581
rect 21637 16572 21649 16575
rect 21508 16544 21649 16572
rect 21508 16532 21514 16544
rect 21637 16541 21649 16544
rect 21683 16541 21695 16575
rect 21637 16535 21695 16541
rect 24578 16532 24584 16584
rect 24636 16572 24642 16584
rect 24765 16575 24823 16581
rect 24765 16572 24777 16575
rect 24636 16544 24777 16572
rect 24636 16532 24642 16544
rect 24765 16541 24777 16544
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 24946 16532 24952 16584
rect 25004 16572 25010 16584
rect 27062 16572 27068 16584
rect 25004 16544 25097 16572
rect 27023 16544 27068 16572
rect 25004 16532 25010 16544
rect 27062 16532 27068 16544
rect 27120 16532 27126 16584
rect 44269 16575 44327 16581
rect 44269 16541 44281 16575
rect 44315 16572 44327 16575
rect 44542 16572 44548 16584
rect 44315 16544 44548 16572
rect 44315 16541 44327 16544
rect 44269 16535 44327 16541
rect 44542 16532 44548 16544
rect 44600 16532 44606 16584
rect 14366 16504 14372 16516
rect 14327 16476 14372 16504
rect 14366 16464 14372 16476
rect 14424 16464 14430 16516
rect 15378 16464 15384 16516
rect 15436 16464 15442 16516
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 18288 16476 24072 16504
rect 18288 16464 18294 16476
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 15841 16439 15899 16445
rect 15841 16436 15853 16439
rect 15252 16408 15853 16436
rect 15252 16396 15258 16408
rect 15841 16405 15853 16408
rect 15887 16405 15899 16439
rect 18598 16436 18604 16448
rect 18559 16408 18604 16436
rect 15841 16399 15899 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 19334 16436 19340 16448
rect 19295 16408 19340 16436
rect 19334 16396 19340 16408
rect 19392 16396 19398 16448
rect 21818 16436 21824 16448
rect 21779 16408 21824 16436
rect 21818 16396 21824 16408
rect 21876 16396 21882 16448
rect 23842 16436 23848 16448
rect 23803 16408 23848 16436
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 24044 16436 24072 16476
rect 24210 16464 24216 16516
rect 24268 16504 24274 16516
rect 24964 16504 24992 16532
rect 24268 16476 24992 16504
rect 44361 16507 44419 16513
rect 24268 16464 24274 16476
rect 44361 16473 44373 16507
rect 44407 16504 44419 16507
rect 45189 16507 45247 16513
rect 45189 16504 45201 16507
rect 44407 16476 45201 16504
rect 44407 16473 44419 16476
rect 44361 16467 44419 16473
rect 45189 16473 45201 16476
rect 45235 16473 45247 16507
rect 45189 16467 45247 16473
rect 45554 16436 45560 16448
rect 24044 16408 45560 16436
rect 45554 16396 45560 16408
rect 45612 16396 45618 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 20346 16232 20352 16244
rect 18472 16204 20352 16232
rect 18472 16192 18478 16204
rect 15010 16164 15016 16176
rect 13832 16136 15016 16164
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 13740 15960 13768 16059
rect 13832 16037 13860 16136
rect 15010 16124 15016 16136
rect 15068 16164 15074 16176
rect 15068 16136 15516 16164
rect 15068 16124 15074 16136
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16096 14703 16099
rect 15102 16096 15108 16108
rect 14691 16068 15108 16096
rect 14691 16065 14703 16068
rect 14645 16059 14703 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 15488 16105 15516 16136
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 18049 16167 18107 16173
rect 18049 16164 18061 16167
rect 18012 16136 18061 16164
rect 18012 16124 18018 16136
rect 18049 16133 18061 16136
rect 18095 16133 18107 16167
rect 19334 16164 19340 16176
rect 19274 16136 19340 16164
rect 18049 16127 18107 16133
rect 19334 16124 19340 16136
rect 19392 16124 19398 16176
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16666 16096 16672 16108
rect 15979 16068 16672 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 13817 16031 13875 16037
rect 13817 15997 13829 16031
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 14366 16028 14372 16040
rect 14139 16000 14372 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15764 16028 15792 16059
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 20088 16105 20116 16204
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 23125 16235 23183 16241
rect 23125 16232 23137 16235
rect 23124 16201 23137 16232
rect 23171 16201 23183 16235
rect 23290 16232 23296 16244
rect 23251 16204 23296 16232
rect 23124 16195 23183 16201
rect 21358 16124 21364 16176
rect 21416 16164 21422 16176
rect 22925 16167 22983 16173
rect 22925 16164 22937 16167
rect 21416 16136 22937 16164
rect 21416 16124 21422 16136
rect 22925 16133 22937 16136
rect 22971 16133 22983 16167
rect 23124 16164 23152 16195
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 23753 16235 23811 16241
rect 23753 16201 23765 16235
rect 23799 16201 23811 16235
rect 23753 16195 23811 16201
rect 23768 16164 23796 16195
rect 25038 16192 25044 16244
rect 25096 16232 25102 16244
rect 26145 16235 26203 16241
rect 26145 16232 26157 16235
rect 25096 16204 26157 16232
rect 25096 16192 25102 16204
rect 26145 16201 26157 16204
rect 26191 16201 26203 16235
rect 26145 16195 26203 16201
rect 24673 16167 24731 16173
rect 24673 16164 24685 16167
rect 23124 16136 23704 16164
rect 23768 16136 24685 16164
rect 22925 16127 22983 16133
rect 20073 16099 20131 16105
rect 20073 16065 20085 16099
rect 20119 16065 20131 16099
rect 20073 16059 20131 16065
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 20990 16096 20996 16108
rect 20947 16068 20996 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21082 16056 21088 16108
rect 21140 16096 21146 16108
rect 21140 16068 21185 16096
rect 21140 16056 21146 16068
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21968 16068 22017 16096
rect 21968 16056 21974 16068
rect 22005 16065 22017 16068
rect 22051 16096 22063 16099
rect 22051 16068 23152 16096
rect 22051 16065 22063 16068
rect 22005 16059 22063 16065
rect 17586 16028 17592 16040
rect 15764 16000 17592 16028
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 17773 16031 17831 16037
rect 17773 15997 17785 16031
rect 17819 16028 17831 16031
rect 18598 16028 18604 16040
rect 17819 16000 18604 16028
rect 17819 15997 17831 16000
rect 17773 15991 17831 15997
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 22094 16028 22100 16040
rect 22055 16000 22100 16028
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 14458 15960 14464 15972
rect 13740 15932 14464 15960
rect 14458 15920 14464 15932
rect 14516 15960 14522 15972
rect 15102 15960 15108 15972
rect 14516 15932 15108 15960
rect 14516 15920 14522 15932
rect 15102 15920 15108 15932
rect 15160 15920 15166 15972
rect 14737 15895 14795 15901
rect 14737 15861 14749 15895
rect 14783 15892 14795 15895
rect 14918 15892 14924 15904
rect 14783 15864 14924 15892
rect 14783 15861 14795 15864
rect 14737 15855 14795 15861
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15010 15852 15016 15904
rect 15068 15892 15074 15904
rect 15289 15895 15347 15901
rect 15289 15892 15301 15895
rect 15068 15864 15301 15892
rect 15068 15852 15074 15864
rect 15289 15861 15301 15864
rect 15335 15861 15347 15895
rect 15289 15855 15347 15861
rect 17862 15852 17868 15904
rect 17920 15892 17926 15904
rect 19521 15895 19579 15901
rect 19521 15892 19533 15895
rect 17920 15864 19533 15892
rect 17920 15852 17926 15864
rect 19521 15861 19533 15864
rect 19567 15861 19579 15895
rect 19521 15855 19579 15861
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 20073 15895 20131 15901
rect 20073 15892 20085 15895
rect 19668 15864 20085 15892
rect 19668 15852 19674 15864
rect 20073 15861 20085 15864
rect 20119 15861 20131 15895
rect 20898 15892 20904 15904
rect 20859 15864 20904 15892
rect 20073 15855 20131 15861
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 23124 15901 23152 16068
rect 23676 16028 23704 16136
rect 24673 16133 24685 16136
rect 24719 16133 24731 16167
rect 24673 16127 24731 16133
rect 25314 16124 25320 16176
rect 25372 16124 25378 16176
rect 23842 16056 23848 16108
rect 23900 16096 23906 16108
rect 23937 16099 23995 16105
rect 23937 16096 23949 16099
rect 23900 16068 23949 16096
rect 23900 16056 23906 16068
rect 23937 16065 23949 16068
rect 23983 16065 23995 16099
rect 41230 16096 41236 16108
rect 41191 16068 41236 16096
rect 23937 16059 23995 16065
rect 41230 16056 41236 16068
rect 41288 16056 41294 16108
rect 46382 16056 46388 16108
rect 46440 16096 46446 16108
rect 47765 16099 47823 16105
rect 47765 16096 47777 16099
rect 46440 16068 47777 16096
rect 46440 16056 46446 16068
rect 47765 16065 47777 16068
rect 47811 16065 47823 16099
rect 47765 16059 47823 16065
rect 24210 16028 24216 16040
rect 23676 16000 24216 16028
rect 24210 15988 24216 16000
rect 24268 15988 24274 16040
rect 24394 16028 24400 16040
rect 24355 16000 24400 16028
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 22373 15895 22431 15901
rect 22373 15892 22385 15895
rect 22152 15864 22385 15892
rect 22152 15852 22158 15864
rect 22373 15861 22385 15864
rect 22419 15861 22431 15895
rect 22373 15855 22431 15861
rect 23109 15895 23167 15901
rect 23109 15861 23121 15895
rect 23155 15892 23167 15895
rect 23566 15892 23572 15904
rect 23155 15864 23572 15892
rect 23155 15861 23167 15864
rect 23109 15855 23167 15861
rect 23566 15852 23572 15864
rect 23624 15852 23630 15904
rect 41325 15895 41383 15901
rect 41325 15861 41337 15895
rect 41371 15892 41383 15895
rect 41414 15892 41420 15904
rect 41371 15864 41420 15892
rect 41371 15861 41383 15864
rect 41325 15855 41383 15861
rect 41414 15852 41420 15864
rect 41472 15852 41478 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 17770 15688 17776 15700
rect 17731 15660 17776 15688
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 17957 15691 18015 15697
rect 17957 15657 17969 15691
rect 18003 15688 18015 15691
rect 22278 15688 22284 15700
rect 18003 15660 22284 15688
rect 18003 15657 18015 15660
rect 17957 15651 18015 15657
rect 22278 15648 22284 15660
rect 22336 15648 22342 15700
rect 23566 15688 23572 15700
rect 23527 15660 23572 15688
rect 23566 15648 23572 15660
rect 23624 15648 23630 15700
rect 24394 15688 24400 15700
rect 24355 15660 24400 15688
rect 24394 15648 24400 15660
rect 24452 15648 24458 15700
rect 25314 15688 25320 15700
rect 25275 15660 25320 15688
rect 25314 15648 25320 15660
rect 25372 15648 25378 15700
rect 21358 15620 21364 15632
rect 21319 15592 21364 15620
rect 21358 15580 21364 15592
rect 21416 15580 21422 15632
rect 43438 15620 43444 15632
rect 41248 15592 43444 15620
rect 15010 15552 15016 15564
rect 14971 15524 15016 15552
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 19610 15552 19616 15564
rect 19571 15524 19616 15552
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 19889 15555 19947 15561
rect 19889 15521 19901 15555
rect 19935 15552 19947 15555
rect 20898 15552 20904 15564
rect 19935 15524 20904 15552
rect 19935 15521 19947 15524
rect 19889 15515 19947 15521
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 21818 15552 21824 15564
rect 21779 15524 21824 15552
rect 21818 15512 21824 15524
rect 21876 15512 21882 15564
rect 22094 15552 22100 15564
rect 22055 15524 22100 15552
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 41248 15561 41276 15592
rect 43438 15580 43444 15592
rect 43496 15580 43502 15632
rect 41233 15555 41291 15561
rect 41233 15521 41245 15555
rect 41279 15521 41291 15555
rect 41233 15515 41291 15521
rect 41414 15512 41420 15564
rect 41472 15552 41478 15564
rect 42886 15552 42892 15564
rect 41472 15524 41517 15552
rect 42847 15524 42892 15552
rect 41472 15512 41478 15524
rect 42886 15512 42892 15524
rect 42944 15512 42950 15564
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 14734 15484 14740 15496
rect 14695 15456 14740 15484
rect 2041 15447 2099 15453
rect 14734 15444 14740 15456
rect 14792 15444 14798 15496
rect 18414 15484 18420 15496
rect 18375 15456 18420 15484
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 23400 15456 24409 15484
rect 14918 15376 14924 15428
rect 14976 15416 14982 15428
rect 17862 15425 17868 15428
rect 17589 15419 17647 15425
rect 14976 15388 15502 15416
rect 14976 15376 14982 15388
rect 17589 15385 17601 15419
rect 17635 15385 17647 15419
rect 17589 15379 17647 15385
rect 17805 15419 17868 15425
rect 17805 15385 17817 15419
rect 17851 15385 17868 15419
rect 17805 15379 17868 15385
rect 16485 15351 16543 15357
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 16666 15348 16672 15360
rect 16531 15320 16672 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 16666 15308 16672 15320
rect 16724 15348 16730 15360
rect 17604 15348 17632 15379
rect 17862 15376 17868 15379
rect 17920 15376 17926 15428
rect 21174 15416 21180 15428
rect 21114 15388 21180 15416
rect 21174 15376 21180 15388
rect 21232 15376 21238 15428
rect 23106 15376 23112 15428
rect 23164 15376 23170 15428
rect 16724 15320 17632 15348
rect 16724 15308 16730 15320
rect 18046 15308 18052 15360
rect 18104 15348 18110 15360
rect 18601 15351 18659 15357
rect 18601 15348 18613 15351
rect 18104 15320 18613 15348
rect 18104 15308 18110 15320
rect 18601 15317 18613 15320
rect 18647 15317 18659 15351
rect 18601 15311 18659 15317
rect 21450 15308 21456 15360
rect 21508 15348 21514 15360
rect 23400 15348 23428 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 25222 15484 25228 15496
rect 25135 15456 25228 15484
rect 24397 15447 24455 15453
rect 25222 15444 25228 15456
rect 25280 15484 25286 15496
rect 26050 15484 26056 15496
rect 25280 15456 26056 15484
rect 25280 15444 25286 15456
rect 26050 15444 26056 15456
rect 26108 15444 26114 15496
rect 21508 15320 23428 15348
rect 21508 15308 21514 15320
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14792 15116 14933 15144
rect 14792 15104 14798 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 17402 15104 17408 15156
rect 17460 15153 17466 15156
rect 17460 15147 17479 15153
rect 17467 15113 17479 15147
rect 17586 15144 17592 15156
rect 17547 15116 17592 15144
rect 17460 15107 17479 15113
rect 17460 15104 17466 15107
rect 17586 15104 17592 15116
rect 17644 15104 17650 15156
rect 19797 15147 19855 15153
rect 19797 15144 19809 15147
rect 17788 15116 19809 15144
rect 17788 15088 17816 15116
rect 19797 15113 19809 15116
rect 19843 15113 19855 15147
rect 21174 15144 21180 15156
rect 21135 15116 21180 15144
rect 19797 15107 19855 15113
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 23017 15147 23075 15153
rect 23017 15113 23029 15147
rect 23063 15144 23075 15147
rect 23106 15144 23112 15156
rect 23063 15116 23112 15144
rect 23063 15113 23075 15116
rect 23017 15107 23075 15113
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 17221 15079 17279 15085
rect 17221 15045 17233 15079
rect 17267 15076 17279 15079
rect 17770 15076 17776 15088
rect 17267 15048 17776 15076
rect 17267 15045 17279 15048
rect 17221 15039 17279 15045
rect 17770 15036 17776 15048
rect 17828 15036 17834 15088
rect 21358 15036 21364 15088
rect 21416 15076 21422 15088
rect 21818 15076 21824 15088
rect 21416 15048 21824 15076
rect 21416 15036 21422 15048
rect 21818 15036 21824 15048
rect 21876 15036 21882 15088
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14737 15011 14795 15017
rect 14737 15008 14749 15011
rect 14608 14980 14749 15008
rect 14608 14968 14614 14980
rect 14737 14977 14749 14980
rect 14783 14977 14795 15011
rect 18046 15008 18052 15020
rect 18007 14980 18052 15008
rect 14737 14971 14795 14977
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 19426 14968 19432 15020
rect 19484 14968 19490 15020
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 18322 14940 18328 14952
rect 2832 14912 2877 14940
rect 18283 14912 18328 14940
rect 2832 14900 2838 14912
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 21100 14940 21128 14971
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22186 15008 22192 15020
rect 22143 14980 22192 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 22925 15011 22983 15017
rect 22925 14977 22937 15011
rect 22971 15008 22983 15011
rect 25222 15008 25228 15020
rect 22971 14980 25228 15008
rect 22971 14977 22983 14980
rect 22925 14971 22983 14977
rect 22940 14940 22968 14971
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 19392 14912 22968 14940
rect 19392 14900 19398 14912
rect 17862 14872 17868 14884
rect 17420 14844 17868 14872
rect 17420 14813 17448 14844
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 20990 14832 20996 14884
rect 21048 14872 21054 14884
rect 21821 14875 21879 14881
rect 21821 14872 21833 14875
rect 21048 14844 21833 14872
rect 21048 14832 21054 14844
rect 21821 14841 21833 14844
rect 21867 14841 21879 14875
rect 21821 14835 21879 14841
rect 17405 14807 17463 14813
rect 17405 14773 17417 14807
rect 17451 14773 17463 14807
rect 17405 14767 17463 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 18049 14603 18107 14609
rect 18049 14569 18061 14603
rect 18095 14600 18107 14603
rect 18322 14600 18328 14612
rect 18095 14572 18328 14600
rect 18095 14569 18107 14572
rect 18049 14563 18107 14569
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 19426 14600 19432 14612
rect 19387 14572 19432 14600
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 17402 14532 17408 14544
rect 16960 14504 17408 14532
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14396 2194 14408
rect 2866 14396 2872 14408
rect 2188 14368 2872 14396
rect 2188 14356 2194 14368
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 16960 14405 16988 14504
rect 17402 14492 17408 14504
rect 17460 14492 17466 14544
rect 17037 14467 17095 14473
rect 17037 14433 17049 14467
rect 17083 14464 17095 14467
rect 17681 14467 17739 14473
rect 17681 14464 17693 14467
rect 17083 14436 17693 14464
rect 17083 14433 17095 14436
rect 17037 14427 17095 14433
rect 17681 14433 17693 14436
rect 17727 14433 17739 14467
rect 17681 14427 17739 14433
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14365 17187 14399
rect 17770 14396 17776 14408
rect 17731 14368 17776 14396
rect 17129 14359 17187 14365
rect 17144 14328 17172 14359
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 19334 14396 19340 14408
rect 19295 14368 19340 14396
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 22189 14399 22247 14405
rect 22189 14365 22201 14399
rect 22235 14396 22247 14399
rect 22554 14396 22560 14408
rect 22235 14368 22560 14396
rect 22235 14365 22247 14368
rect 22189 14359 22247 14365
rect 22554 14356 22560 14368
rect 22612 14396 22618 14408
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22612 14368 22845 14396
rect 22612 14356 22618 14368
rect 22833 14365 22845 14368
rect 22879 14396 22891 14399
rect 30558 14396 30564 14408
rect 22879 14368 30564 14396
rect 22879 14365 22891 14368
rect 22833 14359 22891 14365
rect 30558 14356 30564 14368
rect 30616 14356 30622 14408
rect 17862 14328 17868 14340
rect 17144 14300 17868 14328
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 22278 14260 22284 14272
rect 22239 14232 22284 14260
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 22922 14260 22928 14272
rect 22883 14232 22928 14260
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 3694 13948 3700 14000
rect 3752 13988 3758 14000
rect 3752 13960 21772 13988
rect 3752 13948 3758 13960
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 15160 13892 16681 13920
rect 15160 13880 15166 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 18506 13852 18512 13864
rect 18467 13824 18512 13852
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 14274 13784 14280 13796
rect 4028 13756 14280 13784
rect 4028 13744 4034 13756
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 21744 13784 21772 13960
rect 21818 13948 21824 14000
rect 21876 13948 21882 14000
rect 22005 13991 22063 13997
rect 22005 13957 22017 13991
rect 22051 13988 22063 13991
rect 22922 13988 22928 14000
rect 22051 13960 22928 13988
rect 22051 13957 22063 13960
rect 22005 13951 22063 13957
rect 22922 13948 22928 13960
rect 22980 13948 22986 14000
rect 21836 13861 21864 13948
rect 45094 13880 45100 13932
rect 45152 13920 45158 13932
rect 46845 13923 46903 13929
rect 46845 13920 46857 13923
rect 45152 13892 46857 13920
rect 45152 13880 45158 13892
rect 46845 13889 46857 13892
rect 46891 13889 46903 13923
rect 46845 13883 46903 13889
rect 21821 13855 21879 13861
rect 21821 13821 21833 13855
rect 21867 13821 21879 13855
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 21821 13815 21879 13821
rect 21928 13824 22293 13852
rect 21928 13784 21956 13824
rect 22281 13821 22293 13824
rect 22327 13821 22339 13855
rect 22281 13815 22339 13821
rect 21744 13756 21956 13784
rect 46934 13716 46940 13728
rect 46895 13688 46940 13716
rect 46934 13676 46940 13688
rect 46992 13676 46998 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 15838 13472 15844 13524
rect 15896 13512 15902 13524
rect 24854 13512 24860 13524
rect 15896 13484 24860 13512
rect 15896 13472 15902 13484
rect 24854 13472 24860 13484
rect 24912 13472 24918 13524
rect 17770 13444 17776 13456
rect 16224 13416 17776 13444
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 16224 13308 16252 13416
rect 17770 13404 17776 13416
rect 17828 13404 17834 13456
rect 30466 13444 30472 13456
rect 22066 13416 30472 13444
rect 16942 13376 16948 13388
rect 16903 13348 16948 13376
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17954 13336 17960 13388
rect 18012 13376 18018 13388
rect 19429 13379 19487 13385
rect 19429 13376 19441 13379
rect 18012 13348 19441 13376
rect 18012 13336 18018 13348
rect 19429 13345 19441 13348
rect 19475 13345 19487 13379
rect 19429 13339 19487 13345
rect 21085 13379 21143 13385
rect 21085 13345 21097 13379
rect 21131 13376 21143 13379
rect 22066 13376 22094 13416
rect 30466 13404 30472 13416
rect 30524 13404 30530 13456
rect 22462 13376 22468 13388
rect 21131 13348 22094 13376
rect 22423 13348 22468 13376
rect 21131 13345 21143 13348
rect 21085 13339 21143 13345
rect 22462 13336 22468 13348
rect 22520 13336 22526 13388
rect 46477 13379 46535 13385
rect 46477 13345 46489 13379
rect 46523 13376 46535 13379
rect 46934 13376 46940 13388
rect 46523 13348 46940 13376
rect 46523 13345 46535 13348
rect 46477 13339 46535 13345
rect 46934 13336 46940 13348
rect 46992 13336 46998 13388
rect 16393 13311 16451 13317
rect 16393 13308 16405 13311
rect 16224 13280 16405 13308
rect 15749 13271 15807 13277
rect 16393 13277 16405 13280
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 15764 13172 15792 13271
rect 17862 13268 17868 13320
rect 17920 13308 17926 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 17920 13280 19257 13308
rect 17920 13268 17926 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 22002 13308 22008 13320
rect 21963 13280 22008 13308
rect 19245 13271 19303 13277
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 46290 13308 46296 13320
rect 46251 13280 46296 13308
rect 46290 13268 46296 13280
rect 46348 13268 46354 13320
rect 15841 13243 15899 13249
rect 15841 13209 15853 13243
rect 15887 13240 15899 13243
rect 16577 13243 16635 13249
rect 16577 13240 16589 13243
rect 15887 13212 16589 13240
rect 15887 13209 15899 13212
rect 15841 13203 15899 13209
rect 16577 13209 16589 13212
rect 16623 13209 16635 13243
rect 22186 13240 22192 13252
rect 22147 13212 22192 13240
rect 16577 13203 16635 13209
rect 22186 13200 22192 13212
rect 22244 13200 22250 13252
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 16758 13172 16764 13184
rect 15764 13144 16764 13172
rect 16758 13132 16764 13144
rect 16816 13132 16822 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 1596 12900 1624 12931
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 22462 12968 22468 12980
rect 3384 12940 22468 12968
rect 3384 12928 3390 12940
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 15838 12900 15844 12912
rect 1596 12872 15844 12900
rect 15838 12860 15844 12872
rect 15896 12860 15902 12912
rect 16025 12903 16083 12909
rect 16025 12869 16037 12903
rect 16071 12900 16083 12903
rect 16853 12903 16911 12909
rect 16853 12900 16865 12903
rect 16071 12872 16865 12900
rect 16071 12869 16083 12872
rect 16025 12863 16083 12869
rect 16853 12869 16865 12872
rect 16899 12869 16911 12903
rect 16853 12863 16911 12869
rect 22005 12903 22063 12909
rect 22005 12869 22017 12903
rect 22051 12900 22063 12903
rect 22278 12900 22284 12912
rect 22051 12872 22284 12900
rect 22051 12869 22063 12872
rect 22005 12863 22063 12869
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12801 15991 12835
rect 16666 12832 16672 12844
rect 16627 12804 16672 12832
rect 15933 12795 15991 12801
rect 15948 12764 15976 12795
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 21818 12832 21824 12844
rect 21779 12804 21824 12832
rect 21818 12792 21824 12804
rect 21876 12792 21882 12844
rect 46290 12792 46296 12844
rect 46348 12832 46354 12844
rect 47765 12835 47823 12841
rect 47765 12832 47777 12835
rect 46348 12804 47777 12832
rect 46348 12792 46354 12804
rect 47765 12801 47777 12804
rect 47811 12801 47823 12835
rect 47765 12795 47823 12801
rect 16574 12764 16580 12776
rect 15948 12736 16580 12764
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 22281 12767 22339 12773
rect 22281 12733 22293 12767
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 3510 12656 3516 12708
rect 3568 12696 3574 12708
rect 22296 12696 22324 12727
rect 3568 12668 22324 12696
rect 3568 12656 3574 12668
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 16942 12628 16948 12640
rect 14884 12600 16948 12628
rect 14884 12588 14890 12600
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 16761 12427 16819 12433
rect 16761 12393 16773 12427
rect 16807 12424 16819 12427
rect 16850 12424 16856 12436
rect 16807 12396 16856 12424
rect 16807 12393 16819 12396
rect 16761 12387 16819 12393
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 17773 12427 17831 12433
rect 17773 12393 17785 12427
rect 17819 12424 17831 12427
rect 17954 12424 17960 12436
rect 17819 12396 17960 12424
rect 17819 12393 17831 12396
rect 17773 12387 17831 12393
rect 17954 12384 17960 12396
rect 18012 12384 18018 12436
rect 22186 12384 22192 12436
rect 22244 12424 22250 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 22244 12396 22661 12424
rect 22244 12384 22250 12396
rect 22649 12393 22661 12396
rect 22695 12393 22707 12427
rect 22649 12387 22707 12393
rect 16669 12223 16727 12229
rect 16669 12189 16681 12223
rect 16715 12220 16727 12223
rect 16758 12220 16764 12232
rect 16715 12192 16764 12220
rect 16715 12189 16727 12192
rect 16669 12183 16727 12189
rect 16758 12180 16764 12192
rect 16816 12220 16822 12232
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 16816 12192 17693 12220
rect 16816 12180 16822 12192
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 22554 12220 22560 12232
rect 22515 12192 22560 12220
rect 17681 12183 17739 12189
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 46477 11067 46535 11073
rect 46477 11033 46489 11067
rect 46523 11064 46535 11067
rect 46934 11064 46940 11076
rect 46523 11036 46940 11064
rect 46523 11033 46535 11036
rect 46477 11027 46535 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 10778 10996 10784 11008
rect 3476 10968 10784 10996
rect 3476 10956 3482 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 46934 10792 46940 10804
rect 46895 10764 46940 10792
rect 46934 10752 46940 10764
rect 46992 10752 46998 10804
rect 45646 10616 45652 10668
rect 45704 10656 45710 10668
rect 46658 10656 46664 10668
rect 45704 10628 46664 10656
rect 45704 10616 45710 10628
rect 46658 10616 46664 10628
rect 46716 10656 46722 10668
rect 46845 10659 46903 10665
rect 46845 10656 46857 10659
rect 46716 10628 46857 10656
rect 46716 10616 46722 10628
rect 46845 10625 46857 10628
rect 46891 10625 46903 10659
rect 47578 10656 47584 10668
rect 47539 10628 47584 10656
rect 46845 10619 46903 10625
rect 47578 10616 47584 10628
rect 47636 10616 47642 10668
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 46385 10455 46443 10461
rect 46385 10452 46397 10455
rect 46348 10424 46397 10452
rect 46348 10412 46354 10424
rect 46385 10421 46397 10424
rect 46431 10421 46443 10455
rect 46385 10415 46443 10421
rect 46474 10412 46480 10464
rect 46532 10452 46538 10464
rect 47673 10455 47731 10461
rect 47673 10452 47685 10455
rect 46532 10424 47685 10452
rect 46532 10412 46538 10424
rect 47673 10421 47685 10424
rect 47719 10421 47731 10455
rect 47673 10415 47731 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 46474 10112 46480 10124
rect 46435 10084 46480 10112
rect 46474 10072 46480 10084
rect 46532 10072 46538 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 47854 9568 47860 9580
rect 47815 9540 47860 9568
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 46106 9392 46112 9444
rect 46164 9432 46170 9444
rect 48041 9435 48099 9441
rect 48041 9432 48053 9435
rect 46164 9404 48053 9432
rect 46164 9392 46170 9404
rect 48041 9401 48053 9404
rect 48087 9401 48099 9435
rect 48041 9395 48099 9401
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47762 8888 47768 8900
rect 47723 8860 47768 8888
rect 47762 8848 47768 8860
rect 47820 8848 47826 8900
rect 29730 8780 29736 8832
rect 29788 8820 29794 8832
rect 47857 8823 47915 8829
rect 47857 8820 47869 8823
rect 29788 8792 47869 8820
rect 29788 8780 29794 8792
rect 47857 8789 47869 8792
rect 47903 8789 47915 8823
rect 47857 8783 47915 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 45094 8480 45100 8492
rect 45055 8452 45100 8480
rect 45094 8440 45100 8452
rect 45152 8440 45158 8492
rect 44836 8316 45416 8344
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 18046 8276 18052 8288
rect 3476 8248 18052 8276
rect 3476 8236 3482 8248
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 44836 8276 44864 8316
rect 18564 8248 44864 8276
rect 44913 8279 44971 8285
rect 18564 8236 18570 8248
rect 44913 8245 44925 8279
rect 44959 8276 44971 8279
rect 45278 8276 45284 8288
rect 44959 8248 45284 8276
rect 44959 8245 44971 8248
rect 44913 8239 44971 8245
rect 45278 8236 45284 8248
rect 45336 8236 45342 8288
rect 45388 8276 45416 8316
rect 45554 8276 45560 8288
rect 45388 8248 45560 8276
rect 45554 8236 45560 8248
rect 45612 8236 45618 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 43625 8075 43683 8081
rect 43625 8072 43637 8075
rect 1912 8044 43637 8072
rect 1912 8032 1918 8044
rect 43625 8041 43637 8044
rect 43671 8072 43683 8075
rect 44085 8075 44143 8081
rect 44085 8072 44097 8075
rect 43671 8044 44097 8072
rect 43671 8041 43683 8044
rect 43625 8035 43683 8041
rect 44085 8041 44097 8044
rect 44131 8041 44143 8075
rect 44085 8035 44143 8041
rect 44453 8075 44511 8081
rect 44453 8041 44465 8075
rect 44499 8072 44511 8075
rect 45094 8072 45100 8084
rect 44499 8044 45100 8072
rect 44499 8041 44511 8044
rect 44453 8035 44511 8041
rect 45094 8032 45100 8044
rect 45152 8032 45158 8084
rect 45370 7896 45376 7948
rect 45428 7936 45434 7948
rect 45557 7939 45615 7945
rect 45557 7936 45569 7939
rect 45428 7908 45569 7936
rect 45428 7896 45434 7908
rect 45557 7905 45569 7908
rect 45603 7905 45615 7939
rect 45557 7899 45615 7905
rect 47581 7939 47639 7945
rect 47581 7905 47593 7939
rect 47627 7936 47639 7939
rect 47670 7936 47676 7948
rect 47627 7908 47676 7936
rect 47627 7905 47639 7908
rect 47581 7899 47639 7905
rect 47670 7896 47676 7908
rect 47728 7896 47734 7948
rect 43993 7871 44051 7877
rect 43993 7837 44005 7871
rect 44039 7868 44051 7871
rect 44818 7868 44824 7880
rect 44039 7840 44824 7868
rect 44039 7837 44051 7840
rect 43993 7831 44051 7837
rect 44818 7828 44824 7840
rect 44876 7828 44882 7880
rect 47302 7868 47308 7880
rect 47263 7840 47308 7868
rect 47302 7828 47308 7840
rect 47360 7828 47366 7880
rect 45186 7800 45192 7812
rect 45147 7772 45192 7800
rect 45186 7760 45192 7772
rect 45244 7760 45250 7812
rect 45278 7760 45284 7812
rect 45336 7800 45342 7812
rect 45336 7772 45381 7800
rect 45336 7760 45342 7772
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 32490 7732 32496 7744
rect 16908 7704 32496 7732
rect 16908 7692 16914 7704
rect 32490 7692 32496 7704
rect 32548 7692 32554 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 45186 7488 45192 7540
rect 45244 7528 45250 7540
rect 47949 7531 48007 7537
rect 47949 7528 47961 7531
rect 45244 7500 47961 7528
rect 45244 7488 45250 7500
rect 47949 7497 47961 7500
rect 47995 7497 48007 7531
rect 47949 7491 48007 7497
rect 44818 7460 44824 7472
rect 44779 7432 44824 7460
rect 44818 7420 44824 7432
rect 44876 7420 44882 7472
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 42886 7284 42892 7336
rect 42944 7324 42950 7336
rect 44729 7327 44787 7333
rect 44729 7324 44741 7327
rect 42944 7296 44741 7324
rect 42944 7284 42950 7296
rect 44729 7293 44741 7296
rect 44775 7293 44787 7327
rect 44729 7287 44787 7293
rect 45370 7284 45376 7336
rect 45428 7324 45434 7336
rect 45557 7327 45615 7333
rect 45557 7324 45569 7327
rect 45428 7296 45569 7324
rect 45428 7284 45434 7296
rect 45557 7293 45569 7296
rect 45603 7293 45615 7327
rect 45557 7287 45615 7293
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 43070 6400 43076 6452
rect 43128 6440 43134 6452
rect 48041 6443 48099 6449
rect 48041 6440 48053 6443
rect 43128 6412 48053 6440
rect 43128 6400 43134 6412
rect 48041 6409 48053 6412
rect 48087 6409 48099 6443
rect 48041 6403 48099 6409
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 32214 6236 32220 6248
rect 15620 6208 32220 6236
rect 15620 6196 15626 6208
rect 32214 6196 32220 6208
rect 32272 6196 32278 6248
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 28442 6168 28448 6180
rect 3292 6140 28448 6168
rect 3292 6128 3298 6140
rect 28442 6128 28448 6140
rect 28500 6128 28506 6180
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 40218 5692 40224 5704
rect 40179 5664 40224 5692
rect 40218 5652 40224 5664
rect 40276 5652 40282 5704
rect 42797 5695 42855 5701
rect 42797 5661 42809 5695
rect 42843 5692 42855 5695
rect 43530 5692 43536 5704
rect 42843 5664 43536 5692
rect 42843 5661 42855 5664
rect 42797 5655 42855 5661
rect 43530 5652 43536 5664
rect 43588 5652 43594 5704
rect 40310 5556 40316 5568
rect 40271 5528 40316 5556
rect 40310 5516 40316 5528
rect 40368 5516 40374 5568
rect 42610 5556 42616 5568
rect 42571 5528 42616 5556
rect 42610 5516 42616 5528
rect 42668 5516 42674 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 4028 5324 38608 5352
rect 4028 5312 4034 5324
rect 6638 5244 6644 5296
rect 6696 5284 6702 5296
rect 6696 5256 22094 5284
rect 6696 5244 6702 5256
rect 18690 5216 18696 5228
rect 18651 5188 18696 5216
rect 18690 5176 18696 5188
rect 18748 5176 18754 5228
rect 22066 5148 22094 5256
rect 36538 5244 36544 5296
rect 36596 5284 36602 5296
rect 37461 5287 37519 5293
rect 37461 5284 37473 5287
rect 36596 5256 37473 5284
rect 36596 5244 36602 5256
rect 37461 5253 37473 5256
rect 37507 5253 37519 5287
rect 37461 5247 37519 5253
rect 38381 5287 38439 5293
rect 38381 5253 38393 5287
rect 38427 5284 38439 5287
rect 38470 5284 38476 5296
rect 38427 5256 38476 5284
rect 38427 5253 38439 5256
rect 38381 5247 38439 5253
rect 38470 5244 38476 5256
rect 38528 5244 38534 5296
rect 38580 5284 38608 5324
rect 40218 5312 40224 5364
rect 40276 5352 40282 5364
rect 41049 5355 41107 5361
rect 41049 5352 41061 5355
rect 40276 5324 41061 5352
rect 40276 5312 40282 5324
rect 41049 5321 41061 5324
rect 41095 5321 41107 5355
rect 41049 5315 41107 5321
rect 42610 5284 42616 5296
rect 38580 5256 41414 5284
rect 42571 5256 42616 5284
rect 39669 5219 39727 5225
rect 39669 5185 39681 5219
rect 39715 5216 39727 5219
rect 40310 5216 40316 5228
rect 39715 5188 40316 5216
rect 39715 5185 39727 5188
rect 39669 5179 39727 5185
rect 40310 5176 40316 5188
rect 40368 5176 40374 5228
rect 40497 5219 40555 5225
rect 40497 5185 40509 5219
rect 40543 5216 40555 5219
rect 40770 5216 40776 5228
rect 40543 5188 40776 5216
rect 40543 5185 40555 5188
rect 40497 5179 40555 5185
rect 40770 5176 40776 5188
rect 40828 5176 40834 5228
rect 40954 5216 40960 5228
rect 40915 5188 40960 5216
rect 40954 5176 40960 5188
rect 41012 5176 41018 5228
rect 37369 5151 37427 5157
rect 37369 5148 37381 5151
rect 22066 5120 37381 5148
rect 37369 5117 37381 5120
rect 37415 5148 37427 5151
rect 38657 5151 38715 5157
rect 38657 5148 38669 5151
rect 37415 5120 38669 5148
rect 37415 5117 37427 5120
rect 37369 5111 37427 5117
rect 38657 5117 38669 5120
rect 38703 5117 38715 5151
rect 41386 5148 41414 5256
rect 42610 5244 42616 5256
rect 42668 5244 42674 5296
rect 43533 5287 43591 5293
rect 43533 5253 43545 5287
rect 43579 5284 43591 5287
rect 44358 5284 44364 5296
rect 43579 5256 44364 5284
rect 43579 5253 43591 5256
rect 43533 5247 43591 5253
rect 44358 5244 44364 5256
rect 44416 5244 44422 5296
rect 43809 5219 43867 5225
rect 43809 5216 43821 5219
rect 43364 5188 43821 5216
rect 42521 5151 42579 5157
rect 42521 5148 42533 5151
rect 41386 5120 42533 5148
rect 38657 5111 38715 5117
rect 42521 5117 42533 5120
rect 42567 5148 42579 5151
rect 43364 5148 43392 5188
rect 43809 5185 43821 5188
rect 43855 5185 43867 5219
rect 47854 5216 47860 5228
rect 47815 5188 47860 5216
rect 43809 5179 43867 5185
rect 47854 5176 47860 5188
rect 47912 5176 47918 5228
rect 42567 5120 43392 5148
rect 42567 5117 42579 5120
rect 42521 5111 42579 5117
rect 25590 5040 25596 5092
rect 25648 5080 25654 5092
rect 48041 5083 48099 5089
rect 48041 5080 48053 5083
rect 25648 5052 48053 5080
rect 25648 5040 25654 5052
rect 48041 5049 48053 5052
rect 48087 5049 48099 5083
rect 48041 5043 48099 5049
rect 18785 5015 18843 5021
rect 18785 4981 18797 5015
rect 18831 5012 18843 5015
rect 19242 5012 19248 5024
rect 18831 4984 19248 5012
rect 18831 4981 18843 4984
rect 18785 4975 18843 4981
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 39758 5012 39764 5024
rect 39719 4984 39764 5012
rect 39758 4972 39764 4984
rect 39816 4972 39822 5024
rect 40313 5015 40371 5021
rect 40313 4981 40325 5015
rect 40359 5012 40371 5015
rect 40494 5012 40500 5024
rect 40359 4984 40500 5012
rect 40359 4981 40371 4984
rect 40313 4975 40371 4981
rect 40494 4972 40500 4984
rect 40552 4972 40558 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 40218 4768 40224 4820
rect 40276 4808 40282 4820
rect 46566 4808 46572 4820
rect 40276 4780 46572 4808
rect 40276 4768 40282 4780
rect 46566 4768 46572 4780
rect 46624 4768 46630 4820
rect 18874 4700 18880 4752
rect 18932 4740 18938 4752
rect 18932 4712 25636 4740
rect 18932 4700 18938 4712
rect 25608 4684 25636 4712
rect 22186 4672 22192 4684
rect 21376 4644 22192 4672
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 18046 4604 18052 4616
rect 18007 4576 18052 4604
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 19334 4604 19340 4616
rect 19295 4576 19340 4604
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 19981 4607 20039 4613
rect 19981 4604 19993 4607
rect 19475 4576 19993 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 19981 4573 19993 4576
rect 20027 4573 20039 4607
rect 20622 4604 20628 4616
rect 20583 4576 20628 4604
rect 19981 4567 20039 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 21376 4613 21404 4644
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 25590 4672 25596 4684
rect 25503 4644 25596 4672
rect 25590 4632 25596 4644
rect 25648 4632 25654 4684
rect 27246 4672 27252 4684
rect 27207 4644 27252 4672
rect 27246 4632 27252 4644
rect 27304 4632 27310 4684
rect 39758 4632 39764 4684
rect 39816 4672 39822 4684
rect 40313 4675 40371 4681
rect 40313 4672 40325 4675
rect 39816 4644 40325 4672
rect 39816 4632 39822 4644
rect 40313 4641 40325 4644
rect 40359 4641 40371 4675
rect 40494 4672 40500 4684
rect 40455 4644 40500 4672
rect 40313 4635 40371 4641
rect 40494 4632 40500 4644
rect 40552 4632 40558 4684
rect 42150 4672 42156 4684
rect 42111 4644 42156 4672
rect 42150 4632 42156 4644
rect 42208 4632 42214 4684
rect 42886 4672 42892 4684
rect 42847 4644 42892 4672
rect 42886 4632 42892 4644
rect 42944 4632 42950 4684
rect 43901 4675 43959 4681
rect 43901 4641 43913 4675
rect 43947 4672 43959 4675
rect 44358 4672 44364 4684
rect 43947 4644 44364 4672
rect 43947 4641 43959 4644
rect 43901 4635 43959 4641
rect 44358 4632 44364 4644
rect 44416 4632 44422 4684
rect 44818 4632 44824 4684
rect 44876 4672 44882 4684
rect 47581 4675 47639 4681
rect 47581 4672 47593 4675
rect 44876 4644 47593 4672
rect 44876 4632 44882 4644
rect 47581 4641 47593 4644
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 21361 4607 21419 4613
rect 21361 4573 21373 4607
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 22554 4604 22560 4616
rect 22051 4576 22560 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 22649 4607 22707 4613
rect 22649 4573 22661 4607
rect 22695 4604 22707 4607
rect 23750 4604 23756 4616
rect 22695 4576 23756 4604
rect 22695 4573 22707 4576
rect 22649 4567 22707 4573
rect 23750 4564 23756 4576
rect 23808 4564 23814 4616
rect 25409 4607 25467 4613
rect 25409 4573 25421 4607
rect 25455 4573 25467 4607
rect 46658 4604 46664 4616
rect 46619 4576 46664 4604
rect 25409 4567 25467 4573
rect 21453 4539 21511 4545
rect 21453 4505 21465 4539
rect 21499 4536 21511 4539
rect 22462 4536 22468 4548
rect 21499 4508 22468 4536
rect 21499 4505 21511 4508
rect 21453 4499 21511 4505
rect 22462 4496 22468 4508
rect 22520 4496 22526 4548
rect 18138 4468 18144 4480
rect 18099 4440 18144 4468
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 20073 4471 20131 4477
rect 20073 4437 20085 4471
rect 20119 4468 20131 4471
rect 20346 4468 20352 4480
rect 20119 4440 20352 4468
rect 20119 4437 20131 4440
rect 20073 4431 20131 4437
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 20717 4471 20775 4477
rect 20717 4437 20729 4471
rect 20763 4468 20775 4471
rect 20990 4468 20996 4480
rect 20763 4440 20996 4468
rect 20763 4437 20775 4440
rect 20717 4431 20775 4437
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 22097 4471 22155 4477
rect 22097 4437 22109 4471
rect 22143 4468 22155 4471
rect 22278 4468 22284 4480
rect 22143 4440 22284 4468
rect 22143 4437 22155 4440
rect 22097 4431 22155 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 22738 4468 22744 4480
rect 22699 4440 22744 4468
rect 22738 4428 22744 4440
rect 22796 4428 22802 4480
rect 25314 4428 25320 4480
rect 25372 4468 25378 4480
rect 25424 4468 25452 4567
rect 46658 4564 46664 4576
rect 46716 4564 46722 4616
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47305 4607 47363 4613
rect 47305 4604 47317 4607
rect 46900 4576 47317 4604
rect 46900 4564 46906 4576
rect 47305 4573 47317 4576
rect 47351 4573 47363 4607
rect 47305 4567 47363 4573
rect 39482 4496 39488 4548
rect 39540 4536 39546 4548
rect 42886 4536 42892 4548
rect 39540 4508 42892 4536
rect 39540 4496 39546 4508
rect 42886 4496 42892 4508
rect 42944 4496 42950 4548
rect 42981 4539 43039 4545
rect 42981 4505 42993 4539
rect 43027 4536 43039 4539
rect 43070 4536 43076 4548
rect 43027 4508 43076 4536
rect 43027 4505 43039 4508
rect 42981 4499 43039 4505
rect 43070 4496 43076 4508
rect 43128 4496 43134 4548
rect 32122 4468 32128 4480
rect 25372 4440 32128 4468
rect 25372 4428 25378 4440
rect 32122 4428 32128 4440
rect 32180 4428 32186 4480
rect 46474 4428 46480 4480
rect 46532 4468 46538 4480
rect 46753 4471 46811 4477
rect 46753 4468 46765 4471
rect 46532 4440 46765 4468
rect 46532 4428 46538 4440
rect 46753 4437 46765 4440
rect 46799 4437 46811 4471
rect 46753 4431 46811 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19797 4267 19855 4273
rect 19797 4264 19809 4267
rect 19392 4236 19809 4264
rect 19392 4224 19398 4236
rect 19797 4233 19809 4236
rect 19843 4233 19855 4267
rect 19797 4227 19855 4233
rect 20441 4267 20499 4273
rect 20441 4233 20453 4267
rect 20487 4264 20499 4267
rect 20622 4264 20628 4276
rect 20487 4236 20628 4264
rect 20487 4233 20499 4236
rect 20441 4227 20499 4233
rect 20622 4224 20628 4236
rect 20680 4224 20686 4276
rect 38378 4264 38384 4276
rect 37476 4236 38384 4264
rect 37476 4205 37504 4236
rect 38378 4224 38384 4236
rect 38436 4224 38442 4276
rect 39684 4236 40724 4264
rect 37461 4199 37519 4205
rect 37461 4196 37473 4199
rect 17696 4168 18000 4196
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 13722 4128 13728 4140
rect 13683 4100 13728 4128
rect 10137 4091 10195 4097
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 2958 4060 2964 4072
rect 2271 4032 2964 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2056 3992 2084 4023
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 7374 4060 7380 4072
rect 3108 4032 3153 4060
rect 7335 4032 7380 4060
rect 3108 4020 3114 4032
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7558 4060 7564 4072
rect 7519 4032 7564 4060
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4029 7895 4063
rect 10152 4060 10180 4091
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17221 4131 17279 4137
rect 17221 4128 17233 4131
rect 17092 4100 17233 4128
rect 17092 4088 17098 4100
rect 17221 4097 17233 4100
rect 17267 4097 17279 4131
rect 17221 4091 17279 4097
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17696 4128 17724 4168
rect 17552 4100 17724 4128
rect 17552 4088 17558 4100
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 17828 4100 17877 4128
rect 17828 4088 17834 4100
rect 17865 4097 17877 4100
rect 17911 4097 17923 4131
rect 17972 4128 18000 4168
rect 28966 4168 36492 4196
rect 19061 4131 19119 4137
rect 17972 4100 19012 4128
rect 17865 4091 17923 4097
rect 16022 4060 16028 4072
rect 10152 4032 16028 4060
rect 7837 4023 7895 4029
rect 3970 3992 3976 4004
rect 2056 3964 3976 3992
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 7852 3992 7880 4023
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4060 17371 4063
rect 18690 4060 18696 4072
rect 17359 4032 18696 4060
rect 17359 4029 17371 4032
rect 17313 4023 17371 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 18984 4060 19012 4100
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 19334 4128 19340 4140
rect 19107 4100 19340 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19702 4128 19708 4140
rect 19663 4100 19708 4128
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 20346 4128 20352 4140
rect 20307 4100 20352 4128
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20990 4128 20996 4140
rect 20951 4100 20996 4128
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 21542 4088 21548 4140
rect 21600 4128 21606 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21600 4100 21833 4128
rect 21600 4088 21606 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 22462 4128 22468 4140
rect 22423 4100 22468 4128
rect 21821 4091 21879 4097
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 23109 4131 23167 4137
rect 22612 4100 22657 4128
rect 22612 4088 22618 4100
rect 23109 4097 23121 4131
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 23753 4131 23811 4137
rect 23753 4097 23765 4131
rect 23799 4097 23811 4131
rect 23753 4091 23811 4097
rect 20530 4060 20536 4072
rect 18984 4032 20536 4060
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 23124 4060 23152 4091
rect 20772 4032 23152 4060
rect 20772 4020 20778 4032
rect 7156 3964 7880 3992
rect 7156 3952 7162 3964
rect 12066 3952 12072 4004
rect 12124 3992 12130 4004
rect 18598 3992 18604 4004
rect 12124 3964 18604 3992
rect 12124 3952 12130 3964
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 18782 3952 18788 4004
rect 18840 3992 18846 4004
rect 23201 3995 23259 4001
rect 23201 3992 23213 3995
rect 18840 3964 23213 3992
rect 18840 3952 18846 3964
rect 23201 3961 23213 3964
rect 23247 3961 23259 3995
rect 23768 3992 23796 4091
rect 26694 4088 26700 4140
rect 26752 4128 26758 4140
rect 27338 4128 27344 4140
rect 26752 4100 27344 4128
rect 26752 4088 26758 4100
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 28966 3992 28994 4168
rect 31662 4088 31668 4140
rect 31720 4128 31726 4140
rect 31720 4100 32168 4128
rect 31720 4088 31726 4100
rect 32140 4060 32168 4100
rect 36464 4060 36492 4168
rect 37292 4168 37473 4196
rect 36630 4088 36636 4140
rect 36688 4132 36694 4140
rect 36725 4132 36783 4137
rect 36688 4131 36783 4132
rect 36688 4104 36737 4131
rect 36688 4088 36694 4104
rect 36725 4097 36737 4104
rect 36771 4097 36783 4131
rect 36725 4091 36783 4097
rect 36906 4088 36912 4140
rect 36964 4128 36970 4140
rect 37292 4128 37320 4168
rect 37461 4165 37473 4168
rect 37507 4165 37519 4199
rect 37461 4159 37519 4165
rect 37553 4199 37611 4205
rect 37553 4165 37565 4199
rect 37599 4196 37611 4199
rect 37642 4196 37648 4208
rect 37599 4168 37648 4196
rect 37599 4165 37611 4168
rect 37553 4159 37611 4165
rect 37642 4156 37648 4168
rect 37700 4156 37706 4208
rect 38470 4196 38476 4208
rect 38431 4168 38476 4196
rect 38470 4156 38476 4168
rect 38528 4156 38534 4208
rect 39684 4196 39712 4236
rect 40586 4196 40592 4208
rect 39592 4168 39712 4196
rect 40547 4168 40592 4196
rect 39592 4128 39620 4168
rect 40586 4156 40592 4168
rect 40644 4156 40650 4208
rect 40696 4196 40724 4236
rect 40770 4224 40776 4276
rect 40828 4264 40834 4276
rect 40957 4267 41015 4273
rect 40957 4264 40969 4267
rect 40828 4236 40969 4264
rect 40828 4224 40834 4236
rect 40957 4233 40969 4236
rect 41003 4233 41015 4267
rect 40957 4227 41015 4233
rect 41230 4196 41236 4208
rect 40696 4168 41236 4196
rect 41230 4156 41236 4168
rect 41288 4156 41294 4208
rect 47762 4196 47768 4208
rect 47723 4168 47768 4196
rect 47762 4156 47768 4168
rect 47820 4156 47826 4208
rect 40773 4131 40831 4137
rect 40773 4128 40785 4131
rect 36964 4100 37320 4128
rect 38304 4100 39620 4128
rect 39684 4100 40785 4128
rect 36964 4088 36970 4100
rect 38304 4060 38332 4100
rect 39684 4072 39712 4100
rect 40773 4097 40785 4100
rect 40819 4097 40831 4131
rect 40773 4091 40831 4097
rect 40862 4088 40868 4140
rect 40920 4128 40926 4140
rect 42981 4131 43039 4137
rect 42981 4128 42993 4131
rect 40920 4100 42993 4128
rect 40920 4088 40926 4100
rect 42981 4097 42993 4100
rect 43027 4097 43039 4131
rect 46750 4128 46756 4140
rect 46711 4100 46756 4128
rect 42981 4091 43039 4097
rect 46750 4088 46756 4100
rect 46808 4088 46814 4140
rect 32140 4032 36400 4060
rect 36464 4032 38332 4060
rect 23768 3964 28994 3992
rect 23201 3955 23259 3961
rect 32122 3952 32128 4004
rect 32180 3992 32186 4004
rect 36170 3992 36176 4004
rect 32180 3964 36176 3992
rect 32180 3952 32186 3964
rect 36170 3952 36176 3964
rect 36228 3952 36234 4004
rect 10226 3924 10232 3936
rect 10187 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11572 3896 11713 3924
rect 11572 3884 11578 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 13998 3924 14004 3936
rect 13863 3896 14004 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 17954 3924 17960 3936
rect 17915 3896 17960 3924
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 19153 3927 19211 3933
rect 19153 3924 19165 3927
rect 18564 3896 19165 3924
rect 18564 3884 18570 3896
rect 19153 3893 19165 3896
rect 19199 3893 19211 3927
rect 19153 3887 19211 3893
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20864 3896 21097 3924
rect 20864 3884 20870 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 21913 3927 21971 3933
rect 21913 3893 21925 3927
rect 21959 3924 21971 3927
rect 22094 3924 22100 3936
rect 21959 3896 22100 3924
rect 21959 3893 21971 3896
rect 21913 3887 21971 3893
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 23106 3884 23112 3936
rect 23164 3924 23170 3936
rect 23845 3927 23903 3933
rect 23845 3924 23857 3927
rect 23164 3896 23857 3924
rect 23164 3884 23170 3896
rect 23845 3893 23857 3896
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 26234 3884 26240 3936
rect 26292 3924 26298 3936
rect 27522 3924 27528 3936
rect 26292 3896 27528 3924
rect 26292 3884 26298 3896
rect 27522 3884 27528 3896
rect 27580 3884 27586 3936
rect 32766 3884 32772 3936
rect 32824 3924 32830 3936
rect 36262 3924 36268 3936
rect 32824 3896 36268 3924
rect 32824 3884 32830 3896
rect 36262 3884 36268 3896
rect 36320 3884 36326 3936
rect 36372 3924 36400 4032
rect 38378 4020 38384 4072
rect 38436 4060 38442 4072
rect 39482 4060 39488 4072
rect 38436 4032 39488 4060
rect 38436 4020 38442 4032
rect 39482 4020 39488 4032
rect 39540 4020 39546 4072
rect 39666 4060 39672 4072
rect 39627 4032 39672 4060
rect 39666 4020 39672 4032
rect 39724 4020 39730 4072
rect 39942 4020 39948 4072
rect 40000 4060 40006 4072
rect 47210 4060 47216 4072
rect 40000 4032 47216 4060
rect 40000 4020 40006 4032
rect 47210 4020 47216 4032
rect 47268 4020 47274 4072
rect 36538 3992 36544 4004
rect 36499 3964 36544 3992
rect 36538 3952 36544 3964
rect 36596 3952 36602 4004
rect 47949 3995 48007 4001
rect 47949 3992 47961 3995
rect 37476 3964 47961 3992
rect 37476 3924 37504 3964
rect 47949 3961 47961 3964
rect 47995 3961 48007 3995
rect 47949 3955 48007 3961
rect 40126 3924 40132 3936
rect 36372 3896 37504 3924
rect 40087 3896 40132 3924
rect 40126 3884 40132 3896
rect 40184 3884 40190 3936
rect 40402 3884 40408 3936
rect 40460 3924 40466 3936
rect 42794 3924 42800 3936
rect 40460 3896 42800 3924
rect 40460 3884 40466 3896
rect 42794 3884 42800 3896
rect 42852 3884 42858 3936
rect 42978 3884 42984 3936
rect 43036 3924 43042 3936
rect 43073 3927 43131 3933
rect 43073 3924 43085 3927
rect 43036 3896 43085 3924
rect 43036 3884 43042 3896
rect 43073 3893 43085 3896
rect 43119 3893 43131 3927
rect 43806 3924 43812 3936
rect 43767 3896 43812 3924
rect 43073 3887 43131 3893
rect 43806 3884 43812 3896
rect 43864 3884 43870 3936
rect 46290 3924 46296 3936
rect 46251 3896 46296 3924
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 46934 3924 46940 3936
rect 46895 3896 46940 3924
rect 46934 3884 46940 3896
rect 46992 3884 46998 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 2958 3720 2964 3732
rect 2919 3692 2964 3720
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3970 3720 3976 3732
rect 3931 3692 3976 3720
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 17034 3720 17040 3732
rect 16995 3692 17040 3720
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 19702 3720 19708 3732
rect 18647 3692 19708 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 19702 3680 19708 3692
rect 19760 3680 19766 3732
rect 20254 3680 20260 3732
rect 20312 3680 20318 3732
rect 21542 3720 21548 3732
rect 21503 3692 21548 3720
rect 21542 3680 21548 3692
rect 21600 3680 21606 3732
rect 22186 3720 22192 3732
rect 22147 3692 22192 3720
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 23658 3680 23664 3732
rect 23716 3720 23722 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 23716 3692 23765 3720
rect 23716 3680 23722 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 23753 3683 23811 3689
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 25188 3692 27292 3720
rect 25188 3680 25194 3692
rect 5276 3624 11744 3652
rect 5276 3584 5304 3624
rect 6454 3584 6460 3596
rect 2884 3556 5304 3584
rect 6415 3556 6460 3584
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1762 3516 1768 3528
rect 1719 3488 1768 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 2130 3516 2136 3528
rect 2091 3488 2136 3516
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2884 3525 2912 3556
rect 5276 3525 5304 3556
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 9309 3587 9367 3593
rect 9309 3553 9321 3587
rect 9355 3584 9367 3587
rect 9490 3584 9496 3596
rect 9355 3556 9496 3584
rect 9355 3553 9367 3556
rect 9309 3547 9367 3553
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9640 3556 9781 3584
rect 9640 3544 9646 3556
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 11716 3584 11744 3624
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 18414 3652 18420 3664
rect 13780 3624 18420 3652
rect 13780 3612 13786 3624
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 20272 3652 20300 3680
rect 18748 3624 20300 3652
rect 27264 3652 27292 3692
rect 27338 3680 27344 3732
rect 27396 3720 27402 3732
rect 32674 3720 32680 3732
rect 27396 3692 32680 3720
rect 27396 3680 27402 3692
rect 32674 3680 32680 3692
rect 32732 3680 32738 3732
rect 32766 3680 32772 3732
rect 32824 3720 32830 3732
rect 40221 3723 40279 3729
rect 32824 3692 39436 3720
rect 32824 3680 32830 3692
rect 39298 3652 39304 3664
rect 27264 3624 39304 3652
rect 18748 3612 18754 3624
rect 39298 3612 39304 3624
rect 39356 3612 39362 3664
rect 39408 3652 39436 3692
rect 40221 3689 40233 3723
rect 40267 3720 40279 3723
rect 40954 3720 40960 3732
rect 40267 3692 40960 3720
rect 40267 3689 40279 3692
rect 40221 3683 40279 3689
rect 40954 3680 40960 3692
rect 41012 3680 41018 3732
rect 41414 3680 41420 3732
rect 41472 3720 41478 3732
rect 43165 3723 43223 3729
rect 43165 3720 43177 3723
rect 41472 3692 43177 3720
rect 41472 3680 41478 3692
rect 43165 3689 43177 3692
rect 43211 3689 43223 3723
rect 43530 3720 43536 3732
rect 43491 3692 43536 3720
rect 43165 3683 43223 3689
rect 43530 3680 43536 3692
rect 43588 3680 43594 3732
rect 40402 3652 40408 3664
rect 39408 3624 40408 3652
rect 40402 3612 40408 3624
rect 40460 3612 40466 3664
rect 40494 3612 40500 3664
rect 40552 3652 40558 3664
rect 46934 3652 46940 3664
rect 40552 3624 46940 3652
rect 40552 3612 40558 3624
rect 46934 3612 46940 3624
rect 46992 3612 46998 3664
rect 26602 3584 26608 3596
rect 11716 3556 26608 3584
rect 9769 3547 9827 3553
rect 26602 3544 26608 3556
rect 26660 3544 26666 3596
rect 26878 3544 26884 3596
rect 26936 3584 26942 3596
rect 33686 3584 33692 3596
rect 26936 3556 33692 3584
rect 26936 3544 26942 3556
rect 33686 3544 33692 3556
rect 33744 3544 33750 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 40218 3584 40224 3596
rect 33928 3556 40224 3584
rect 33928 3544 33934 3556
rect 40218 3544 40224 3556
rect 40276 3544 40282 3596
rect 42150 3584 42156 3596
rect 42111 3556 42156 3584
rect 42150 3544 42156 3556
rect 42208 3544 42214 3596
rect 46290 3584 46296 3596
rect 44560 3556 45692 3584
rect 46251 3556 46296 3584
rect 44560 3528 44588 3556
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5902 3516 5908 3528
rect 5863 3488 5908 3516
rect 5261 3479 5319 3485
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 8202 3516 8208 3528
rect 8163 3488 8208 3516
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 12066 3516 12072 3528
rect 12027 3488 12072 3516
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13872 3488 14289 3516
rect 13872 3476 13878 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 6089 3451 6147 3457
rect 6089 3448 6101 3451
rect 5399 3420 6101 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 6089 3417 6101 3420
rect 6135 3417 6147 3451
rect 6089 3411 6147 3417
rect 9493 3451 9551 3457
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 10226 3448 10232 3460
rect 9539 3420 10232 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 10226 3408 10232 3420
rect 10284 3408 10290 3460
rect 16960 3448 16988 3479
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17276 3488 17601 3516
rect 17276 3476 17282 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 18506 3516 18512 3528
rect 18467 3488 18512 3516
rect 17589 3479 17647 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 18656 3488 19533 3516
rect 18656 3476 18662 3488
rect 19521 3485 19533 3488
rect 19567 3516 19579 3519
rect 20346 3516 20352 3528
rect 19567 3488 19840 3516
rect 20307 3488 20352 3516
rect 19567 3485 19579 3488
rect 19521 3479 19579 3485
rect 18230 3448 18236 3460
rect 16960 3420 18236 3448
rect 18230 3408 18236 3420
rect 18288 3408 18294 3460
rect 18874 3408 18880 3460
rect 18932 3448 18938 3460
rect 19702 3448 19708 3460
rect 18932 3420 19708 3448
rect 18932 3408 18938 3420
rect 19702 3408 19708 3420
rect 19760 3408 19766 3460
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2004 3352 2237 3380
rect 2004 3340 2010 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 8260 3352 8309 3380
rect 8260 3340 8266 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8297 3343 8355 3349
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12161 3383 12219 3389
rect 12161 3380 12173 3383
rect 11756 3352 12173 3380
rect 11756 3340 11762 3352
rect 12161 3349 12173 3352
rect 12207 3349 12219 3383
rect 17678 3380 17684 3392
rect 17639 3352 17684 3380
rect 12161 3343 12219 3349
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 19484 3352 19625 3380
rect 19484 3340 19490 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19812 3380 19840 3488
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 20806 3516 20812 3528
rect 20767 3488 20812 3516
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3516 20959 3519
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 20947 3488 21465 3516
rect 20947 3485 20959 3488
rect 20901 3479 20959 3485
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 22152 3488 22197 3516
rect 22152 3476 22158 3488
rect 22922 3476 22928 3528
rect 22980 3516 22986 3528
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 22980 3488 23213 3516
rect 22980 3476 22986 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 23661 3519 23719 3525
rect 23661 3485 23673 3519
rect 23707 3485 23719 3519
rect 25406 3516 25412 3528
rect 25367 3488 25412 3516
rect 23661 3479 23719 3485
rect 19886 3408 19892 3460
rect 19944 3448 19950 3460
rect 23676 3448 23704 3479
rect 25406 3476 25412 3488
rect 25464 3476 25470 3528
rect 27246 3516 27252 3528
rect 27207 3488 27252 3516
rect 27246 3476 27252 3488
rect 27304 3476 27310 3528
rect 32674 3476 32680 3528
rect 32732 3516 32738 3528
rect 32950 3516 32956 3528
rect 32732 3488 32956 3516
rect 32732 3476 32738 3488
rect 32950 3476 32956 3488
rect 33008 3476 33014 3528
rect 33134 3476 33140 3528
rect 33192 3516 33198 3528
rect 33781 3519 33839 3525
rect 33781 3516 33793 3519
rect 33192 3488 33793 3516
rect 33192 3476 33198 3488
rect 33781 3485 33793 3488
rect 33827 3485 33839 3519
rect 33781 3479 33839 3485
rect 37826 3476 37832 3528
rect 37884 3516 37890 3528
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 37884 3488 38117 3516
rect 37884 3476 37890 3488
rect 38105 3485 38117 3488
rect 38151 3485 38163 3519
rect 38105 3479 38163 3485
rect 38657 3519 38715 3525
rect 38657 3485 38669 3519
rect 38703 3516 38715 3519
rect 39942 3516 39948 3528
rect 38703 3488 39948 3516
rect 38703 3485 38715 3488
rect 38657 3479 38715 3485
rect 39942 3476 39948 3488
rect 40000 3476 40006 3528
rect 40126 3476 40132 3528
rect 40184 3516 40190 3528
rect 40770 3516 40776 3528
rect 40184 3488 40229 3516
rect 40731 3488 40776 3516
rect 40184 3476 40190 3488
rect 40770 3476 40776 3488
rect 40828 3476 40834 3528
rect 43070 3516 43076 3528
rect 43031 3488 43076 3516
rect 43070 3476 43076 3488
rect 43128 3476 43134 3528
rect 43993 3519 44051 3525
rect 43993 3485 44005 3519
rect 44039 3516 44051 3519
rect 44542 3516 44548 3528
rect 44039 3488 44548 3516
rect 44039 3485 44051 3488
rect 43993 3479 44051 3485
rect 44542 3476 44548 3488
rect 44600 3476 44606 3528
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45664 3525 45692 3556
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 19944 3420 23704 3448
rect 25593 3451 25651 3457
rect 19944 3408 19950 3420
rect 25593 3417 25605 3451
rect 25639 3448 25651 3451
rect 26970 3448 26976 3460
rect 25639 3420 26976 3448
rect 25639 3417 25651 3420
rect 25593 3411 25651 3417
rect 26970 3408 26976 3420
rect 27028 3408 27034 3460
rect 33042 3448 33048 3460
rect 33003 3420 33048 3448
rect 33042 3408 33048 3420
rect 33100 3408 33106 3460
rect 33870 3408 33876 3460
rect 33928 3448 33934 3460
rect 40957 3451 41015 3457
rect 33928 3420 40908 3448
rect 33928 3408 33934 3420
rect 40880 3392 40908 3420
rect 40957 3417 40969 3451
rect 41003 3448 41015 3451
rect 41322 3448 41328 3460
rect 41003 3420 41328 3448
rect 41003 3417 41015 3420
rect 40957 3411 41015 3417
rect 41322 3408 41328 3420
rect 41380 3408 41386 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 26234 3380 26240 3392
rect 19812 3352 26240 3380
rect 19613 3343 19671 3349
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 26326 3340 26332 3392
rect 26384 3380 26390 3392
rect 36538 3380 36544 3392
rect 26384 3352 36544 3380
rect 26384 3340 26390 3352
rect 36538 3340 36544 3352
rect 36596 3340 36602 3392
rect 38010 3340 38016 3392
rect 38068 3380 38074 3392
rect 38749 3383 38807 3389
rect 38749 3380 38761 3383
rect 38068 3352 38761 3380
rect 38068 3340 38074 3352
rect 38749 3349 38761 3352
rect 38795 3349 38807 3383
rect 38749 3343 38807 3349
rect 40862 3340 40868 3392
rect 40920 3340 40926 3392
rect 44082 3380 44088 3392
rect 44043 3352 44088 3380
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 3936 3148 36216 3176
rect 3936 3136 3942 3148
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 8202 3108 8208 3120
rect 8163 3080 8208 3108
rect 8202 3068 8208 3080
rect 8260 3068 8266 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 13998 3108 14004 3120
rect 13959 3080 14004 3108
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 17770 3108 17776 3120
rect 17731 3080 17776 3108
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 18874 3108 18880 3120
rect 18835 3080 18880 3108
rect 18874 3068 18880 3080
rect 18932 3068 18938 3120
rect 32766 3108 32772 3120
rect 19444 3080 32772 3108
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 5960 3012 6561 3040
rect 5960 3000 5966 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7374 3000 7380 3052
rect 7432 3040 7438 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7432 3012 7573 3040
rect 7432 3000 7438 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 7561 3003 7619 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 17494 3040 17500 3052
rect 16899 3012 17500 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 17678 3040 17684 3052
rect 17639 3012 17684 3040
rect 17678 3000 17684 3012
rect 17736 3000 17742 3052
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19444 3040 19472 3080
rect 32766 3068 32772 3080
rect 32824 3068 32830 3120
rect 33042 3108 33048 3120
rect 33003 3080 33048 3108
rect 33042 3068 33048 3080
rect 33100 3068 33106 3120
rect 18892 3012 19472 3040
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 8018 2972 8024 2984
rect 7979 2944 8024 2972
rect 2225 2935 2283 2941
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 8496 2904 8524 2935
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11020 2944 11989 2972
rect 11020 2932 11026 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 15252 2944 16773 2972
rect 15252 2932 15258 2944
rect 16761 2941 16773 2944
rect 16807 2941 16819 2975
rect 17218 2972 17224 2984
rect 17179 2944 17224 2972
rect 16761 2935 16819 2941
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 18892 2972 18920 3012
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 22281 3043 22339 3049
rect 22281 3040 22293 3043
rect 21968 3012 22293 3040
rect 21968 3000 21974 3012
rect 22281 3009 22293 3012
rect 22327 3009 22339 3043
rect 22922 3040 22928 3052
rect 22883 3012 22928 3040
rect 22281 3003 22339 3009
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 25590 3040 25596 3052
rect 25551 3012 25596 3040
rect 25590 3000 25596 3012
rect 25648 3000 25654 3052
rect 26050 3000 26056 3052
rect 26108 3040 26114 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26108 3012 27169 3040
rect 26108 3000 26114 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 17460 2944 18920 2972
rect 19429 2975 19487 2981
rect 17460 2932 17466 2944
rect 19429 2941 19441 2975
rect 19475 2956 19487 2975
rect 19475 2941 19564 2956
rect 19429 2935 19564 2941
rect 19444 2928 19564 2935
rect 19610 2932 19616 2984
rect 19668 2972 19674 2984
rect 19978 2972 19984 2984
rect 19668 2944 19713 2972
rect 19939 2944 19984 2972
rect 19668 2932 19674 2944
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 23106 2972 23112 2984
rect 23067 2944 23112 2972
rect 23106 2932 23112 2944
rect 23164 2932 23170 2984
rect 23385 2975 23443 2981
rect 23385 2941 23397 2975
rect 23431 2941 23443 2975
rect 32861 2975 32919 2981
rect 23385 2935 23443 2941
rect 25792 2944 31754 2972
rect 19536 2904 19564 2928
rect 20346 2904 20352 2916
rect 7800 2876 8524 2904
rect 8956 2876 19012 2904
rect 19536 2876 20352 2904
rect 7800 2864 7806 2876
rect 7558 2796 7564 2848
rect 7616 2836 7622 2848
rect 8956 2836 8984 2876
rect 7616 2808 8984 2836
rect 7616 2796 7622 2808
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9582 2836 9588 2848
rect 9088 2808 9588 2836
rect 9088 2796 9094 2808
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 18984 2836 19012 2876
rect 20346 2864 20352 2876
rect 20404 2864 20410 2916
rect 22462 2904 22468 2916
rect 22423 2876 22468 2904
rect 22462 2864 22468 2876
rect 22520 2864 22526 2916
rect 22554 2864 22560 2916
rect 22612 2904 22618 2916
rect 23400 2904 23428 2935
rect 22612 2876 23428 2904
rect 22612 2864 22618 2876
rect 25792 2836 25820 2944
rect 31726 2904 31754 2944
rect 32861 2941 32873 2975
rect 32907 2972 32919 2975
rect 33134 2972 33140 2984
rect 32907 2944 33140 2972
rect 32907 2941 32919 2944
rect 32861 2935 32919 2941
rect 33134 2932 33140 2944
rect 33192 2932 33198 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 36188 2972 36216 3148
rect 36630 3136 36636 3188
rect 36688 3176 36694 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 36688 3148 36737 3176
rect 36688 3136 36694 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 37642 3176 37648 3188
rect 36725 3139 36783 3145
rect 36832 3148 37648 3176
rect 36832 3108 36860 3148
rect 37642 3136 37648 3148
rect 37700 3176 37706 3188
rect 37700 3148 38424 3176
rect 37700 3136 37706 3148
rect 38010 3108 38016 3120
rect 36280 3080 36860 3108
rect 37971 3080 38016 3108
rect 36280 3049 36308 3080
rect 38010 3068 38016 3080
rect 38068 3068 38074 3120
rect 38396 3108 38424 3148
rect 40770 3136 40776 3188
rect 40828 3176 40834 3188
rect 40865 3179 40923 3185
rect 40865 3176 40877 3179
rect 40828 3148 40877 3176
rect 40828 3136 40834 3148
rect 40865 3145 40877 3148
rect 40911 3145 40923 3179
rect 41322 3176 41328 3188
rect 41283 3148 41328 3176
rect 40865 3139 40923 3145
rect 41322 3136 41328 3148
rect 41380 3136 41386 3188
rect 43806 3176 43812 3188
rect 42812 3148 43812 3176
rect 41598 3108 41604 3120
rect 38396 3080 41604 3108
rect 41598 3068 41604 3080
rect 41656 3068 41662 3120
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3009 36323 3043
rect 37826 3040 37832 3052
rect 37787 3012 37832 3040
rect 36265 3003 36323 3009
rect 37826 3000 37832 3012
rect 37884 3000 37890 3052
rect 39224 3012 41414 3040
rect 39224 2972 39252 3012
rect 36188 2944 39252 2972
rect 39298 2932 39304 2984
rect 39356 2972 39362 2984
rect 39356 2944 39401 2972
rect 39356 2932 39362 2944
rect 39482 2932 39488 2984
rect 39540 2972 39546 2984
rect 40221 2975 40279 2981
rect 40221 2972 40233 2975
rect 39540 2944 40233 2972
rect 39540 2932 39546 2944
rect 40221 2941 40233 2944
rect 40267 2941 40279 2975
rect 40402 2972 40408 2984
rect 40363 2944 40408 2972
rect 40221 2935 40279 2941
rect 40402 2932 40408 2944
rect 40460 2932 40466 2984
rect 41386 2972 41414 3012
rect 41506 3000 41512 3052
rect 41564 3040 41570 3052
rect 42812 3049 42840 3148
rect 43806 3136 43812 3148
rect 43864 3136 43870 3188
rect 48038 3176 48044 3188
rect 47999 3148 48044 3176
rect 48038 3136 48044 3148
rect 48096 3136 48102 3188
rect 42978 3108 42984 3120
rect 42939 3080 42984 3108
rect 42978 3068 42984 3080
rect 43036 3068 43042 3120
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 42797 3043 42855 3049
rect 41564 3012 41609 3040
rect 41564 3000 41570 3012
rect 42797 3009 42809 3043
rect 42843 3009 42855 3043
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 42797 3003 42855 3009
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3040 47823 3043
rect 48314 3040 48320 3052
rect 47811 3012 48320 3040
rect 47811 3009 47823 3012
rect 47765 3003 47823 3009
rect 48314 3000 48320 3012
rect 48372 3000 48378 3052
rect 41874 2972 41880 2984
rect 41386 2944 41880 2972
rect 41874 2932 41880 2944
rect 41932 2932 41938 2984
rect 43162 2932 43168 2984
rect 43220 2972 43226 2984
rect 43257 2975 43315 2981
rect 43257 2972 43269 2975
rect 43220 2944 43269 2972
rect 43220 2932 43226 2944
rect 43257 2941 43269 2944
rect 43303 2941 43315 2975
rect 43257 2935 43315 2941
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 44082 2904 44088 2916
rect 25884 2876 27108 2904
rect 31726 2876 44088 2904
rect 25884 2845 25912 2876
rect 18984 2808 25820 2836
rect 25869 2839 25927 2845
rect 25869 2805 25881 2839
rect 25915 2805 25927 2839
rect 26050 2836 26056 2848
rect 26011 2808 26056 2836
rect 25869 2799 25927 2805
rect 26050 2796 26056 2808
rect 26108 2796 26114 2848
rect 26970 2836 26976 2848
rect 26931 2808 26976 2836
rect 26970 2796 26976 2808
rect 27028 2796 27034 2848
rect 27080 2836 27108 2876
rect 44082 2864 44088 2876
rect 44140 2864 44146 2916
rect 35526 2836 35532 2848
rect 27080 2808 35532 2836
rect 35526 2796 35532 2808
rect 35584 2796 35590 2848
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 36357 2839 36415 2845
rect 36357 2836 36369 2839
rect 36228 2808 36369 2836
rect 36228 2796 36234 2808
rect 36357 2805 36369 2808
rect 36403 2805 36415 2839
rect 36357 2799 36415 2805
rect 36538 2796 36544 2848
rect 36596 2836 36602 2848
rect 47578 2836 47584 2848
rect 36596 2808 47584 2836
rect 36596 2796 36602 2808
rect 47578 2796 47584 2808
rect 47636 2796 47642 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 3234 2632 3240 2644
rect 3099 2604 3240 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 8018 2592 8024 2644
rect 8076 2632 8082 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 8076 2604 8217 2632
rect 8076 2592 8082 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 16850 2632 16856 2644
rect 8205 2595 8263 2601
rect 11716 2604 16712 2632
rect 16811 2604 16856 2632
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 11716 2564 11744 2604
rect 16684 2564 16712 2604
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17589 2635 17647 2641
rect 17589 2601 17601 2635
rect 17635 2632 17647 2635
rect 18046 2632 18052 2644
rect 17635 2604 18052 2632
rect 17635 2601 17647 2604
rect 17589 2595 17647 2601
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18230 2632 18236 2644
rect 18191 2604 18236 2632
rect 18230 2592 18236 2604
rect 18288 2592 18294 2644
rect 19334 2632 19340 2644
rect 19295 2604 19340 2632
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 20165 2635 20223 2641
rect 20165 2601 20177 2635
rect 20211 2632 20223 2635
rect 20714 2632 20720 2644
rect 20211 2604 20720 2632
rect 20211 2601 20223 2604
rect 20165 2595 20223 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 20901 2635 20959 2641
rect 20901 2601 20913 2635
rect 20947 2632 20959 2635
rect 21450 2632 21456 2644
rect 20947 2604 21456 2632
rect 20947 2601 20959 2604
rect 20901 2595 20959 2601
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 23750 2632 23756 2644
rect 23711 2604 23756 2632
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 23934 2592 23940 2644
rect 23992 2632 23998 2644
rect 24949 2635 25007 2641
rect 24949 2632 24961 2635
rect 23992 2604 24961 2632
rect 23992 2592 23998 2604
rect 24949 2601 24961 2604
rect 24995 2601 25007 2635
rect 24949 2595 25007 2601
rect 25406 2592 25412 2644
rect 25464 2632 25470 2644
rect 25501 2635 25559 2641
rect 25501 2632 25513 2635
rect 25464 2604 25513 2632
rect 25464 2592 25470 2604
rect 25501 2601 25513 2604
rect 25547 2601 25559 2635
rect 25501 2595 25559 2601
rect 28166 2592 28172 2644
rect 28224 2632 28230 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 28224 2604 28641 2632
rect 28224 2592 28230 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 31110 2632 31116 2644
rect 28629 2595 28687 2601
rect 29288 2604 31116 2632
rect 27062 2564 27068 2576
rect 2179 2536 11744 2564
rect 15396 2536 16620 2564
rect 16684 2536 27068 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 5307 2468 9076 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8444 2400 8953 2428
rect 8444 2388 8450 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 9048 2428 9076 2468
rect 15194 2428 15200 2440
rect 9048 2400 15200 2428
rect 8941 2391 8999 2397
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 1360 2332 1869 2360
rect 1360 2320 1366 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2648 2332 2789 2360
rect 2648 2320 2654 2332
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 15396 2292 15424 2536
rect 16592 2496 16620 2536
rect 27062 2524 27068 2536
rect 27120 2524 27126 2576
rect 27617 2567 27675 2573
rect 27617 2533 27629 2567
rect 27663 2564 27675 2567
rect 29288 2564 29316 2604
rect 31110 2592 31116 2604
rect 31168 2592 31174 2644
rect 35526 2632 35532 2644
rect 35487 2604 35532 2632
rect 35526 2592 35532 2604
rect 35584 2592 35590 2644
rect 38289 2635 38347 2641
rect 38289 2632 38301 2635
rect 35636 2604 38301 2632
rect 27663 2536 29316 2564
rect 29733 2567 29791 2573
rect 27663 2533 27675 2536
rect 27617 2527 27675 2533
rect 29733 2533 29745 2567
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 22278 2496 22284 2508
rect 16592 2468 16896 2496
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 15528 2332 15669 2360
rect 15528 2320 15534 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 15746 2292 15752 2304
rect 9171 2264 15424 2292
rect 15707 2264 15752 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 16868 2292 16896 2468
rect 20088 2468 22284 2496
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2428 17555 2431
rect 17954 2428 17960 2440
rect 17543 2400 17960 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 19242 2428 19248 2440
rect 19203 2400 19248 2428
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 20088 2437 20116 2468
rect 22278 2456 22284 2468
rect 22336 2456 22342 2508
rect 23017 2499 23075 2505
rect 23017 2465 23029 2499
rect 23063 2496 23075 2499
rect 25314 2496 25320 2508
rect 23063 2468 25320 2496
rect 23063 2465 23075 2468
rect 23017 2459 23075 2465
rect 25314 2456 25320 2468
rect 25372 2456 25378 2508
rect 29748 2496 29776 2527
rect 33778 2524 33784 2576
rect 33836 2564 33842 2576
rect 35636 2564 35664 2604
rect 38289 2601 38301 2604
rect 38335 2601 38347 2635
rect 38289 2595 38347 2601
rect 40405 2635 40463 2641
rect 40405 2601 40417 2635
rect 40451 2632 40463 2635
rect 40586 2632 40592 2644
rect 40451 2604 40592 2632
rect 40451 2601 40463 2604
rect 40405 2595 40463 2601
rect 40586 2592 40592 2604
rect 40644 2592 40650 2644
rect 40770 2592 40776 2644
rect 40828 2632 40834 2644
rect 41506 2632 41512 2644
rect 40828 2604 41512 2632
rect 40828 2592 40834 2604
rect 41506 2592 41512 2604
rect 41564 2592 41570 2644
rect 39301 2567 39359 2573
rect 39301 2564 39313 2567
rect 33836 2536 35664 2564
rect 35820 2536 39313 2564
rect 33836 2524 33842 2536
rect 35618 2496 35624 2508
rect 29748 2468 35624 2496
rect 35618 2456 35624 2468
rect 35676 2456 35682 2508
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 22373 2431 22431 2437
rect 22373 2397 22385 2431
rect 22419 2428 22431 2431
rect 22462 2428 22468 2440
rect 22419 2400 22468 2428
rect 22419 2397 22431 2400
rect 22373 2391 22431 2397
rect 22462 2388 22468 2400
rect 22520 2388 22526 2440
rect 22738 2428 22744 2440
rect 22699 2400 22744 2428
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 23658 2428 23664 2440
rect 23619 2400 23664 2428
rect 23658 2388 23664 2400
rect 23716 2388 23722 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 23768 2400 25697 2428
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 23198 2320 23204 2372
rect 23256 2360 23262 2372
rect 23768 2360 23796 2400
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 23256 2332 23796 2360
rect 23256 2320 23262 2332
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24544 2332 24869 2360
rect 24544 2320 24550 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 26237 2363 26295 2369
rect 26237 2329 26249 2363
rect 26283 2360 26295 2363
rect 26418 2360 26424 2372
rect 26283 2332 26424 2360
rect 26283 2329 26295 2332
rect 26237 2323 26295 2329
rect 26418 2320 26424 2332
rect 26476 2320 26482 2372
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 27120 2332 27445 2360
rect 27120 2320 27126 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 31294 2320 31300 2372
rect 31352 2360 31358 2372
rect 35820 2360 35848 2536
rect 39301 2533 39313 2536
rect 39347 2533 39359 2567
rect 42429 2567 42487 2573
rect 42429 2564 42441 2567
rect 39301 2527 39359 2533
rect 40420 2536 42441 2564
rect 36354 2456 36360 2508
rect 36412 2496 36418 2508
rect 36449 2499 36507 2505
rect 36449 2496 36461 2499
rect 36412 2468 36461 2496
rect 36412 2456 36418 2468
rect 36449 2465 36461 2468
rect 36495 2465 36507 2499
rect 39942 2496 39948 2508
rect 36449 2459 36507 2465
rect 37660 2468 39948 2496
rect 37660 2437 37688 2468
rect 39942 2456 39948 2468
rect 40000 2456 40006 2508
rect 40420 2440 40448 2536
rect 42429 2533 42441 2536
rect 42475 2533 42487 2567
rect 42429 2527 42487 2533
rect 44174 2524 44180 2576
rect 44232 2564 44238 2576
rect 44232 2536 47900 2564
rect 44232 2524 44238 2536
rect 41325 2499 41383 2505
rect 41325 2465 41337 2499
rect 41371 2496 41383 2499
rect 42334 2496 42340 2508
rect 41371 2468 42340 2496
rect 41371 2465 41383 2468
rect 41325 2459 41383 2465
rect 42334 2456 42340 2468
rect 42392 2456 42398 2508
rect 43070 2456 43076 2508
rect 43128 2496 43134 2508
rect 47872 2505 47900 2536
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 43128 2468 46489 2496
rect 43128 2456 43134 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 46477 2459 46535 2465
rect 47857 2499 47915 2505
rect 47857 2465 47869 2499
rect 47903 2465 47915 2499
rect 47857 2459 47915 2465
rect 37645 2431 37703 2437
rect 37645 2397 37657 2431
rect 37691 2397 37703 2431
rect 39666 2428 39672 2440
rect 37645 2391 37703 2397
rect 37936 2400 39672 2428
rect 31352 2332 35848 2360
rect 31352 2320 31358 2332
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 24394 2292 24400 2304
rect 16868 2264 24400 2292
rect 24394 2252 24400 2264
rect 24452 2252 24458 2304
rect 26326 2292 26332 2304
rect 26287 2264 26332 2292
rect 26326 2252 26332 2264
rect 26384 2252 26390 2304
rect 37461 2295 37519 2301
rect 37461 2261 37473 2295
rect 37507 2292 37519 2295
rect 37936 2292 37964 2400
rect 39666 2388 39672 2400
rect 39724 2428 39730 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39724 2400 40049 2428
rect 39724 2388 39730 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40402 2428 40408 2440
rect 40363 2400 40408 2428
rect 40037 2391 40095 2397
rect 40402 2388 40408 2400
rect 40460 2388 40466 2440
rect 40586 2388 40592 2440
rect 40644 2428 40650 2440
rect 41141 2431 41199 2437
rect 41141 2428 41153 2431
rect 40644 2400 41153 2428
rect 40644 2388 40650 2400
rect 41141 2397 41153 2400
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 41230 2388 41236 2440
rect 41288 2428 41294 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 41288 2400 42625 2428
rect 41288 2388 41294 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 46201 2431 46259 2437
rect 46201 2397 46213 2431
rect 46247 2428 46259 2431
rect 47026 2428 47032 2440
rect 46247 2400 47032 2428
rect 46247 2397 46259 2400
rect 46201 2391 46259 2397
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 38197 2363 38255 2369
rect 38197 2360 38209 2363
rect 38068 2332 38209 2360
rect 38068 2320 38074 2332
rect 38197 2329 38209 2332
rect 38243 2329 38255 2363
rect 38197 2323 38255 2329
rect 39117 2363 39175 2369
rect 39117 2329 39129 2363
rect 39163 2360 39175 2363
rect 39298 2360 39304 2372
rect 39163 2332 39304 2360
rect 39163 2329 39175 2332
rect 39117 2323 39175 2329
rect 39298 2320 39304 2332
rect 39356 2320 39362 2372
rect 40678 2320 40684 2372
rect 40736 2360 40742 2372
rect 41414 2360 41420 2372
rect 40736 2332 41420 2360
rect 40736 2320 40742 2332
rect 41414 2320 41420 2332
rect 41472 2320 41478 2372
rect 41598 2320 41604 2372
rect 41656 2360 41662 2372
rect 43916 2360 43944 2391
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 47673 2431 47731 2437
rect 47673 2397 47685 2431
rect 47719 2428 47731 2431
rect 48038 2428 48044 2440
rect 47719 2400 48044 2428
rect 47719 2397 47731 2400
rect 47673 2391 47731 2397
rect 48038 2388 48044 2400
rect 48096 2388 48102 2440
rect 41656 2332 43944 2360
rect 45373 2363 45431 2369
rect 41656 2320 41662 2332
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46382 2360 46388 2372
rect 45419 2332 46388 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 37507 2264 37964 2292
rect 40589 2295 40647 2301
rect 37507 2261 37519 2264
rect 37461 2255 37519 2261
rect 40589 2261 40601 2295
rect 40635 2292 40647 2295
rect 40770 2292 40776 2304
rect 40635 2264 40776 2292
rect 40635 2261 40647 2264
rect 40589 2255 40647 2261
rect 40770 2252 40776 2264
rect 40828 2252 40834 2304
rect 45462 2292 45468 2304
rect 45423 2264 45468 2292
rect 45462 2252 45468 2264
rect 45520 2252 45526 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 35618 2048 35624 2100
rect 35676 2088 35682 2100
rect 40678 2088 40684 2100
rect 35676 2060 40684 2088
rect 35676 2048 35682 2060
rect 40678 2048 40684 2060
rect 40736 2048 40742 2100
rect 23382 1980 23388 2032
rect 23440 2020 23446 2032
rect 45462 2020 45468 2032
rect 23440 1992 45468 2020
rect 23440 1980 23446 1992
rect 45462 1980 45468 1992
rect 45520 1980 45526 2032
rect 26326 1912 26332 1964
rect 26384 1952 26390 1964
rect 40310 1952 40316 1964
rect 26384 1924 40316 1952
rect 26384 1912 26390 1924
rect 40310 1912 40316 1924
rect 40368 1912 40374 1964
rect 15746 1844 15752 1896
rect 15804 1884 15810 1896
rect 36170 1884 36176 1896
rect 15804 1856 36176 1884
rect 15804 1844 15810 1856
rect 36170 1844 36176 1856
rect 36228 1844 36234 1896
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 34244 47200 34296 47252
rect 39764 47132 39816 47184
rect 1952 46996 2004 47048
rect 3240 46996 3292 47048
rect 4712 47039 4764 47048
rect 4712 47005 4721 47039
rect 4721 47005 4755 47039
rect 4755 47005 4764 47039
rect 4712 46996 4764 47005
rect 5816 46996 5868 47048
rect 7288 47039 7340 47048
rect 7288 47005 7297 47039
rect 7297 47005 7331 47039
rect 7331 47005 7340 47039
rect 7288 46996 7340 47005
rect 9036 46996 9088 47048
rect 11612 47039 11664 47048
rect 11612 47005 11621 47039
rect 11621 47005 11655 47039
rect 11655 47005 11664 47039
rect 11612 46996 11664 47005
rect 12256 46996 12308 47048
rect 12900 46996 12952 47048
rect 16488 46996 16540 47048
rect 16948 47039 17000 47048
rect 16948 47005 16957 47039
rect 16957 47005 16991 47039
rect 16991 47005 17000 47039
rect 16948 46996 17000 47005
rect 18696 46996 18748 47048
rect 19984 46996 20036 47048
rect 20352 47039 20404 47048
rect 20352 47005 20361 47039
rect 20361 47005 20395 47039
rect 20395 47005 20404 47039
rect 20352 46996 20404 47005
rect 24860 47039 24912 47048
rect 24860 47005 24869 47039
rect 24869 47005 24903 47039
rect 24903 47005 24912 47039
rect 24860 46996 24912 47005
rect 25504 47039 25556 47048
rect 25504 47005 25513 47039
rect 25513 47005 25547 47039
rect 25547 47005 25556 47039
rect 25504 46996 25556 47005
rect 4068 46971 4120 46980
rect 2596 46860 2648 46912
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 4988 46971 5040 46980
rect 4988 46937 4997 46971
rect 4997 46937 5031 46971
rect 5031 46937 5040 46971
rect 4988 46928 5040 46937
rect 6644 46971 6696 46980
rect 6644 46937 6653 46971
rect 6653 46937 6687 46971
rect 6687 46937 6696 46971
rect 6644 46928 6696 46937
rect 8208 46928 8260 46980
rect 11704 46928 11756 46980
rect 12440 46928 12492 46980
rect 13360 46928 13412 46980
rect 13544 46860 13596 46912
rect 14648 46928 14700 46980
rect 18880 46928 18932 46980
rect 32404 47064 32456 47116
rect 37648 47064 37700 47116
rect 43168 47107 43220 47116
rect 43168 47073 43177 47107
rect 43177 47073 43211 47107
rect 43211 47073 43220 47107
rect 43168 47064 43220 47073
rect 48320 47064 48372 47116
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 30932 46996 30984 47048
rect 38016 46996 38068 47048
rect 40132 46996 40184 47048
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 30196 46928 30248 46980
rect 31024 46928 31076 46980
rect 42708 46971 42760 46980
rect 29920 46903 29972 46912
rect 29920 46869 29929 46903
rect 29929 46869 29963 46903
rect 29963 46869 29972 46903
rect 29920 46860 29972 46869
rect 39304 46860 39356 46912
rect 42708 46937 42717 46971
rect 42717 46937 42751 46971
rect 42751 46937 42760 46971
rect 42708 46928 42760 46937
rect 45468 46928 45520 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1860 46631 1912 46640
rect 1860 46597 1869 46631
rect 1869 46597 1903 46631
rect 1903 46597 1912 46631
rect 1860 46588 1912 46597
rect 24860 46588 24912 46640
rect 27068 46588 27120 46640
rect 34060 46588 34112 46640
rect 47032 46631 47084 46640
rect 47032 46597 47041 46631
rect 47041 46597 47075 46631
rect 47075 46597 47084 46631
rect 47032 46588 47084 46597
rect 38016 46563 38068 46572
rect 38016 46529 38025 46563
rect 38025 46529 38059 46563
rect 38059 46529 38068 46563
rect 38016 46520 38068 46529
rect 47952 46563 48004 46572
rect 47952 46529 47961 46563
rect 47961 46529 47995 46563
rect 47995 46529 48004 46563
rect 47952 46520 48004 46529
rect 3884 46452 3936 46504
rect 3976 46452 4028 46504
rect 13728 46495 13780 46504
rect 13728 46461 13737 46495
rect 13737 46461 13771 46495
rect 13771 46461 13780 46495
rect 13728 46452 13780 46461
rect 14188 46495 14240 46504
rect 14188 46461 14197 46495
rect 14197 46461 14231 46495
rect 14231 46461 14240 46495
rect 14188 46452 14240 46461
rect 19432 46495 19484 46504
rect 19432 46461 19441 46495
rect 19441 46461 19475 46495
rect 19475 46461 19484 46495
rect 19432 46452 19484 46461
rect 20168 46452 20220 46504
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32496 46495 32548 46504
rect 32496 46461 32505 46495
rect 32505 46461 32539 46495
rect 32539 46461 32548 46495
rect 32496 46452 32548 46461
rect 33416 46452 33468 46504
rect 38200 46495 38252 46504
rect 4620 46384 4672 46436
rect 32220 46384 32272 46436
rect 38200 46461 38209 46495
rect 38209 46461 38243 46495
rect 38243 46461 38252 46495
rect 38200 46452 38252 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 45376 46495 45428 46504
rect 42248 46384 42300 46436
rect 45376 46461 45385 46495
rect 45385 46461 45419 46495
rect 45419 46461 45428 46495
rect 45376 46452 45428 46461
rect 45652 46384 45704 46436
rect 2320 46316 2372 46368
rect 2780 46316 2832 46368
rect 10416 46316 10468 46368
rect 20720 46316 20772 46368
rect 41052 46316 41104 46368
rect 47216 46316 47268 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3884 46155 3936 46164
rect 3884 46121 3893 46155
rect 3893 46121 3927 46155
rect 3927 46121 3936 46155
rect 3884 46112 3936 46121
rect 4620 46155 4672 46164
rect 4620 46121 4629 46155
rect 4629 46121 4663 46155
rect 4663 46121 4672 46155
rect 4620 46112 4672 46121
rect 19432 46112 19484 46164
rect 20168 46155 20220 46164
rect 20168 46121 20177 46155
rect 20177 46121 20211 46155
rect 20211 46121 20220 46155
rect 20168 46112 20220 46121
rect 24768 46112 24820 46164
rect 32496 46112 32548 46164
rect 33416 46155 33468 46164
rect 33416 46121 33425 46155
rect 33425 46121 33459 46155
rect 33459 46121 33468 46155
rect 33416 46112 33468 46121
rect 38200 46155 38252 46164
rect 38200 46121 38209 46155
rect 38209 46121 38243 46155
rect 38243 46121 38252 46155
rect 38200 46112 38252 46121
rect 10416 46019 10468 46028
rect 10416 45985 10425 46019
rect 10425 45985 10459 46019
rect 10459 45985 10468 46019
rect 10416 45976 10468 45985
rect 10968 45976 11020 46028
rect 20720 46019 20772 46028
rect 20720 45985 20729 46019
rect 20729 45985 20763 46019
rect 20763 45985 20772 46019
rect 20720 45976 20772 45985
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25504 45976 25556 46028
rect 25780 46019 25832 46028
rect 25780 45985 25789 46019
rect 25789 45985 25823 46019
rect 25823 45985 25832 46019
rect 25780 45976 25832 45985
rect 45836 46044 45888 46096
rect 41052 46019 41104 46028
rect 41052 45985 41061 46019
rect 41061 45985 41095 46019
rect 41095 45985 41104 46019
rect 41052 45976 41104 45985
rect 42524 46019 42576 46028
rect 42524 45985 42533 46019
rect 42533 45985 42567 46019
rect 42567 45985 42576 46019
rect 42524 45976 42576 45985
rect 48136 46019 48188 46028
rect 48136 45985 48145 46019
rect 48145 45985 48179 46019
rect 48179 45985 48188 46019
rect 48136 45976 48188 45985
rect 3056 45908 3108 45960
rect 20076 45951 20128 45960
rect 20076 45917 20085 45951
rect 20085 45917 20119 45951
rect 20119 45917 20128 45951
rect 20076 45908 20128 45917
rect 24860 45908 24912 45960
rect 38108 45951 38160 45960
rect 10600 45883 10652 45892
rect 2872 45815 2924 45824
rect 2872 45781 2881 45815
rect 2881 45781 2915 45815
rect 2915 45781 2924 45815
rect 2872 45772 2924 45781
rect 10600 45849 10609 45883
rect 10609 45849 10643 45883
rect 10643 45849 10652 45883
rect 10600 45840 10652 45849
rect 20904 45883 20956 45892
rect 20904 45849 20913 45883
rect 20913 45849 20947 45883
rect 20947 45849 20956 45883
rect 20904 45840 20956 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 38108 45917 38117 45951
rect 38117 45917 38151 45951
rect 38151 45917 38160 45951
rect 38108 45908 38160 45917
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 46296 45951 46348 45960
rect 46296 45917 46305 45951
rect 46305 45917 46339 45951
rect 46339 45917 46348 45951
rect 46296 45908 46348 45917
rect 40040 45840 40092 45892
rect 41236 45883 41288 45892
rect 41236 45849 41245 45883
rect 41245 45849 41279 45883
rect 41279 45849 41288 45883
rect 41236 45840 41288 45849
rect 44456 45840 44508 45892
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 10508 45772 10560 45824
rect 45560 45772 45612 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 10600 45611 10652 45620
rect 10600 45577 10609 45611
rect 10609 45577 10643 45611
rect 10643 45577 10652 45611
rect 10600 45568 10652 45577
rect 13728 45611 13780 45620
rect 13728 45577 13737 45611
rect 13737 45577 13771 45611
rect 13771 45577 13780 45611
rect 13728 45568 13780 45577
rect 16120 45568 16172 45620
rect 17408 45568 17460 45620
rect 20904 45568 20956 45620
rect 25412 45611 25464 45620
rect 25412 45577 25421 45611
rect 25421 45577 25455 45611
rect 25455 45577 25464 45611
rect 25412 45568 25464 45577
rect 42616 45568 42668 45620
rect 45100 45568 45152 45620
rect 2872 45500 2924 45552
rect 10508 45475 10560 45484
rect 10508 45441 10517 45475
rect 10517 45441 10551 45475
rect 10551 45441 10560 45475
rect 24860 45500 24912 45552
rect 42708 45543 42760 45552
rect 42708 45509 42717 45543
rect 42717 45509 42751 45543
rect 42751 45509 42760 45543
rect 42708 45500 42760 45509
rect 10508 45432 10560 45441
rect 2780 45364 2832 45416
rect 2964 45407 3016 45416
rect 2964 45373 2973 45407
rect 2973 45373 3007 45407
rect 3007 45373 3016 45407
rect 2964 45364 3016 45373
rect 26056 45432 26108 45484
rect 43996 45500 44048 45552
rect 46204 45568 46256 45620
rect 44180 45432 44232 45484
rect 27344 45364 27396 45416
rect 38660 45407 38712 45416
rect 38660 45373 38669 45407
rect 38669 45373 38703 45407
rect 38703 45373 38712 45407
rect 38660 45364 38712 45373
rect 38844 45407 38896 45416
rect 38844 45373 38853 45407
rect 38853 45373 38887 45407
rect 38887 45373 38896 45407
rect 38844 45364 38896 45373
rect 39856 45407 39908 45416
rect 39856 45373 39865 45407
rect 39865 45373 39899 45407
rect 39899 45373 39908 45407
rect 39856 45364 39908 45373
rect 45100 45364 45152 45416
rect 40684 45296 40736 45348
rect 42800 45296 42852 45348
rect 44088 45271 44140 45280
rect 44088 45237 44097 45271
rect 44097 45237 44131 45271
rect 44131 45237 44140 45271
rect 44088 45228 44140 45237
rect 44272 45296 44324 45348
rect 47584 45296 47636 45348
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 38844 45067 38896 45076
rect 38844 45033 38853 45067
rect 38853 45033 38887 45067
rect 38887 45033 38896 45067
rect 38844 45024 38896 45033
rect 41236 45024 41288 45076
rect 45100 45067 45152 45076
rect 45100 45033 45109 45067
rect 45109 45033 45143 45067
rect 45143 45033 45152 45067
rect 45100 45024 45152 45033
rect 46480 45024 46532 45076
rect 45376 44956 45428 45008
rect 47032 44888 47084 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 28632 44820 28684 44872
rect 40040 44820 40092 44872
rect 40316 44863 40368 44872
rect 40316 44829 40325 44863
rect 40325 44829 40359 44863
rect 40359 44829 40368 44863
rect 40316 44820 40368 44829
rect 44272 44863 44324 44872
rect 44272 44829 44281 44863
rect 44281 44829 44315 44863
rect 44315 44829 44324 44863
rect 44272 44820 44324 44829
rect 45008 44863 45060 44872
rect 45008 44829 45017 44863
rect 45017 44829 45051 44863
rect 45051 44829 45060 44863
rect 45008 44820 45060 44829
rect 38660 44684 38712 44736
rect 47676 44752 47728 44804
rect 45836 44684 45888 44736
rect 46756 44684 46808 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 45468 44480 45520 44532
rect 47676 44523 47728 44532
rect 47676 44489 47685 44523
rect 47685 44489 47719 44523
rect 47719 44489 47728 44523
rect 47676 44480 47728 44489
rect 40684 44412 40736 44464
rect 20076 44344 20128 44396
rect 45192 44344 45244 44396
rect 45744 44387 45796 44396
rect 45744 44353 45753 44387
rect 45753 44353 45787 44387
rect 45787 44353 45796 44387
rect 45744 44344 45796 44353
rect 46572 44344 46624 44396
rect 45928 44276 45980 44328
rect 46940 44183 46992 44192
rect 46940 44149 46949 44183
rect 46949 44149 46983 44183
rect 46983 44149 46992 44183
rect 46940 44140 46992 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 46940 43800 46992 43852
rect 48228 43800 48280 43852
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 1676 43231 1728 43240
rect 1676 43197 1685 43231
rect 1685 43197 1719 43231
rect 1719 43197 1728 43231
rect 1676 43188 1728 43197
rect 46296 43188 46348 43240
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 46296 42687 46348 42696
rect 46296 42653 46305 42687
rect 46305 42653 46339 42687
rect 46339 42653 46348 42687
rect 46296 42644 46348 42653
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 46296 42168 46348 42220
rect 47584 42211 47636 42220
rect 47584 42177 47593 42211
rect 47593 42177 47627 42211
rect 47627 42177 47636 42211
rect 47584 42168 47636 42177
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47676 41624 47728 41676
rect 48136 41599 48188 41608
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46940 41488 46992 41540
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46940 41259 46992 41268
rect 46940 41225 46949 41259
rect 46949 41225 46983 41259
rect 46983 41225 46992 41259
rect 46940 41216 46992 41225
rect 2136 41123 2188 41132
rect 2136 41089 2145 41123
rect 2145 41089 2179 41123
rect 2179 41089 2188 41123
rect 2136 41080 2188 41089
rect 20076 41080 20128 41132
rect 46756 41080 46808 41132
rect 48044 41080 48096 41132
rect 47952 40876 48004 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 1768 40332 1820 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 46940 39312 46992 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 3332 39040 3384 39092
rect 7564 39040 7616 39092
rect 26148 39083 26200 39092
rect 26148 39049 26157 39083
rect 26157 39049 26191 39083
rect 26191 39049 26200 39083
rect 46940 39083 46992 39092
rect 26148 39040 26200 39049
rect 25320 38904 25372 38956
rect 25964 38947 26016 38956
rect 25964 38913 25973 38947
rect 25973 38913 26007 38947
rect 26007 38913 26016 38947
rect 25964 38904 26016 38913
rect 46940 39049 46949 39083
rect 46949 39049 46983 39083
rect 46983 39049 46992 39083
rect 46940 39040 46992 39049
rect 46020 38904 46072 38956
rect 47676 38947 47728 38956
rect 47676 38913 47685 38947
rect 47685 38913 47719 38947
rect 47719 38913 47728 38947
rect 47676 38904 47728 38913
rect 8208 38836 8260 38888
rect 38108 38836 38160 38888
rect 47860 38879 47912 38888
rect 25964 38768 26016 38820
rect 47860 38845 47869 38879
rect 47869 38845 47903 38879
rect 47903 38845 47912 38879
rect 47860 38836 47912 38845
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 26148 38335 26200 38344
rect 26148 38301 26157 38335
rect 26157 38301 26191 38335
rect 26191 38301 26200 38335
rect 26148 38292 26200 38301
rect 46940 38292 46992 38344
rect 26332 38156 26384 38208
rect 44272 38156 44324 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 26148 37816 26200 37868
rect 47584 37859 47636 37868
rect 25412 37748 25464 37800
rect 26056 37791 26108 37800
rect 26056 37757 26065 37791
rect 26065 37757 26099 37791
rect 26099 37757 26108 37791
rect 26056 37748 26108 37757
rect 26792 37748 26844 37800
rect 27344 37791 27396 37800
rect 27344 37757 27353 37791
rect 27353 37757 27387 37791
rect 27387 37757 27396 37791
rect 47584 37825 47593 37859
rect 47593 37825 47627 37859
rect 47627 37825 47636 37859
rect 47584 37816 47636 37825
rect 27344 37748 27396 37757
rect 47676 37655 47728 37664
rect 47676 37621 47685 37655
rect 47685 37621 47719 37655
rect 47719 37621 47728 37655
rect 47676 37612 47728 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 26148 37247 26200 37256
rect 26148 37213 26157 37247
rect 26157 37213 26191 37247
rect 26191 37213 26200 37247
rect 26148 37204 26200 37213
rect 26700 37136 26752 37188
rect 40316 37136 40368 37188
rect 47676 37136 47728 37188
rect 46940 37068 46992 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 27528 36796 27580 36848
rect 12440 36728 12492 36780
rect 26976 36660 27028 36712
rect 27528 36703 27580 36712
rect 27528 36669 27537 36703
rect 27537 36669 27571 36703
rect 27571 36669 27580 36703
rect 27528 36660 27580 36669
rect 26424 36567 26476 36576
rect 26424 36533 26433 36567
rect 26433 36533 26467 36567
rect 26467 36533 26476 36567
rect 26424 36524 26476 36533
rect 26516 36524 26568 36576
rect 45560 36524 45612 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 26976 36363 27028 36372
rect 26976 36329 26985 36363
rect 26985 36329 27019 36363
rect 27019 36329 27028 36363
rect 26976 36320 27028 36329
rect 2780 36227 2832 36236
rect 2780 36193 2789 36227
rect 2789 36193 2823 36227
rect 2823 36193 2832 36227
rect 2780 36184 2832 36193
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 26516 36184 26568 36236
rect 27436 36184 27488 36236
rect 25780 36116 25832 36168
rect 26608 36159 26660 36168
rect 26608 36125 26617 36159
rect 26617 36125 26651 36159
rect 26651 36125 26660 36159
rect 26608 36116 26660 36125
rect 2228 36048 2280 36100
rect 23480 36023 23532 36032
rect 23480 35989 23489 36023
rect 23489 35989 23523 36023
rect 23523 35989 23532 36023
rect 23480 35980 23532 35989
rect 25688 35980 25740 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 26608 35776 26660 35828
rect 22836 35708 22888 35760
rect 25688 35708 25740 35760
rect 30932 35708 30984 35760
rect 1400 35640 1452 35692
rect 26424 35640 26476 35692
rect 23480 35572 23532 35624
rect 24676 35615 24728 35624
rect 24676 35581 24685 35615
rect 24685 35581 24719 35615
rect 24719 35581 24728 35615
rect 24676 35572 24728 35581
rect 24952 35615 25004 35624
rect 24952 35581 24961 35615
rect 24961 35581 24995 35615
rect 24995 35581 25004 35615
rect 24952 35572 25004 35581
rect 28448 35572 28500 35624
rect 29920 35615 29972 35624
rect 23480 35436 23532 35488
rect 24676 35436 24728 35488
rect 26516 35436 26568 35488
rect 26976 35479 27028 35488
rect 26976 35445 26985 35479
rect 26985 35445 27019 35479
rect 27019 35445 27028 35479
rect 26976 35436 27028 35445
rect 27436 35436 27488 35488
rect 29920 35581 29929 35615
rect 29929 35581 29963 35615
rect 29963 35581 29972 35615
rect 29920 35572 29972 35581
rect 30288 35572 30340 35624
rect 31116 35436 31168 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 2228 35275 2280 35284
rect 2228 35241 2237 35275
rect 2237 35241 2271 35275
rect 2271 35241 2280 35275
rect 2228 35232 2280 35241
rect 22836 35275 22888 35284
rect 22836 35241 22845 35275
rect 22845 35241 22879 35275
rect 22879 35241 22888 35275
rect 22836 35232 22888 35241
rect 24952 35232 25004 35284
rect 24676 35164 24728 35216
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 1584 35028 1636 35037
rect 2228 35028 2280 35080
rect 22008 35028 22060 35080
rect 24492 35071 24544 35080
rect 24492 35037 24501 35071
rect 24501 35037 24535 35071
rect 24535 35037 24544 35071
rect 24492 35028 24544 35037
rect 26424 35164 26476 35216
rect 29920 35232 29972 35284
rect 30196 35275 30248 35284
rect 30196 35241 30205 35275
rect 30205 35241 30239 35275
rect 30239 35241 30248 35275
rect 30196 35232 30248 35241
rect 30932 35232 30984 35284
rect 29736 35096 29788 35148
rect 1492 34892 1544 34944
rect 24952 34892 25004 34944
rect 26976 35028 27028 35080
rect 30104 35028 30156 35080
rect 48136 35071 48188 35080
rect 26516 34960 26568 35012
rect 27804 34960 27856 35012
rect 28816 34960 28868 35012
rect 28908 34960 28960 35012
rect 48136 35037 48145 35071
rect 48145 35037 48179 35071
rect 48179 35037 48188 35071
rect 48136 35028 48188 35037
rect 27344 34892 27396 34944
rect 29184 34892 29236 34944
rect 29828 34935 29880 34944
rect 29828 34901 29837 34935
rect 29837 34901 29871 34935
rect 29871 34901 29880 34935
rect 29828 34892 29880 34901
rect 31852 34892 31904 34944
rect 47124 34892 47176 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 23480 34688 23532 34740
rect 27988 34688 28040 34740
rect 28816 34731 28868 34740
rect 28816 34697 28825 34731
rect 28825 34697 28859 34731
rect 28859 34697 28868 34731
rect 28816 34688 28868 34697
rect 30104 34731 30156 34740
rect 30104 34697 30113 34731
rect 30113 34697 30147 34731
rect 30147 34697 30156 34731
rect 30104 34688 30156 34697
rect 26516 34620 26568 34672
rect 23204 34552 23256 34604
rect 24952 34552 25004 34604
rect 25780 34552 25832 34604
rect 23572 34484 23624 34536
rect 24492 34484 24544 34536
rect 25136 34484 25188 34536
rect 26884 34552 26936 34604
rect 28908 34552 28960 34604
rect 33508 34620 33560 34672
rect 30288 34552 30340 34604
rect 48136 34595 48188 34604
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 27252 34416 27304 34468
rect 29184 34416 29236 34468
rect 20812 34348 20864 34400
rect 22652 34348 22704 34400
rect 22836 34348 22888 34400
rect 24952 34348 25004 34400
rect 25964 34348 26016 34400
rect 30104 34348 30156 34400
rect 30380 34348 30432 34400
rect 47860 34348 47912 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 22652 34187 22704 34196
rect 22652 34153 22661 34187
rect 22661 34153 22695 34187
rect 22695 34153 22704 34187
rect 22652 34144 22704 34153
rect 23204 34187 23256 34196
rect 23204 34153 23213 34187
rect 23213 34153 23247 34187
rect 23247 34153 23256 34187
rect 23204 34144 23256 34153
rect 26516 34144 26568 34196
rect 29828 34144 29880 34196
rect 20812 34076 20864 34128
rect 22008 34076 22060 34128
rect 16948 34008 17000 34060
rect 20812 33983 20864 33992
rect 20812 33949 20821 33983
rect 20821 33949 20855 33983
rect 20855 33949 20864 33983
rect 20812 33940 20864 33949
rect 21916 33983 21968 33992
rect 21916 33949 21925 33983
rect 21925 33949 21959 33983
rect 21959 33949 21968 33983
rect 21916 33940 21968 33949
rect 20904 33847 20956 33856
rect 20904 33813 20913 33847
rect 20913 33813 20947 33847
rect 20947 33813 20956 33847
rect 20904 33804 20956 33813
rect 22744 33940 22796 33992
rect 29552 34076 29604 34128
rect 24216 34008 24268 34060
rect 24676 34008 24728 34060
rect 26516 34008 26568 34060
rect 26148 33940 26200 33992
rect 27252 34008 27304 34060
rect 29000 34008 29052 34060
rect 30380 34008 30432 34060
rect 31116 34051 31168 34060
rect 31116 34017 31125 34051
rect 31125 34017 31159 34051
rect 31159 34017 31168 34051
rect 31116 34008 31168 34017
rect 28448 33983 28500 33992
rect 28448 33949 28457 33983
rect 28457 33949 28491 33983
rect 28491 33949 28500 33983
rect 28448 33940 28500 33949
rect 29644 33940 29696 33992
rect 22836 33872 22888 33924
rect 24676 33915 24728 33924
rect 24676 33881 24685 33915
rect 24685 33881 24719 33915
rect 24719 33881 24728 33915
rect 24676 33872 24728 33881
rect 25136 33872 25188 33924
rect 22284 33804 22336 33856
rect 29368 33872 29420 33924
rect 26148 33847 26200 33856
rect 26148 33813 26157 33847
rect 26157 33813 26191 33847
rect 26191 33813 26200 33847
rect 26148 33804 26200 33813
rect 27068 33847 27120 33856
rect 27068 33813 27077 33847
rect 27077 33813 27111 33847
rect 27111 33813 27120 33847
rect 27068 33804 27120 33813
rect 27160 33804 27212 33856
rect 33324 33983 33376 33992
rect 29828 33872 29880 33924
rect 33324 33949 33333 33983
rect 33333 33949 33367 33983
rect 33367 33949 33376 33983
rect 33324 33940 33376 33949
rect 33508 33983 33560 33992
rect 33508 33949 33517 33983
rect 33517 33949 33551 33983
rect 33551 33949 33560 33983
rect 33508 33940 33560 33949
rect 47952 33940 48004 33992
rect 30104 33872 30156 33924
rect 31392 33915 31444 33924
rect 31392 33881 31401 33915
rect 31401 33881 31435 33915
rect 31435 33881 31444 33915
rect 31392 33872 31444 33881
rect 31852 33872 31904 33924
rect 30288 33804 30340 33856
rect 31300 33804 31352 33856
rect 32404 33804 32456 33856
rect 33508 33847 33560 33856
rect 33508 33813 33517 33847
rect 33517 33813 33551 33847
rect 33551 33813 33560 33847
rect 33508 33804 33560 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 16028 33575 16080 33584
rect 16028 33541 16037 33575
rect 16037 33541 16071 33575
rect 16071 33541 16080 33575
rect 16028 33532 16080 33541
rect 2688 33507 2740 33516
rect 2688 33473 2697 33507
rect 2697 33473 2731 33507
rect 2731 33473 2740 33507
rect 2688 33464 2740 33473
rect 23480 33600 23532 33652
rect 24676 33600 24728 33652
rect 20904 33464 20956 33516
rect 27160 33600 27212 33652
rect 27344 33643 27396 33652
rect 27344 33609 27353 33643
rect 27353 33609 27387 33643
rect 27387 33609 27396 33643
rect 27344 33600 27396 33609
rect 27804 33600 27856 33652
rect 29000 33600 29052 33652
rect 29828 33643 29880 33652
rect 29828 33609 29837 33643
rect 29837 33609 29871 33643
rect 29871 33609 29880 33643
rect 29828 33600 29880 33609
rect 31392 33600 31444 33652
rect 27068 33532 27120 33584
rect 25872 33464 25924 33516
rect 26884 33464 26936 33516
rect 27252 33464 27304 33516
rect 29460 33532 29512 33584
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 13636 33396 13688 33448
rect 14372 33439 14424 33448
rect 14372 33405 14381 33439
rect 14381 33405 14415 33439
rect 14415 33405 14424 33439
rect 14372 33396 14424 33405
rect 22008 33396 22060 33448
rect 24308 33396 24360 33448
rect 26148 33396 26200 33448
rect 22376 33328 22428 33380
rect 28080 33439 28132 33448
rect 28080 33405 28089 33439
rect 28089 33405 28123 33439
rect 28123 33405 28132 33439
rect 28080 33396 28132 33405
rect 28448 33464 28500 33516
rect 29000 33507 29052 33516
rect 29000 33473 29009 33507
rect 29009 33473 29043 33507
rect 29043 33473 29052 33507
rect 29184 33507 29236 33516
rect 29000 33464 29052 33473
rect 29184 33473 29193 33507
rect 29193 33473 29227 33507
rect 29227 33473 29236 33507
rect 29184 33464 29236 33473
rect 30196 33464 30248 33516
rect 30840 33507 30892 33516
rect 30840 33473 30849 33507
rect 30849 33473 30883 33507
rect 30883 33473 30892 33507
rect 30840 33464 30892 33473
rect 31300 33464 31352 33516
rect 33140 33600 33192 33652
rect 32956 33532 33008 33584
rect 28540 33396 28592 33448
rect 31668 33396 31720 33448
rect 32404 33507 32456 33516
rect 32404 33473 32413 33507
rect 32413 33473 32447 33507
rect 32447 33473 32456 33507
rect 32404 33464 32456 33473
rect 32772 33464 32824 33516
rect 35440 33532 35492 33584
rect 46112 33532 46164 33584
rect 32956 33396 33008 33448
rect 33692 33396 33744 33448
rect 34428 33439 34480 33448
rect 34428 33405 34437 33439
rect 34437 33405 34471 33439
rect 34471 33405 34480 33439
rect 34428 33396 34480 33405
rect 33416 33371 33468 33380
rect 2780 33303 2832 33312
rect 2780 33269 2789 33303
rect 2789 33269 2823 33303
rect 2823 33269 2832 33303
rect 2780 33260 2832 33269
rect 3976 33260 4028 33312
rect 21732 33260 21784 33312
rect 21916 33260 21968 33312
rect 23388 33260 23440 33312
rect 25136 33260 25188 33312
rect 26976 33303 27028 33312
rect 26976 33269 26985 33303
rect 26985 33269 27019 33303
rect 27019 33269 27028 33303
rect 26976 33260 27028 33269
rect 28172 33260 28224 33312
rect 28448 33260 28500 33312
rect 33416 33337 33425 33371
rect 33425 33337 33459 33371
rect 33459 33337 33468 33371
rect 33416 33328 33468 33337
rect 30288 33260 30340 33312
rect 32588 33303 32640 33312
rect 32588 33269 32597 33303
rect 32597 33269 32631 33303
rect 32631 33269 32640 33303
rect 32588 33260 32640 33269
rect 32680 33260 32732 33312
rect 47308 33260 47360 33312
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 11704 33056 11756 33108
rect 22008 33056 22060 33108
rect 25136 33099 25188 33108
rect 25136 33065 25145 33099
rect 25145 33065 25179 33099
rect 25179 33065 25188 33099
rect 25136 33056 25188 33065
rect 26056 33099 26108 33108
rect 26056 33065 26065 33099
rect 26065 33065 26099 33099
rect 26099 33065 26108 33099
rect 26056 33056 26108 33065
rect 29092 33056 29144 33108
rect 30840 33056 30892 33108
rect 32404 33056 32456 33108
rect 32772 33099 32824 33108
rect 32772 33065 32781 33099
rect 32781 33065 32815 33099
rect 32815 33065 32824 33099
rect 32772 33056 32824 33065
rect 33324 33056 33376 33108
rect 34428 33056 34480 33108
rect 35440 33056 35492 33108
rect 1492 32988 1544 33040
rect 23572 32988 23624 33040
rect 28080 32988 28132 33040
rect 28540 32988 28592 33040
rect 29828 32988 29880 33040
rect 33140 32988 33192 33040
rect 11704 32963 11756 32972
rect 11704 32929 11713 32963
rect 11713 32929 11747 32963
rect 11747 32929 11756 32963
rect 11704 32920 11756 32929
rect 16120 32920 16172 32972
rect 25872 32963 25924 32972
rect 25872 32929 25881 32963
rect 25881 32929 25915 32963
rect 25915 32929 25924 32963
rect 25872 32920 25924 32929
rect 26240 32920 26292 32972
rect 26884 32963 26936 32972
rect 26884 32929 26893 32963
rect 26893 32929 26927 32963
rect 26927 32929 26936 32963
rect 26884 32920 26936 32929
rect 27804 32920 27856 32972
rect 30104 32920 30156 32972
rect 3976 32895 4028 32904
rect 3976 32861 3985 32895
rect 3985 32861 4019 32895
rect 4019 32861 4028 32895
rect 3976 32852 4028 32861
rect 13268 32852 13320 32904
rect 3240 32827 3292 32836
rect 3240 32793 3249 32827
rect 3249 32793 3283 32827
rect 3283 32793 3292 32827
rect 3240 32784 3292 32793
rect 9680 32784 9732 32836
rect 13544 32852 13596 32904
rect 20352 32852 20404 32904
rect 22376 32895 22428 32904
rect 22376 32861 22385 32895
rect 22385 32861 22419 32895
rect 22419 32861 22428 32895
rect 22376 32852 22428 32861
rect 22468 32895 22520 32904
rect 22468 32861 22477 32895
rect 22477 32861 22511 32895
rect 22511 32861 22520 32895
rect 22468 32852 22520 32861
rect 22652 32852 22704 32904
rect 24952 32895 25004 32904
rect 11796 32716 11848 32768
rect 22008 32784 22060 32836
rect 24952 32861 24961 32895
rect 24961 32861 24995 32895
rect 24995 32861 25004 32895
rect 24952 32852 25004 32861
rect 25228 32895 25280 32904
rect 25228 32861 25237 32895
rect 25237 32861 25271 32895
rect 25271 32861 25280 32895
rect 25228 32852 25280 32861
rect 26148 32852 26200 32904
rect 27252 32852 27304 32904
rect 25780 32827 25832 32836
rect 25780 32793 25789 32827
rect 25789 32793 25823 32827
rect 25823 32793 25832 32827
rect 25780 32784 25832 32793
rect 27988 32827 28040 32836
rect 27988 32793 28013 32827
rect 28013 32793 28040 32827
rect 29000 32852 29052 32904
rect 30380 32852 30432 32904
rect 31300 32920 31352 32972
rect 32956 32963 33008 32972
rect 32956 32929 32965 32963
rect 32965 32929 32999 32963
rect 32999 32929 33008 32963
rect 32956 32920 33008 32929
rect 33508 32920 33560 32972
rect 27988 32784 28040 32793
rect 29184 32784 29236 32836
rect 29644 32784 29696 32836
rect 31208 32852 31260 32904
rect 32680 32895 32732 32904
rect 32680 32861 32689 32895
rect 32689 32861 32723 32895
rect 32723 32861 32732 32895
rect 32680 32852 32732 32861
rect 33416 32895 33468 32904
rect 33416 32861 33425 32895
rect 33425 32861 33459 32895
rect 33459 32861 33468 32895
rect 33416 32852 33468 32861
rect 33600 32895 33652 32904
rect 33600 32861 33609 32895
rect 33609 32861 33643 32895
rect 33643 32861 33652 32895
rect 33600 32852 33652 32861
rect 33876 32852 33928 32904
rect 47124 32963 47176 32972
rect 47124 32929 47133 32963
rect 47133 32929 47167 32963
rect 47167 32929 47176 32963
rect 47124 32920 47176 32929
rect 47400 32963 47452 32972
rect 47400 32929 47409 32963
rect 47409 32929 47443 32963
rect 47443 32929 47452 32963
rect 47400 32920 47452 32929
rect 34704 32852 34756 32904
rect 46296 32852 46348 32904
rect 46480 32784 46532 32836
rect 47308 32784 47360 32836
rect 22192 32716 22244 32768
rect 23204 32716 23256 32768
rect 26240 32759 26292 32768
rect 26240 32725 26249 32759
rect 26249 32725 26283 32759
rect 26283 32725 26292 32759
rect 26240 32716 26292 32725
rect 27436 32716 27488 32768
rect 28540 32716 28592 32768
rect 29368 32716 29420 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 14372 32512 14424 32564
rect 22468 32512 22520 32564
rect 23388 32555 23440 32564
rect 23388 32521 23397 32555
rect 23397 32521 23431 32555
rect 23431 32521 23440 32555
rect 23388 32512 23440 32521
rect 28540 32512 28592 32564
rect 2688 32487 2740 32496
rect 2688 32453 2697 32487
rect 2697 32453 2731 32487
rect 2731 32453 2740 32487
rect 2688 32444 2740 32453
rect 11796 32487 11848 32496
rect 11796 32453 11805 32487
rect 11805 32453 11839 32487
rect 11839 32453 11848 32487
rect 11796 32444 11848 32453
rect 12808 32444 12860 32496
rect 22652 32444 22704 32496
rect 24584 32444 24636 32496
rect 25136 32444 25188 32496
rect 26056 32444 26108 32496
rect 27988 32444 28040 32496
rect 29276 32512 29328 32564
rect 29552 32512 29604 32564
rect 29644 32512 29696 32564
rect 33416 32512 33468 32564
rect 37648 32555 37700 32564
rect 37648 32521 37657 32555
rect 37657 32521 37691 32555
rect 37691 32521 37700 32555
rect 37648 32512 37700 32521
rect 28816 32444 28868 32496
rect 29000 32444 29052 32496
rect 13544 32376 13596 32428
rect 21732 32376 21784 32428
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 22376 32376 22428 32428
rect 24952 32376 25004 32428
rect 3240 32351 3292 32360
rect 3240 32317 3249 32351
rect 3249 32317 3283 32351
rect 3283 32317 3292 32351
rect 3240 32308 3292 32317
rect 11520 32351 11572 32360
rect 11520 32317 11529 32351
rect 11529 32317 11563 32351
rect 11563 32317 11572 32351
rect 11520 32308 11572 32317
rect 1952 32172 2004 32224
rect 9404 32240 9456 32292
rect 14096 32308 14148 32360
rect 22468 32308 22520 32360
rect 23112 32351 23164 32360
rect 23112 32317 23121 32351
rect 23121 32317 23155 32351
rect 23155 32317 23164 32351
rect 23112 32308 23164 32317
rect 25872 32308 25924 32360
rect 28908 32376 28960 32428
rect 29460 32487 29512 32496
rect 29460 32453 29477 32487
rect 29477 32453 29511 32487
rect 29511 32453 29512 32487
rect 29460 32444 29512 32453
rect 30104 32419 30156 32428
rect 30104 32385 30119 32419
rect 30119 32385 30153 32419
rect 30153 32385 30156 32419
rect 32588 32444 32640 32496
rect 32956 32444 33008 32496
rect 30104 32376 30156 32385
rect 31208 32419 31260 32428
rect 29184 32308 29236 32360
rect 29644 32351 29696 32360
rect 29644 32317 29653 32351
rect 29653 32317 29687 32351
rect 29687 32317 29696 32351
rect 31208 32385 31217 32419
rect 31217 32385 31251 32419
rect 31251 32385 31260 32419
rect 31208 32376 31260 32385
rect 33232 32419 33284 32428
rect 33232 32385 33241 32419
rect 33241 32385 33275 32419
rect 33275 32385 33284 32419
rect 33232 32376 33284 32385
rect 45928 32444 45980 32496
rect 46480 32419 46532 32428
rect 32404 32351 32456 32360
rect 29644 32308 29696 32317
rect 32404 32317 32413 32351
rect 32413 32317 32447 32351
rect 32447 32317 32456 32351
rect 32404 32308 32456 32317
rect 32588 32308 32640 32360
rect 22008 32240 22060 32292
rect 22652 32240 22704 32292
rect 26792 32240 26844 32292
rect 27528 32240 27580 32292
rect 27988 32240 28040 32292
rect 29460 32240 29512 32292
rect 29828 32240 29880 32292
rect 33600 32240 33652 32292
rect 34520 32240 34572 32292
rect 46480 32385 46489 32419
rect 46489 32385 46523 32419
rect 46523 32385 46532 32419
rect 46480 32376 46532 32385
rect 47492 32376 47544 32428
rect 37740 32351 37792 32360
rect 37740 32317 37749 32351
rect 37749 32317 37783 32351
rect 37783 32317 37792 32351
rect 37740 32308 37792 32317
rect 46204 32351 46256 32360
rect 13268 32215 13320 32224
rect 13268 32181 13277 32215
rect 13277 32181 13311 32215
rect 13311 32181 13320 32215
rect 13268 32172 13320 32181
rect 13728 32172 13780 32224
rect 23204 32215 23256 32224
rect 23204 32181 23213 32215
rect 23213 32181 23247 32215
rect 23247 32181 23256 32215
rect 23204 32172 23256 32181
rect 27804 32172 27856 32224
rect 28540 32172 28592 32224
rect 31024 32172 31076 32224
rect 31760 32172 31812 32224
rect 36176 32172 36228 32224
rect 46204 32317 46213 32351
rect 46213 32317 46247 32351
rect 46247 32317 46256 32351
rect 46204 32308 46256 32317
rect 46480 32172 46532 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2780 31968 2832 32020
rect 8300 31968 8352 32020
rect 9864 31968 9916 32020
rect 11704 31968 11756 32020
rect 12808 31968 12860 32020
rect 3056 31900 3108 31952
rect 25504 31968 25556 32020
rect 23572 31900 23624 31952
rect 9404 31875 9456 31884
rect 9404 31841 9413 31875
rect 9413 31841 9447 31875
rect 9447 31841 9456 31875
rect 9404 31832 9456 31841
rect 9772 31832 9824 31884
rect 9864 31875 9916 31884
rect 9864 31841 9873 31875
rect 9873 31841 9907 31875
rect 9907 31841 9916 31875
rect 9864 31832 9916 31841
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 3056 31764 3108 31816
rect 12900 31832 12952 31884
rect 15200 31832 15252 31884
rect 12624 31807 12676 31816
rect 12624 31773 12633 31807
rect 12633 31773 12667 31807
rect 12667 31773 12676 31807
rect 12624 31764 12676 31773
rect 16580 31764 16632 31816
rect 20812 31832 20864 31884
rect 20444 31764 20496 31816
rect 24768 31832 24820 31884
rect 22376 31764 22428 31816
rect 22652 31764 22704 31816
rect 23664 31764 23716 31816
rect 24676 31764 24728 31816
rect 27988 31943 28040 31952
rect 27988 31909 27997 31943
rect 27997 31909 28031 31943
rect 28031 31909 28040 31943
rect 27988 31900 28040 31909
rect 28080 31900 28132 31952
rect 28632 31900 28684 31952
rect 12532 31696 12584 31748
rect 2872 31671 2924 31680
rect 2872 31637 2881 31671
rect 2881 31637 2915 31671
rect 2915 31637 2924 31671
rect 2872 31628 2924 31637
rect 15384 31671 15436 31680
rect 15384 31637 15393 31671
rect 15393 31637 15427 31671
rect 15427 31637 15436 31671
rect 15384 31628 15436 31637
rect 20812 31628 20864 31680
rect 21916 31628 21968 31680
rect 22008 31628 22060 31680
rect 22192 31671 22244 31680
rect 22192 31637 22201 31671
rect 22201 31637 22235 31671
rect 22235 31637 22244 31671
rect 22192 31628 22244 31637
rect 24400 31628 24452 31680
rect 24492 31628 24544 31680
rect 25688 31807 25740 31816
rect 25688 31773 25697 31807
rect 25697 31773 25731 31807
rect 25731 31773 25740 31807
rect 25688 31764 25740 31773
rect 25964 31832 26016 31884
rect 26792 31764 26844 31816
rect 26976 31764 27028 31816
rect 27804 31807 27856 31816
rect 27804 31773 27813 31807
rect 27813 31773 27847 31807
rect 27847 31773 27856 31807
rect 27804 31764 27856 31773
rect 29092 31832 29144 31884
rect 25780 31696 25832 31748
rect 27068 31696 27120 31748
rect 30472 31764 30524 31816
rect 31208 31764 31260 31816
rect 31760 31807 31812 31816
rect 31760 31773 31769 31807
rect 31769 31773 31803 31807
rect 31803 31773 31812 31807
rect 31760 31764 31812 31773
rect 32680 31832 32732 31884
rect 32588 31807 32640 31816
rect 32588 31773 32595 31807
rect 32595 31773 32640 31807
rect 32588 31764 32640 31773
rect 32220 31696 32272 31748
rect 32772 31739 32824 31748
rect 32772 31705 32781 31739
rect 32781 31705 32815 31739
rect 32815 31705 32824 31739
rect 33416 31900 33468 31952
rect 33692 31832 33744 31884
rect 36176 31875 36228 31884
rect 36176 31841 36185 31875
rect 36185 31841 36219 31875
rect 36219 31841 36228 31875
rect 36176 31832 36228 31841
rect 36636 31832 36688 31884
rect 46296 31875 46348 31884
rect 46296 31841 46305 31875
rect 46305 31841 46339 31875
rect 46339 31841 46348 31875
rect 46296 31832 46348 31841
rect 46480 31875 46532 31884
rect 46480 31841 46489 31875
rect 46489 31841 46523 31875
rect 46523 31841 46532 31875
rect 46480 31832 46532 31841
rect 48136 31875 48188 31884
rect 48136 31841 48145 31875
rect 48145 31841 48179 31875
rect 48179 31841 48188 31875
rect 48136 31832 48188 31841
rect 34704 31807 34756 31816
rect 34704 31773 34713 31807
rect 34713 31773 34747 31807
rect 34747 31773 34756 31807
rect 34704 31764 34756 31773
rect 34796 31807 34848 31816
rect 34796 31773 34805 31807
rect 34805 31773 34839 31807
rect 34839 31773 34848 31807
rect 34796 31764 34848 31773
rect 32772 31696 32824 31705
rect 37464 31696 37516 31748
rect 32956 31628 33008 31680
rect 37556 31628 37608 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 9772 31467 9824 31476
rect 9772 31433 9781 31467
rect 9781 31433 9815 31467
rect 9815 31433 9824 31467
rect 9772 31424 9824 31433
rect 11520 31424 11572 31476
rect 14096 31424 14148 31476
rect 25504 31424 25556 31476
rect 26424 31424 26476 31476
rect 32588 31424 32640 31476
rect 37464 31424 37516 31476
rect 2872 31356 2924 31408
rect 20444 31356 20496 31408
rect 21824 31356 21876 31408
rect 24492 31399 24544 31408
rect 24492 31365 24501 31399
rect 24501 31365 24535 31399
rect 24535 31365 24544 31399
rect 24492 31356 24544 31365
rect 25964 31356 26016 31408
rect 26608 31356 26660 31408
rect 28448 31356 28500 31408
rect 29184 31356 29236 31408
rect 29368 31356 29420 31408
rect 30564 31356 30616 31408
rect 1952 31331 2004 31340
rect 1952 31297 1961 31331
rect 1961 31297 1995 31331
rect 1995 31297 2004 31331
rect 1952 31288 2004 31297
rect 9680 31331 9732 31340
rect 9680 31297 9689 31331
rect 9689 31297 9723 31331
rect 9723 31297 9732 31331
rect 9680 31288 9732 31297
rect 10968 31288 11020 31340
rect 15568 31288 15620 31340
rect 2964 31263 3016 31272
rect 2964 31229 2973 31263
rect 2973 31229 3007 31263
rect 3007 31229 3016 31263
rect 2964 31220 3016 31229
rect 13912 31263 13964 31272
rect 13912 31229 13921 31263
rect 13921 31229 13955 31263
rect 13955 31229 13964 31263
rect 13912 31220 13964 31229
rect 19156 31263 19208 31272
rect 19156 31229 19165 31263
rect 19165 31229 19199 31263
rect 19199 31229 19208 31263
rect 19156 31220 19208 31229
rect 20720 31220 20772 31272
rect 22008 31263 22060 31272
rect 22008 31229 22017 31263
rect 22017 31229 22051 31263
rect 22051 31229 22060 31263
rect 22008 31220 22060 31229
rect 22376 31220 22428 31272
rect 22560 31220 22612 31272
rect 26424 31288 26476 31340
rect 24216 31263 24268 31272
rect 24216 31229 24225 31263
rect 24225 31229 24259 31263
rect 24259 31229 24268 31263
rect 24216 31220 24268 31229
rect 24492 31220 24544 31272
rect 31116 31288 31168 31340
rect 31392 31288 31444 31340
rect 33692 31356 33744 31408
rect 34796 31356 34848 31408
rect 34704 31288 34756 31340
rect 36176 31288 36228 31340
rect 36636 31288 36688 31340
rect 37556 31356 37608 31408
rect 46112 31399 46164 31408
rect 46112 31365 46121 31399
rect 46121 31365 46155 31399
rect 46155 31365 46164 31399
rect 46112 31356 46164 31365
rect 27896 31220 27948 31272
rect 33140 31263 33192 31272
rect 33140 31229 33149 31263
rect 33149 31229 33183 31263
rect 33183 31229 33192 31263
rect 33140 31220 33192 31229
rect 33416 31263 33468 31272
rect 33416 31229 33425 31263
rect 33425 31229 33459 31263
rect 33459 31229 33468 31263
rect 33416 31220 33468 31229
rect 14648 31084 14700 31136
rect 16764 31084 16816 31136
rect 20904 31127 20956 31136
rect 20904 31093 20913 31127
rect 20913 31093 20947 31127
rect 20947 31093 20956 31127
rect 20904 31084 20956 31093
rect 21824 31084 21876 31136
rect 22468 31084 22520 31136
rect 25780 31084 25832 31136
rect 29092 31084 29144 31136
rect 37740 31220 37792 31272
rect 44180 31220 44232 31272
rect 47400 31356 47452 31408
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 15200 30923 15252 30932
rect 15200 30889 15209 30923
rect 15209 30889 15243 30923
rect 15243 30889 15252 30923
rect 15200 30880 15252 30889
rect 20720 30880 20772 30932
rect 22468 30880 22520 30932
rect 25688 30880 25740 30932
rect 26424 30923 26476 30932
rect 26424 30889 26433 30923
rect 26433 30889 26467 30923
rect 26467 30889 26476 30923
rect 26424 30880 26476 30889
rect 12900 30812 12952 30864
rect 14096 30855 14148 30864
rect 13268 30744 13320 30796
rect 14096 30821 14105 30855
rect 14105 30821 14139 30855
rect 14139 30821 14148 30855
rect 14096 30812 14148 30821
rect 10968 30719 11020 30728
rect 10968 30685 10977 30719
rect 10977 30685 11011 30719
rect 11011 30685 11020 30719
rect 10968 30676 11020 30685
rect 11704 30719 11756 30728
rect 11704 30685 11713 30719
rect 11713 30685 11747 30719
rect 11747 30685 11756 30719
rect 11704 30676 11756 30685
rect 13084 30676 13136 30728
rect 11060 30651 11112 30660
rect 11060 30617 11069 30651
rect 11069 30617 11103 30651
rect 11103 30617 11112 30651
rect 11060 30608 11112 30617
rect 12716 30651 12768 30660
rect 12716 30617 12725 30651
rect 12725 30617 12759 30651
rect 12759 30617 12768 30651
rect 13728 30676 13780 30728
rect 15384 30744 15436 30796
rect 19156 30744 19208 30796
rect 24216 30744 24268 30796
rect 25688 30744 25740 30796
rect 26056 30744 26108 30796
rect 15752 30719 15804 30728
rect 12716 30608 12768 30617
rect 13544 30608 13596 30660
rect 15752 30685 15761 30719
rect 15761 30685 15795 30719
rect 15795 30685 15804 30719
rect 15752 30676 15804 30685
rect 21824 30719 21876 30728
rect 21824 30685 21833 30719
rect 21833 30685 21867 30719
rect 21867 30685 21876 30719
rect 21824 30676 21876 30685
rect 21916 30719 21968 30728
rect 21916 30685 21925 30719
rect 21925 30685 21959 30719
rect 21959 30685 21968 30719
rect 21916 30676 21968 30685
rect 22376 30676 22428 30728
rect 16764 30608 16816 30660
rect 11796 30583 11848 30592
rect 11796 30549 11805 30583
rect 11805 30549 11839 30583
rect 11839 30549 11848 30583
rect 11796 30540 11848 30549
rect 12532 30540 12584 30592
rect 12900 30583 12952 30592
rect 12900 30549 12909 30583
rect 12909 30549 12943 30583
rect 12943 30549 12952 30583
rect 12900 30540 12952 30549
rect 13084 30583 13136 30592
rect 13084 30549 13093 30583
rect 13093 30549 13127 30583
rect 13127 30549 13136 30583
rect 13084 30540 13136 30549
rect 13268 30540 13320 30592
rect 14740 30540 14792 30592
rect 16672 30540 16724 30592
rect 17500 30583 17552 30592
rect 17500 30549 17509 30583
rect 17509 30549 17543 30583
rect 17543 30549 17552 30583
rect 17500 30540 17552 30549
rect 20812 30608 20864 30660
rect 21088 30608 21140 30660
rect 21732 30608 21784 30660
rect 25780 30676 25832 30728
rect 28632 30676 28684 30728
rect 30196 30676 30248 30728
rect 33232 30676 33284 30728
rect 24860 30608 24912 30660
rect 31300 30651 31352 30660
rect 31300 30617 31309 30651
rect 31309 30617 31343 30651
rect 31343 30617 31352 30651
rect 31300 30608 31352 30617
rect 33692 30608 33744 30660
rect 20996 30583 21048 30592
rect 20996 30549 21005 30583
rect 21005 30549 21039 30583
rect 21039 30549 21048 30583
rect 21456 30583 21508 30592
rect 20996 30540 21048 30549
rect 21456 30549 21465 30583
rect 21465 30549 21499 30583
rect 21499 30549 21508 30583
rect 21456 30540 21508 30549
rect 22652 30540 22704 30592
rect 24216 30540 24268 30592
rect 25044 30540 25096 30592
rect 28356 30583 28408 30592
rect 28356 30549 28365 30583
rect 28365 30549 28399 30583
rect 28399 30549 28408 30583
rect 28356 30540 28408 30549
rect 30380 30540 30432 30592
rect 31392 30583 31444 30592
rect 31392 30549 31401 30583
rect 31401 30549 31435 30583
rect 31435 30549 31444 30583
rect 31392 30540 31444 30549
rect 33324 30540 33376 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 13268 30379 13320 30388
rect 13268 30345 13277 30379
rect 13277 30345 13311 30379
rect 13311 30345 13320 30379
rect 13268 30336 13320 30345
rect 13912 30336 13964 30388
rect 15752 30336 15804 30388
rect 24492 30379 24544 30388
rect 24492 30345 24501 30379
rect 24501 30345 24535 30379
rect 24535 30345 24544 30379
rect 24492 30336 24544 30345
rect 25320 30336 25372 30388
rect 46848 30336 46900 30388
rect 11796 30311 11848 30320
rect 11796 30277 11805 30311
rect 11805 30277 11839 30311
rect 11839 30277 11848 30311
rect 11796 30268 11848 30277
rect 12440 30268 12492 30320
rect 14648 30268 14700 30320
rect 21088 30268 21140 30320
rect 11060 30200 11112 30252
rect 13084 30132 13136 30184
rect 16120 30200 16172 30252
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 22100 30243 22152 30252
rect 22100 30209 22109 30243
rect 22109 30209 22143 30243
rect 22143 30209 22152 30243
rect 22100 30200 22152 30209
rect 22284 30243 22336 30252
rect 22284 30209 22293 30243
rect 22293 30209 22327 30243
rect 22327 30209 22336 30243
rect 22284 30200 22336 30209
rect 22744 30200 22796 30252
rect 23020 30200 23072 30252
rect 26424 30268 26476 30320
rect 28356 30268 28408 30320
rect 25044 30200 25096 30252
rect 30380 30268 30432 30320
rect 33140 30268 33192 30320
rect 32496 30200 32548 30252
rect 33324 30243 33376 30252
rect 33324 30209 33333 30243
rect 33333 30209 33367 30243
rect 33367 30209 33376 30243
rect 33324 30200 33376 30209
rect 33508 30243 33560 30252
rect 33508 30209 33517 30243
rect 33517 30209 33551 30243
rect 33551 30209 33560 30243
rect 33508 30200 33560 30209
rect 33876 30243 33928 30252
rect 33876 30209 33885 30243
rect 33885 30209 33919 30243
rect 33919 30209 33928 30243
rect 33876 30200 33928 30209
rect 35348 30268 35400 30320
rect 14096 30064 14148 30116
rect 15200 30132 15252 30184
rect 20996 30175 21048 30184
rect 20996 30141 21005 30175
rect 21005 30141 21039 30175
rect 21039 30141 21048 30175
rect 22376 30175 22428 30184
rect 20996 30132 21048 30141
rect 22376 30141 22385 30175
rect 22385 30141 22419 30175
rect 22419 30141 22428 30175
rect 22376 30132 22428 30141
rect 23388 30132 23440 30184
rect 24952 30175 25004 30184
rect 24952 30141 24961 30175
rect 24961 30141 24995 30175
rect 24995 30141 25004 30175
rect 24952 30132 25004 30141
rect 27620 30175 27672 30184
rect 27620 30141 27629 30175
rect 27629 30141 27663 30175
rect 27663 30141 27672 30175
rect 27620 30132 27672 30141
rect 30656 30132 30708 30184
rect 31116 30132 31168 30184
rect 33232 30132 33284 30184
rect 33600 30175 33652 30184
rect 33600 30141 33609 30175
rect 33609 30141 33643 30175
rect 33643 30141 33652 30175
rect 33600 30132 33652 30141
rect 21732 30064 21784 30116
rect 24308 30107 24360 30116
rect 24308 30073 24317 30107
rect 24317 30073 24351 30107
rect 24351 30073 24360 30107
rect 24308 30064 24360 30073
rect 26240 30064 26292 30116
rect 28632 30064 28684 30116
rect 21272 30039 21324 30048
rect 21272 30005 21281 30039
rect 21281 30005 21315 30039
rect 21315 30005 21324 30039
rect 21272 29996 21324 30005
rect 24768 29996 24820 30048
rect 27068 29996 27120 30048
rect 27344 29996 27396 30048
rect 29092 30039 29144 30048
rect 29092 30005 29101 30039
rect 29101 30005 29135 30039
rect 29135 30005 29144 30039
rect 29092 29996 29144 30005
rect 32404 30064 32456 30116
rect 31576 30039 31628 30048
rect 31576 30005 31585 30039
rect 31585 30005 31619 30039
rect 31619 30005 31628 30039
rect 31576 29996 31628 30005
rect 44456 30064 44508 30116
rect 36268 30039 36320 30048
rect 36268 30005 36277 30039
rect 36277 30005 36311 30039
rect 36311 30005 36320 30039
rect 36268 29996 36320 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 11704 29792 11756 29844
rect 12440 29835 12492 29844
rect 12440 29801 12449 29835
rect 12449 29801 12483 29835
rect 12483 29801 12492 29835
rect 21456 29835 21508 29844
rect 12440 29792 12492 29801
rect 21456 29801 21465 29835
rect 21465 29801 21499 29835
rect 21499 29801 21508 29835
rect 21456 29792 21508 29801
rect 22468 29792 22520 29844
rect 22652 29835 22704 29844
rect 22652 29801 22661 29835
rect 22661 29801 22695 29835
rect 22695 29801 22704 29835
rect 22652 29792 22704 29801
rect 24952 29792 25004 29844
rect 26240 29792 26292 29844
rect 27620 29792 27672 29844
rect 22100 29724 22152 29776
rect 24308 29724 24360 29776
rect 29000 29835 29052 29844
rect 29000 29801 29009 29835
rect 29009 29801 29043 29835
rect 29043 29801 29052 29835
rect 30840 29835 30892 29844
rect 29000 29792 29052 29801
rect 30840 29801 30849 29835
rect 30849 29801 30883 29835
rect 30883 29801 30892 29835
rect 30840 29792 30892 29801
rect 31116 29792 31168 29844
rect 32496 29835 32548 29844
rect 32496 29801 32505 29835
rect 32505 29801 32539 29835
rect 32539 29801 32548 29835
rect 32496 29792 32548 29801
rect 33600 29792 33652 29844
rect 35348 29792 35400 29844
rect 36452 29792 36504 29844
rect 12716 29656 12768 29708
rect 11244 29588 11296 29640
rect 9128 29520 9180 29572
rect 12624 29588 12676 29640
rect 15568 29588 15620 29640
rect 16120 29656 16172 29708
rect 24952 29656 25004 29708
rect 25688 29699 25740 29708
rect 25688 29665 25697 29699
rect 25697 29665 25731 29699
rect 25731 29665 25740 29699
rect 25688 29656 25740 29665
rect 26056 29656 26108 29708
rect 28632 29699 28684 29708
rect 28632 29665 28641 29699
rect 28641 29665 28675 29699
rect 28675 29665 28684 29699
rect 28632 29656 28684 29665
rect 29092 29724 29144 29776
rect 13268 29520 13320 29572
rect 15936 29520 15988 29572
rect 17040 29520 17092 29572
rect 22192 29588 22244 29640
rect 23112 29588 23164 29640
rect 25780 29631 25832 29640
rect 23020 29520 23072 29572
rect 24676 29520 24728 29572
rect 25780 29597 25789 29631
rect 25789 29597 25823 29631
rect 25823 29597 25832 29631
rect 25780 29588 25832 29597
rect 27160 29631 27212 29640
rect 27160 29597 27169 29631
rect 27169 29597 27203 29631
rect 27203 29597 27212 29631
rect 27160 29588 27212 29597
rect 27252 29631 27304 29640
rect 27252 29597 27262 29631
rect 27262 29597 27296 29631
rect 27296 29597 27304 29631
rect 27252 29588 27304 29597
rect 28264 29588 28316 29640
rect 28816 29631 28868 29640
rect 28816 29597 28825 29631
rect 28825 29597 28859 29631
rect 28859 29597 28868 29631
rect 28816 29588 28868 29597
rect 46848 29724 46900 29776
rect 30380 29656 30432 29708
rect 31392 29656 31444 29708
rect 31576 29656 31628 29708
rect 30288 29588 30340 29640
rect 31024 29588 31076 29640
rect 32404 29631 32456 29640
rect 32404 29597 32413 29631
rect 32413 29597 32447 29631
rect 32447 29597 32456 29631
rect 32404 29588 32456 29597
rect 33416 29588 33468 29640
rect 33692 29588 33744 29640
rect 34428 29656 34480 29708
rect 36084 29699 36136 29708
rect 36084 29665 36093 29699
rect 36093 29665 36127 29699
rect 36127 29665 36136 29699
rect 36084 29656 36136 29665
rect 33968 29588 34020 29640
rect 36176 29631 36228 29640
rect 36176 29597 36185 29631
rect 36185 29597 36219 29631
rect 36219 29597 36228 29631
rect 36176 29588 36228 29597
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 47768 29588 47820 29640
rect 26148 29520 26200 29572
rect 27068 29520 27120 29572
rect 28080 29520 28132 29572
rect 28356 29520 28408 29572
rect 12440 29452 12492 29504
rect 18052 29452 18104 29504
rect 21548 29452 21600 29504
rect 25872 29452 25924 29504
rect 27252 29452 27304 29504
rect 30840 29452 30892 29504
rect 30932 29452 30984 29504
rect 31484 29452 31536 29504
rect 32404 29452 32456 29504
rect 33968 29452 34020 29504
rect 34428 29520 34480 29572
rect 36268 29520 36320 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 17040 29291 17092 29300
rect 17040 29257 17049 29291
rect 17049 29257 17083 29291
rect 17083 29257 17092 29291
rect 17040 29248 17092 29257
rect 1768 29180 1820 29232
rect 9036 29180 9088 29232
rect 9128 29155 9180 29164
rect 9128 29121 9137 29155
rect 9137 29121 9171 29155
rect 9171 29121 9180 29155
rect 9128 29112 9180 29121
rect 9772 29044 9824 29096
rect 12900 29180 12952 29232
rect 13452 29112 13504 29164
rect 14464 29155 14516 29164
rect 14464 29121 14473 29155
rect 14473 29121 14507 29155
rect 14507 29121 14516 29155
rect 14464 29112 14516 29121
rect 15476 29112 15528 29164
rect 18052 29180 18104 29232
rect 24308 29180 24360 29232
rect 15752 29112 15804 29164
rect 21272 29112 21324 29164
rect 21640 29112 21692 29164
rect 22560 29112 22612 29164
rect 27344 29248 27396 29300
rect 28816 29248 28868 29300
rect 30380 29248 30432 29300
rect 30656 29291 30708 29300
rect 30656 29257 30665 29291
rect 30665 29257 30699 29291
rect 30699 29257 30708 29291
rect 30656 29248 30708 29257
rect 29828 29180 29880 29232
rect 33968 29248 34020 29300
rect 24584 29155 24636 29164
rect 24584 29121 24593 29155
rect 24593 29121 24627 29155
rect 24627 29121 24636 29155
rect 24584 29112 24636 29121
rect 24676 29155 24728 29164
rect 24676 29121 24685 29155
rect 24685 29121 24719 29155
rect 24719 29121 24728 29155
rect 24676 29112 24728 29121
rect 14280 29087 14332 29096
rect 14280 29053 14289 29087
rect 14289 29053 14323 29087
rect 14323 29053 14332 29087
rect 14280 29044 14332 29053
rect 15200 29044 15252 29096
rect 15660 29087 15712 29096
rect 15660 29053 15669 29087
rect 15669 29053 15703 29087
rect 15703 29053 15712 29087
rect 15660 29044 15712 29053
rect 15936 29087 15988 29096
rect 15936 29053 15945 29087
rect 15945 29053 15979 29087
rect 15979 29053 15988 29087
rect 15936 29044 15988 29053
rect 18144 29087 18196 29096
rect 18144 29053 18153 29087
rect 18153 29053 18187 29087
rect 18187 29053 18196 29087
rect 18144 29044 18196 29053
rect 18328 29087 18380 29096
rect 18328 29053 18337 29087
rect 18337 29053 18371 29087
rect 18371 29053 18380 29087
rect 18328 29044 18380 29053
rect 25872 29155 25924 29164
rect 25872 29121 25881 29155
rect 25881 29121 25915 29155
rect 25915 29121 25924 29155
rect 25872 29112 25924 29121
rect 25964 29112 26016 29164
rect 27712 29155 27764 29164
rect 27712 29121 27721 29155
rect 27721 29121 27755 29155
rect 27755 29121 27764 29155
rect 27712 29112 27764 29121
rect 29000 29112 29052 29164
rect 29736 29112 29788 29164
rect 29920 29155 29972 29164
rect 29920 29121 29929 29155
rect 29929 29121 29963 29155
rect 29963 29121 29972 29155
rect 29920 29112 29972 29121
rect 30380 29112 30432 29164
rect 27068 29044 27120 29096
rect 29460 29044 29512 29096
rect 30840 29112 30892 29164
rect 31024 29112 31076 29164
rect 31392 29155 31444 29164
rect 31392 29121 31401 29155
rect 31401 29121 31435 29155
rect 31435 29121 31444 29155
rect 31392 29112 31444 29121
rect 31576 29112 31628 29164
rect 32588 29155 32640 29164
rect 32588 29121 32597 29155
rect 32597 29121 32631 29155
rect 32631 29121 32640 29155
rect 32588 29112 32640 29121
rect 12624 28908 12676 28960
rect 14648 28908 14700 28960
rect 22100 28908 22152 28960
rect 24768 28908 24820 28960
rect 25136 28951 25188 28960
rect 25136 28917 25145 28951
rect 25145 28917 25179 28951
rect 25179 28917 25188 28951
rect 25136 28908 25188 28917
rect 25688 28951 25740 28960
rect 25688 28917 25697 28951
rect 25697 28917 25731 28951
rect 25731 28917 25740 28951
rect 25688 28908 25740 28917
rect 28908 28908 28960 28960
rect 33232 28976 33284 29028
rect 33876 29112 33928 29164
rect 34428 29155 34480 29164
rect 34428 29121 34437 29155
rect 34437 29121 34471 29155
rect 34471 29121 34480 29155
rect 34428 29112 34480 29121
rect 33508 28976 33560 29028
rect 33692 29044 33744 29096
rect 36084 29112 36136 29164
rect 34612 28976 34664 29028
rect 31208 28908 31260 28960
rect 31576 28951 31628 28960
rect 31576 28917 31585 28951
rect 31585 28917 31619 28951
rect 31619 28917 31628 28951
rect 31576 28908 31628 28917
rect 32312 28951 32364 28960
rect 32312 28917 32321 28951
rect 32321 28917 32355 28951
rect 32355 28917 32364 28951
rect 32312 28908 32364 28917
rect 33600 28908 33652 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 9772 28747 9824 28756
rect 9772 28713 9781 28747
rect 9781 28713 9815 28747
rect 9815 28713 9824 28747
rect 9772 28704 9824 28713
rect 13360 28704 13412 28756
rect 23480 28704 23532 28756
rect 11244 28636 11296 28688
rect 14648 28636 14700 28688
rect 11796 28568 11848 28620
rect 14556 28568 14608 28620
rect 23020 28636 23072 28688
rect 25688 28704 25740 28756
rect 26148 28747 26200 28756
rect 26148 28713 26157 28747
rect 26157 28713 26191 28747
rect 26191 28713 26200 28747
rect 26148 28704 26200 28713
rect 27804 28704 27856 28756
rect 29736 28747 29788 28756
rect 29736 28713 29745 28747
rect 29745 28713 29779 28747
rect 29779 28713 29788 28747
rect 29736 28704 29788 28713
rect 29828 28704 29880 28756
rect 32588 28704 32640 28756
rect 36084 28704 36136 28756
rect 26516 28636 26568 28688
rect 9680 28543 9732 28552
rect 9680 28509 9689 28543
rect 9689 28509 9723 28543
rect 9723 28509 9732 28543
rect 9680 28500 9732 28509
rect 12440 28500 12492 28552
rect 13544 28500 13596 28552
rect 15200 28500 15252 28552
rect 15384 28543 15436 28552
rect 15384 28509 15393 28543
rect 15393 28509 15427 28543
rect 15427 28509 15436 28543
rect 15384 28500 15436 28509
rect 16120 28543 16172 28552
rect 16120 28509 16129 28543
rect 16129 28509 16163 28543
rect 16163 28509 16172 28543
rect 16120 28500 16172 28509
rect 19340 28543 19392 28552
rect 19340 28509 19349 28543
rect 19349 28509 19383 28543
rect 19383 28509 19392 28543
rect 19340 28500 19392 28509
rect 21088 28500 21140 28552
rect 22100 28568 22152 28620
rect 25136 28568 25188 28620
rect 27068 28568 27120 28620
rect 30288 28636 30340 28688
rect 31024 28636 31076 28688
rect 32312 28636 32364 28688
rect 24400 28543 24452 28552
rect 13360 28475 13412 28484
rect 13360 28441 13369 28475
rect 13369 28441 13403 28475
rect 13403 28441 13412 28475
rect 13360 28432 13412 28441
rect 13912 28432 13964 28484
rect 14740 28432 14792 28484
rect 13452 28407 13504 28416
rect 13452 28373 13461 28407
rect 13461 28373 13495 28407
rect 13495 28373 13504 28407
rect 13452 28364 13504 28373
rect 14280 28407 14332 28416
rect 14280 28373 14289 28407
rect 14289 28373 14323 28407
rect 14323 28373 14332 28407
rect 14280 28364 14332 28373
rect 14464 28407 14516 28416
rect 14464 28373 14473 28407
rect 14473 28373 14507 28407
rect 14507 28373 14516 28407
rect 15016 28432 15068 28484
rect 14464 28364 14516 28373
rect 15292 28407 15344 28416
rect 15292 28373 15301 28407
rect 15301 28373 15335 28407
rect 15335 28373 15344 28407
rect 15292 28364 15344 28373
rect 15568 28364 15620 28416
rect 16672 28364 16724 28416
rect 20628 28432 20680 28484
rect 21180 28432 21232 28484
rect 21824 28475 21876 28484
rect 21824 28441 21833 28475
rect 21833 28441 21867 28475
rect 21867 28441 21876 28475
rect 21824 28432 21876 28441
rect 20996 28364 21048 28416
rect 21272 28364 21324 28416
rect 22008 28364 22060 28416
rect 22284 28364 22336 28416
rect 24400 28509 24409 28543
rect 24409 28509 24443 28543
rect 24443 28509 24452 28543
rect 24400 28500 24452 28509
rect 27252 28543 27304 28552
rect 27252 28509 27261 28543
rect 27261 28509 27295 28543
rect 27295 28509 27304 28543
rect 27252 28500 27304 28509
rect 24768 28432 24820 28484
rect 25964 28432 26016 28484
rect 26240 28432 26292 28484
rect 26976 28364 27028 28416
rect 27252 28364 27304 28416
rect 31208 28568 31260 28620
rect 28632 28500 28684 28552
rect 28448 28432 28500 28484
rect 31392 28500 31444 28552
rect 31760 28500 31812 28552
rect 34428 28568 34480 28620
rect 34612 28568 34664 28620
rect 30288 28432 30340 28484
rect 33416 28543 33468 28552
rect 33416 28509 33425 28543
rect 33425 28509 33459 28543
rect 33459 28509 33468 28543
rect 33416 28500 33468 28509
rect 34704 28500 34756 28552
rect 46940 28500 46992 28552
rect 33692 28432 33744 28484
rect 36084 28432 36136 28484
rect 29736 28364 29788 28416
rect 32496 28364 32548 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 10968 28092 11020 28144
rect 11796 28135 11848 28144
rect 11796 28101 11805 28135
rect 11805 28101 11839 28135
rect 11839 28101 11848 28135
rect 11796 28092 11848 28101
rect 12440 28092 12492 28144
rect 13544 28135 13596 28144
rect 13544 28101 13553 28135
rect 13553 28101 13587 28135
rect 13587 28101 13596 28135
rect 13544 28092 13596 28101
rect 15568 28160 15620 28212
rect 18236 28160 18288 28212
rect 20628 28160 20680 28212
rect 21180 28203 21232 28212
rect 21180 28169 21189 28203
rect 21189 28169 21223 28203
rect 21223 28169 21232 28203
rect 21180 28160 21232 28169
rect 21824 28160 21876 28212
rect 24768 28160 24820 28212
rect 24860 28160 24912 28212
rect 27160 28160 27212 28212
rect 27436 28160 27488 28212
rect 17960 28092 18012 28144
rect 14740 28024 14792 28076
rect 15016 28024 15068 28076
rect 15476 28067 15528 28076
rect 15476 28033 15485 28067
rect 15485 28033 15519 28067
rect 15519 28033 15528 28067
rect 15476 28024 15528 28033
rect 15660 28024 15712 28076
rect 16672 28067 16724 28076
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 22100 28092 22152 28144
rect 24400 28092 24452 28144
rect 24952 28092 25004 28144
rect 28908 28092 28960 28144
rect 31300 28092 31352 28144
rect 21272 28067 21324 28076
rect 18144 27956 18196 28008
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 21272 28024 21324 28033
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 20996 27956 21048 28008
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22284 28024 22336 28033
rect 23480 28024 23532 28076
rect 26240 28067 26292 28076
rect 26240 28033 26249 28067
rect 26249 28033 26283 28067
rect 26283 28033 26292 28067
rect 26240 28024 26292 28033
rect 27436 28067 27488 28076
rect 21272 27888 21324 27940
rect 20628 27820 20680 27872
rect 25872 27820 25924 27872
rect 27436 28033 27445 28067
rect 27445 28033 27479 28067
rect 27479 28033 27488 28067
rect 27436 28024 27488 28033
rect 28356 28067 28408 28076
rect 28356 28033 28371 28067
rect 28371 28033 28405 28067
rect 28405 28033 28408 28067
rect 28356 28024 28408 28033
rect 27804 27956 27856 28008
rect 29276 28024 29328 28076
rect 29920 28024 29972 28076
rect 32128 28024 32180 28076
rect 32496 28067 32548 28076
rect 32496 28033 32505 28067
rect 32505 28033 32539 28067
rect 32539 28033 32548 28067
rect 32496 28024 32548 28033
rect 33968 28160 34020 28212
rect 34796 28160 34848 28212
rect 36084 28160 36136 28212
rect 34520 28092 34572 28144
rect 34428 28067 34480 28076
rect 34428 28033 34437 28067
rect 34437 28033 34471 28067
rect 34471 28033 34480 28067
rect 34428 28024 34480 28033
rect 45652 28024 45704 28076
rect 47584 28067 47636 28076
rect 47584 28033 47593 28067
rect 47593 28033 47627 28067
rect 47627 28033 47636 28067
rect 47584 28024 47636 28033
rect 30564 27956 30616 28008
rect 47400 27956 47452 28008
rect 28540 27888 28592 27940
rect 32036 27888 32088 27940
rect 32404 27888 32456 27940
rect 34336 27888 34388 27940
rect 36084 27888 36136 27940
rect 27620 27820 27672 27872
rect 27988 27820 28040 27872
rect 31852 27820 31904 27872
rect 31944 27820 31996 27872
rect 33324 27820 33376 27872
rect 34428 27820 34480 27872
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3332 27616 3384 27668
rect 21640 27659 21692 27668
rect 12440 27548 12492 27600
rect 11520 27480 11572 27532
rect 21640 27625 21649 27659
rect 21649 27625 21683 27659
rect 21683 27625 21692 27659
rect 21640 27616 21692 27625
rect 22284 27616 22336 27668
rect 24768 27616 24820 27668
rect 28080 27616 28132 27668
rect 18328 27548 18380 27600
rect 19248 27548 19300 27600
rect 25780 27548 25832 27600
rect 25964 27591 26016 27600
rect 25964 27557 25973 27591
rect 25973 27557 26007 27591
rect 26007 27557 26016 27591
rect 25964 27548 26016 27557
rect 26332 27548 26384 27600
rect 26976 27548 27028 27600
rect 27252 27591 27304 27600
rect 27252 27557 27261 27591
rect 27261 27557 27295 27591
rect 27295 27557 27304 27591
rect 27252 27548 27304 27557
rect 27436 27548 27488 27600
rect 28540 27616 28592 27668
rect 30564 27616 30616 27668
rect 30288 27548 30340 27600
rect 30380 27548 30432 27600
rect 31852 27616 31904 27668
rect 33324 27616 33376 27668
rect 36452 27591 36504 27600
rect 36452 27557 36461 27591
rect 36461 27557 36495 27591
rect 36495 27557 36504 27591
rect 36452 27548 36504 27557
rect 22560 27523 22612 27532
rect 12532 27412 12584 27464
rect 13820 27412 13872 27464
rect 14096 27455 14148 27464
rect 14096 27421 14105 27455
rect 14105 27421 14139 27455
rect 14139 27421 14148 27455
rect 14096 27412 14148 27421
rect 17592 27412 17644 27464
rect 21272 27412 21324 27464
rect 21640 27412 21692 27464
rect 21916 27412 21968 27464
rect 22560 27489 22569 27523
rect 22569 27489 22603 27523
rect 22603 27489 22612 27523
rect 22560 27480 22612 27489
rect 22468 27455 22520 27464
rect 22468 27421 22477 27455
rect 22477 27421 22511 27455
rect 22511 27421 22520 27455
rect 22468 27412 22520 27421
rect 24860 27455 24912 27464
rect 24860 27421 24869 27455
rect 24869 27421 24903 27455
rect 24903 27421 24912 27455
rect 24860 27412 24912 27421
rect 27344 27480 27396 27532
rect 27068 27455 27120 27464
rect 27068 27421 27077 27455
rect 27077 27421 27111 27455
rect 27111 27421 27120 27455
rect 27068 27412 27120 27421
rect 29828 27480 29880 27532
rect 33416 27480 33468 27532
rect 34704 27523 34756 27532
rect 34704 27489 34713 27523
rect 34713 27489 34747 27523
rect 34747 27489 34756 27523
rect 34704 27480 34756 27489
rect 46940 27548 46992 27600
rect 47676 27480 47728 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 29368 27412 29420 27464
rect 29552 27412 29604 27464
rect 9772 27344 9824 27396
rect 7564 27276 7616 27328
rect 20812 27387 20864 27396
rect 20812 27353 20821 27387
rect 20821 27353 20855 27387
rect 20855 27353 20864 27387
rect 20812 27344 20864 27353
rect 14372 27276 14424 27328
rect 15476 27276 15528 27328
rect 30932 27412 30984 27464
rect 31208 27455 31260 27464
rect 31208 27421 31217 27455
rect 31217 27421 31251 27455
rect 31251 27421 31260 27455
rect 31208 27412 31260 27421
rect 31944 27455 31996 27464
rect 31944 27421 31953 27455
rect 31953 27421 31987 27455
rect 31987 27421 31996 27455
rect 31944 27412 31996 27421
rect 31484 27344 31536 27396
rect 31760 27344 31812 27396
rect 32220 27455 32272 27464
rect 32220 27421 32229 27455
rect 32229 27421 32263 27455
rect 32263 27421 32272 27455
rect 32220 27412 32272 27421
rect 32496 27412 32548 27464
rect 36084 27412 36136 27464
rect 45652 27455 45704 27464
rect 45652 27421 45661 27455
rect 45661 27421 45695 27455
rect 45695 27421 45704 27455
rect 45652 27412 45704 27421
rect 22836 27319 22888 27328
rect 22836 27285 22845 27319
rect 22845 27285 22879 27319
rect 22879 27285 22888 27319
rect 22836 27276 22888 27285
rect 24952 27319 25004 27328
rect 24952 27285 24961 27319
rect 24961 27285 24995 27319
rect 24995 27285 25004 27319
rect 24952 27276 25004 27285
rect 27160 27276 27212 27328
rect 32312 27387 32364 27396
rect 32312 27353 32321 27387
rect 32321 27353 32355 27387
rect 32355 27353 32364 27387
rect 32312 27344 32364 27353
rect 32772 27344 32824 27396
rect 45744 27319 45796 27328
rect 45744 27285 45753 27319
rect 45753 27285 45787 27319
rect 45787 27285 45796 27319
rect 45744 27276 45796 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9772 27115 9824 27124
rect 9772 27081 9781 27115
rect 9781 27081 9815 27115
rect 9815 27081 9824 27115
rect 9772 27072 9824 27081
rect 14464 27072 14516 27124
rect 14740 27072 14792 27124
rect 11888 27004 11940 27056
rect 14096 27004 14148 27056
rect 15568 27072 15620 27124
rect 17960 27072 18012 27124
rect 9680 26979 9732 26988
rect 9680 26945 9689 26979
rect 9689 26945 9723 26979
rect 9723 26945 9732 26979
rect 9680 26936 9732 26945
rect 10784 26979 10836 26988
rect 10784 26945 10793 26979
rect 10793 26945 10827 26979
rect 10827 26945 10836 26979
rect 10784 26936 10836 26945
rect 10968 26936 11020 26988
rect 14556 26936 14608 26988
rect 15384 26936 15436 26988
rect 17408 26936 17460 26988
rect 17960 26979 18012 26988
rect 17960 26945 17969 26979
rect 17969 26945 18003 26979
rect 18003 26945 18012 26979
rect 17960 26936 18012 26945
rect 21180 27004 21232 27056
rect 21088 26979 21140 26988
rect 21088 26945 21097 26979
rect 21097 26945 21131 26979
rect 21131 26945 21140 26979
rect 21088 26936 21140 26945
rect 22008 26979 22060 26988
rect 22008 26945 22017 26979
rect 22017 26945 22051 26979
rect 22051 26945 22060 26979
rect 22008 26936 22060 26945
rect 22192 26979 22244 26988
rect 22192 26945 22201 26979
rect 22201 26945 22235 26979
rect 22235 26945 22244 26979
rect 22192 26936 22244 26945
rect 11060 26800 11112 26852
rect 14832 26868 14884 26920
rect 18144 26911 18196 26920
rect 18144 26877 18153 26911
rect 18153 26877 18187 26911
rect 18187 26877 18196 26911
rect 18144 26868 18196 26877
rect 20260 26868 20312 26920
rect 21456 26868 21508 26920
rect 13820 26800 13872 26852
rect 17592 26800 17644 26852
rect 21088 26800 21140 26852
rect 22744 26868 22796 26920
rect 25780 27004 25832 27056
rect 27160 27004 27212 27056
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 26056 26936 26108 26988
rect 24860 26868 24912 26920
rect 31760 27072 31812 27124
rect 36452 27072 36504 27124
rect 46572 27115 46624 27124
rect 46572 27081 46581 27115
rect 46581 27081 46615 27115
rect 46615 27081 46624 27115
rect 46572 27072 46624 27081
rect 29184 27004 29236 27056
rect 32864 27004 32916 27056
rect 29368 26979 29420 26988
rect 29368 26945 29377 26979
rect 29377 26945 29411 26979
rect 29411 26945 29420 26979
rect 29368 26936 29420 26945
rect 29000 26868 29052 26920
rect 29184 26911 29236 26920
rect 29184 26877 29193 26911
rect 29193 26877 29227 26911
rect 29227 26877 29236 26911
rect 29184 26868 29236 26877
rect 22836 26800 22888 26852
rect 24676 26800 24728 26852
rect 26148 26800 26200 26852
rect 31024 26936 31076 26988
rect 45652 26936 45704 26988
rect 29828 26868 29880 26920
rect 31852 26868 31904 26920
rect 33048 26868 33100 26920
rect 46388 26868 46440 26920
rect 29552 26800 29604 26852
rect 30472 26800 30524 26852
rect 32772 26800 32824 26852
rect 13084 26732 13136 26784
rect 15292 26775 15344 26784
rect 15292 26741 15301 26775
rect 15301 26741 15335 26775
rect 15335 26741 15344 26775
rect 15292 26732 15344 26741
rect 19432 26732 19484 26784
rect 20720 26732 20772 26784
rect 20996 26732 21048 26784
rect 25136 26732 25188 26784
rect 26056 26732 26108 26784
rect 27896 26732 27948 26784
rect 28356 26775 28408 26784
rect 28356 26741 28365 26775
rect 28365 26741 28399 26775
rect 28399 26741 28408 26775
rect 28356 26732 28408 26741
rect 28540 26775 28592 26784
rect 28540 26741 28549 26775
rect 28549 26741 28583 26775
rect 28583 26741 28592 26775
rect 28540 26732 28592 26741
rect 30840 26732 30892 26784
rect 46664 26732 46716 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 11060 26571 11112 26580
rect 11060 26537 11069 26571
rect 11069 26537 11103 26571
rect 11103 26537 11112 26571
rect 11060 26528 11112 26537
rect 11888 26571 11940 26580
rect 11888 26537 11897 26571
rect 11897 26537 11931 26571
rect 11931 26537 11940 26571
rect 11888 26528 11940 26537
rect 15384 26528 15436 26580
rect 18144 26528 18196 26580
rect 20996 26528 21048 26580
rect 21088 26528 21140 26580
rect 21456 26528 21508 26580
rect 20720 26460 20772 26512
rect 11060 26367 11112 26376
rect 11060 26333 11069 26367
rect 11069 26333 11103 26367
rect 11103 26333 11112 26367
rect 11060 26324 11112 26333
rect 11244 26367 11296 26376
rect 11244 26333 11253 26367
rect 11253 26333 11287 26367
rect 11287 26333 11296 26367
rect 11244 26324 11296 26333
rect 12532 26324 12584 26376
rect 13452 26324 13504 26376
rect 14924 26324 14976 26376
rect 15660 26367 15712 26376
rect 15660 26333 15669 26367
rect 15669 26333 15703 26367
rect 15703 26333 15712 26367
rect 15660 26324 15712 26333
rect 17592 26324 17644 26376
rect 19340 26392 19392 26444
rect 20076 26392 20128 26444
rect 22468 26528 22520 26580
rect 24216 26528 24268 26580
rect 26516 26571 26568 26580
rect 22100 26460 22152 26512
rect 22284 26435 22336 26444
rect 22284 26401 22293 26435
rect 22293 26401 22327 26435
rect 22327 26401 22336 26435
rect 22284 26392 22336 26401
rect 14832 26299 14884 26308
rect 14832 26265 14841 26299
rect 14841 26265 14875 26299
rect 14875 26265 14884 26299
rect 14832 26256 14884 26265
rect 15568 26256 15620 26308
rect 15936 26299 15988 26308
rect 15936 26265 15945 26299
rect 15945 26265 15979 26299
rect 15979 26265 15988 26299
rect 15936 26256 15988 26265
rect 18788 26256 18840 26308
rect 14556 26188 14608 26240
rect 20720 26256 20772 26308
rect 21640 26256 21692 26308
rect 25228 26460 25280 26512
rect 25320 26460 25372 26512
rect 26516 26537 26525 26571
rect 26525 26537 26559 26571
rect 26559 26537 26568 26571
rect 26516 26528 26568 26537
rect 27344 26528 27396 26580
rect 29828 26528 29880 26580
rect 45468 26528 45520 26580
rect 45652 26571 45704 26580
rect 45652 26537 45661 26571
rect 45661 26537 45695 26571
rect 45695 26537 45704 26571
rect 45652 26528 45704 26537
rect 27068 26460 27120 26512
rect 27804 26460 27856 26512
rect 28724 26460 28776 26512
rect 30288 26460 30340 26512
rect 31944 26460 31996 26512
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 27160 26324 27212 26376
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 27620 26324 27672 26376
rect 30472 26392 30524 26444
rect 28540 26324 28592 26376
rect 32128 26392 32180 26444
rect 33324 26392 33376 26444
rect 31852 26367 31904 26376
rect 31852 26333 31861 26367
rect 31861 26333 31895 26367
rect 31895 26333 31904 26367
rect 31852 26324 31904 26333
rect 23756 26256 23808 26308
rect 25044 26256 25096 26308
rect 21456 26188 21508 26240
rect 23296 26188 23348 26240
rect 25412 26188 25464 26240
rect 26516 26188 26568 26240
rect 28632 26256 28684 26308
rect 32588 26367 32640 26376
rect 32588 26333 32597 26367
rect 32597 26333 32631 26367
rect 32631 26333 32640 26367
rect 32772 26367 32824 26376
rect 32588 26324 32640 26333
rect 32772 26333 32781 26367
rect 32781 26333 32815 26367
rect 32815 26333 32824 26367
rect 32772 26324 32824 26333
rect 32864 26367 32916 26376
rect 32864 26333 32873 26367
rect 32873 26333 32907 26367
rect 32907 26333 32916 26367
rect 47584 26460 47636 26512
rect 40132 26392 40184 26444
rect 32864 26324 32916 26333
rect 33508 26324 33560 26376
rect 33968 26367 34020 26376
rect 33232 26256 33284 26308
rect 33968 26333 33977 26367
rect 33977 26333 34011 26367
rect 34011 26333 34020 26367
rect 33968 26324 34020 26333
rect 45652 26392 45704 26444
rect 43996 26324 44048 26376
rect 45468 26367 45520 26376
rect 34152 26299 34204 26308
rect 34152 26265 34161 26299
rect 34161 26265 34195 26299
rect 34195 26265 34204 26299
rect 34152 26256 34204 26265
rect 45468 26333 45477 26367
rect 45477 26333 45511 26367
rect 45511 26333 45520 26367
rect 45468 26324 45520 26333
rect 47308 26392 47360 26444
rect 46020 26324 46072 26376
rect 47676 26256 47728 26308
rect 48136 26299 48188 26308
rect 48136 26265 48145 26299
rect 48145 26265 48179 26299
rect 48179 26265 48188 26299
rect 48136 26256 48188 26265
rect 30932 26188 30984 26240
rect 31392 26231 31444 26240
rect 31392 26197 31401 26231
rect 31401 26197 31435 26231
rect 31435 26197 31444 26231
rect 31392 26188 31444 26197
rect 31484 26188 31536 26240
rect 36544 26188 36596 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2320 25984 2372 26036
rect 11520 25959 11572 25968
rect 11520 25925 11529 25959
rect 11529 25925 11563 25959
rect 11563 25925 11572 25959
rect 13084 25959 13136 25968
rect 11520 25916 11572 25925
rect 13084 25925 13093 25959
rect 13093 25925 13127 25959
rect 13127 25925 13136 25959
rect 13084 25916 13136 25925
rect 14832 25984 14884 26036
rect 15200 25984 15252 26036
rect 15476 25984 15528 26036
rect 15660 25984 15712 26036
rect 17408 25984 17460 26036
rect 18788 26027 18840 26036
rect 11428 25848 11480 25900
rect 12072 25848 12124 25900
rect 13176 25848 13228 25900
rect 10784 25780 10836 25832
rect 14648 25848 14700 25900
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 15568 25848 15620 25900
rect 16120 25848 16172 25900
rect 9680 25712 9732 25764
rect 9864 25644 9916 25696
rect 11060 25712 11112 25764
rect 14372 25780 14424 25832
rect 15016 25712 15068 25764
rect 18788 25993 18797 26027
rect 18797 25993 18831 26027
rect 18831 25993 18840 26027
rect 18788 25984 18840 25993
rect 20720 26027 20772 26036
rect 20720 25993 20729 26027
rect 20729 25993 20763 26027
rect 20763 25993 20772 26027
rect 20720 25984 20772 25993
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 22192 25848 22244 25900
rect 23296 25712 23348 25764
rect 13268 25687 13320 25696
rect 13268 25653 13277 25687
rect 13277 25653 13311 25687
rect 13311 25653 13320 25687
rect 13268 25644 13320 25653
rect 17408 25644 17460 25696
rect 18144 25687 18196 25696
rect 18144 25653 18153 25687
rect 18153 25653 18187 25687
rect 18187 25653 18196 25687
rect 18144 25644 18196 25653
rect 22376 25644 22428 25696
rect 26056 25984 26108 26036
rect 26608 25984 26660 26036
rect 23756 25916 23808 25968
rect 28540 25984 28592 26036
rect 31944 25984 31996 26036
rect 32036 25984 32088 26036
rect 23848 25891 23900 25900
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 24860 25891 24912 25900
rect 24860 25857 24869 25891
rect 24869 25857 24903 25891
rect 24903 25857 24912 25891
rect 24860 25848 24912 25857
rect 25044 25891 25096 25900
rect 25044 25857 25053 25891
rect 25053 25857 25087 25891
rect 25087 25857 25096 25891
rect 25044 25848 25096 25857
rect 27896 25916 27948 25968
rect 31484 25916 31536 25968
rect 26792 25848 26844 25900
rect 27436 25823 27488 25832
rect 27436 25789 27445 25823
rect 27445 25789 27479 25823
rect 27479 25789 27488 25823
rect 27436 25780 27488 25789
rect 27620 25823 27672 25832
rect 27620 25789 27629 25823
rect 27629 25789 27663 25823
rect 27663 25789 27672 25823
rect 27620 25780 27672 25789
rect 28448 25848 28500 25900
rect 28632 25891 28684 25900
rect 28632 25857 28641 25891
rect 28641 25857 28675 25891
rect 28675 25857 28684 25891
rect 28632 25848 28684 25857
rect 29552 25891 29604 25900
rect 29552 25857 29561 25891
rect 29561 25857 29595 25891
rect 29595 25857 29604 25891
rect 29552 25848 29604 25857
rect 30840 25891 30892 25900
rect 30840 25857 30849 25891
rect 30849 25857 30883 25891
rect 30883 25857 30892 25891
rect 30840 25848 30892 25857
rect 30932 25891 30984 25900
rect 30932 25857 30941 25891
rect 30941 25857 30975 25891
rect 30975 25857 30984 25891
rect 31208 25891 31260 25900
rect 30932 25848 30984 25857
rect 31208 25857 31217 25891
rect 31217 25857 31251 25891
rect 31251 25857 31260 25891
rect 31208 25848 31260 25857
rect 32864 25916 32916 25968
rect 36544 25984 36596 26036
rect 45836 25984 45888 26036
rect 33876 25848 33928 25900
rect 34704 25916 34756 25968
rect 35348 25916 35400 25968
rect 45744 25916 45796 25968
rect 45928 25916 45980 25968
rect 30104 25780 30156 25832
rect 32772 25780 32824 25832
rect 34612 25823 34664 25832
rect 25320 25712 25372 25764
rect 26608 25712 26660 25764
rect 32128 25712 32180 25764
rect 34612 25789 34621 25823
rect 34621 25789 34655 25823
rect 34655 25789 34664 25823
rect 34612 25780 34664 25789
rect 45192 25823 45244 25832
rect 45192 25789 45201 25823
rect 45201 25789 45235 25823
rect 45235 25789 45244 25823
rect 45192 25780 45244 25789
rect 46848 25823 46900 25832
rect 46848 25789 46857 25823
rect 46857 25789 46891 25823
rect 46891 25789 46900 25823
rect 46848 25780 46900 25789
rect 25872 25644 25924 25696
rect 28356 25687 28408 25696
rect 28356 25653 28365 25687
rect 28365 25653 28399 25687
rect 28399 25653 28408 25687
rect 28356 25644 28408 25653
rect 31300 25644 31352 25696
rect 31484 25644 31536 25696
rect 33784 25644 33836 25696
rect 36084 25687 36136 25696
rect 36084 25653 36093 25687
rect 36093 25653 36127 25687
rect 36127 25653 36136 25687
rect 36084 25644 36136 25653
rect 46296 25644 46348 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 11428 25440 11480 25492
rect 13268 25440 13320 25492
rect 14372 25440 14424 25492
rect 15568 25440 15620 25492
rect 15936 25440 15988 25492
rect 17592 25483 17644 25492
rect 17592 25449 17601 25483
rect 17601 25449 17635 25483
rect 17635 25449 17644 25483
rect 17592 25440 17644 25449
rect 23756 25440 23808 25492
rect 26608 25483 26660 25492
rect 26608 25449 26617 25483
rect 26617 25449 26651 25483
rect 26651 25449 26660 25483
rect 26608 25440 26660 25449
rect 28080 25440 28132 25492
rect 29000 25440 29052 25492
rect 31208 25440 31260 25492
rect 31392 25483 31444 25492
rect 31392 25449 31401 25483
rect 31401 25449 31435 25483
rect 31435 25449 31444 25483
rect 31392 25440 31444 25449
rect 31852 25440 31904 25492
rect 32864 25483 32916 25492
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 12532 25236 12584 25288
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 10140 25211 10192 25220
rect 10140 25177 10149 25211
rect 10149 25177 10183 25211
rect 10183 25177 10192 25211
rect 10140 25168 10192 25177
rect 15108 25304 15160 25356
rect 19248 25304 19300 25356
rect 22376 25347 22428 25356
rect 22376 25313 22385 25347
rect 22385 25313 22419 25347
rect 22419 25313 22428 25347
rect 22376 25304 22428 25313
rect 29736 25372 29788 25424
rect 32864 25449 32873 25483
rect 32873 25449 32907 25483
rect 32907 25449 32916 25483
rect 32864 25440 32916 25449
rect 34612 25440 34664 25492
rect 35348 25440 35400 25492
rect 46020 25440 46072 25492
rect 1952 25143 2004 25152
rect 1952 25109 1961 25143
rect 1961 25109 1995 25143
rect 1995 25109 2004 25143
rect 1952 25100 2004 25109
rect 11520 25100 11572 25152
rect 13176 25100 13228 25152
rect 13728 25100 13780 25152
rect 15292 25236 15344 25288
rect 15844 25279 15896 25288
rect 15844 25245 15853 25279
rect 15853 25245 15887 25279
rect 15887 25245 15896 25279
rect 15844 25236 15896 25245
rect 14556 25168 14608 25220
rect 14648 25168 14700 25220
rect 18144 25236 18196 25288
rect 20076 25236 20128 25288
rect 14464 25143 14516 25152
rect 14464 25109 14473 25143
rect 14473 25109 14507 25143
rect 14507 25109 14516 25143
rect 14464 25100 14516 25109
rect 25044 25236 25096 25288
rect 27160 25304 27212 25356
rect 31484 25304 31536 25356
rect 31760 25304 31812 25356
rect 32772 25372 32824 25424
rect 33784 25372 33836 25424
rect 45192 25372 45244 25424
rect 25596 25236 25648 25288
rect 26424 25279 26476 25288
rect 26424 25245 26433 25279
rect 26433 25245 26467 25279
rect 26467 25245 26476 25279
rect 26424 25236 26476 25245
rect 29368 25236 29420 25288
rect 22652 25168 22704 25220
rect 25780 25168 25832 25220
rect 27436 25168 27488 25220
rect 29920 25279 29972 25288
rect 29920 25245 29929 25279
rect 29929 25245 29963 25279
rect 29963 25245 29972 25279
rect 30104 25279 30156 25288
rect 29920 25236 29972 25245
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 31116 25236 31168 25288
rect 32588 25304 32640 25356
rect 36084 25304 36136 25356
rect 46296 25347 46348 25356
rect 46296 25313 46305 25347
rect 46305 25313 46339 25347
rect 46339 25313 46348 25347
rect 46296 25304 46348 25313
rect 47952 25347 48004 25356
rect 47952 25313 47961 25347
rect 47961 25313 47995 25347
rect 47995 25313 48004 25347
rect 47952 25304 48004 25313
rect 32772 25279 32824 25288
rect 32772 25245 32781 25279
rect 32781 25245 32815 25279
rect 32815 25245 32824 25279
rect 32772 25236 32824 25245
rect 33324 25236 33376 25288
rect 33508 25236 33560 25288
rect 33784 25279 33836 25288
rect 33784 25245 33793 25279
rect 33793 25245 33827 25279
rect 33827 25245 33836 25279
rect 33784 25236 33836 25245
rect 33968 25279 34020 25288
rect 33968 25245 33977 25279
rect 33977 25245 34011 25279
rect 34011 25245 34020 25279
rect 33968 25236 34020 25245
rect 34704 25236 34756 25288
rect 45468 25279 45520 25288
rect 45468 25245 45477 25279
rect 45477 25245 45511 25279
rect 45511 25245 45520 25279
rect 45468 25236 45520 25245
rect 45928 25236 45980 25288
rect 31024 25211 31076 25220
rect 22744 25100 22796 25152
rect 24768 25143 24820 25152
rect 24768 25109 24777 25143
rect 24777 25109 24811 25143
rect 24811 25109 24820 25143
rect 24768 25100 24820 25109
rect 30472 25100 30524 25152
rect 31024 25177 31033 25211
rect 31033 25177 31067 25211
rect 31067 25177 31076 25211
rect 31024 25168 31076 25177
rect 31852 25211 31904 25220
rect 31852 25177 31861 25211
rect 31861 25177 31895 25211
rect 31895 25177 31904 25211
rect 31852 25168 31904 25177
rect 32220 25100 32272 25152
rect 45560 25143 45612 25152
rect 45560 25109 45569 25143
rect 45569 25109 45603 25143
rect 45603 25109 45612 25143
rect 45560 25100 45612 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 28356 24896 28408 24948
rect 11520 24871 11572 24880
rect 11520 24837 11529 24871
rect 11529 24837 11563 24871
rect 11563 24837 11572 24871
rect 11520 24828 11572 24837
rect 11980 24760 12032 24812
rect 12716 24760 12768 24812
rect 14464 24828 14516 24880
rect 15844 24760 15896 24812
rect 18328 24803 18380 24812
rect 8576 24735 8628 24744
rect 8576 24701 8585 24735
rect 8585 24701 8619 24735
rect 8619 24701 8628 24735
rect 8576 24692 8628 24701
rect 8944 24692 8996 24744
rect 3608 24556 3660 24608
rect 11428 24624 11480 24676
rect 14188 24692 14240 24744
rect 14464 24735 14516 24744
rect 14464 24701 14473 24735
rect 14473 24701 14507 24735
rect 14507 24701 14516 24735
rect 14464 24692 14516 24701
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 23480 24828 23532 24880
rect 26424 24828 26476 24880
rect 29920 24896 29972 24948
rect 31024 24896 31076 24948
rect 32220 24896 32272 24948
rect 44088 24896 44140 24948
rect 29368 24871 29420 24880
rect 29368 24837 29377 24871
rect 29377 24837 29411 24871
rect 29411 24837 29420 24871
rect 29368 24828 29420 24837
rect 30380 24828 30432 24880
rect 34796 24828 34848 24880
rect 19340 24760 19392 24812
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 22100 24803 22152 24812
rect 22100 24769 22109 24803
rect 22109 24769 22143 24803
rect 22143 24769 22152 24803
rect 22100 24760 22152 24769
rect 25136 24803 25188 24812
rect 18512 24692 18564 24744
rect 19984 24692 20036 24744
rect 22744 24735 22796 24744
rect 22744 24701 22753 24735
rect 22753 24701 22787 24735
rect 22787 24701 22796 24735
rect 22744 24692 22796 24701
rect 24768 24692 24820 24744
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25136 24760 25188 24769
rect 25228 24803 25280 24812
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 28540 24760 28592 24812
rect 30472 24803 30524 24812
rect 30472 24769 30481 24803
rect 30481 24769 30515 24803
rect 30515 24769 30524 24803
rect 30472 24760 30524 24769
rect 31484 24803 31536 24812
rect 31484 24769 31493 24803
rect 31493 24769 31527 24803
rect 31527 24769 31536 24803
rect 33876 24803 33928 24812
rect 31484 24760 31536 24769
rect 33876 24769 33885 24803
rect 33885 24769 33919 24803
rect 33919 24769 33928 24803
rect 33876 24760 33928 24769
rect 40040 24760 40092 24812
rect 44272 24760 44324 24812
rect 45100 24803 45152 24812
rect 45100 24769 45109 24803
rect 45109 24769 45143 24803
rect 45143 24769 45152 24803
rect 45100 24760 45152 24769
rect 45652 24760 45704 24812
rect 46388 24760 46440 24812
rect 47492 24760 47544 24812
rect 28080 24692 28132 24744
rect 28632 24735 28684 24744
rect 28632 24701 28641 24735
rect 28641 24701 28675 24735
rect 28675 24701 28684 24735
rect 28632 24692 28684 24701
rect 30656 24692 30708 24744
rect 31760 24692 31812 24744
rect 34152 24735 34204 24744
rect 34152 24701 34161 24735
rect 34161 24701 34195 24735
rect 34195 24701 34204 24735
rect 34152 24692 34204 24701
rect 13912 24624 13964 24676
rect 16120 24624 16172 24676
rect 11704 24599 11756 24608
rect 11704 24565 11713 24599
rect 11713 24565 11747 24599
rect 11747 24565 11756 24599
rect 11704 24556 11756 24565
rect 12072 24556 12124 24608
rect 17776 24556 17828 24608
rect 22652 24624 22704 24676
rect 24860 24624 24912 24676
rect 25044 24624 25096 24676
rect 27712 24624 27764 24676
rect 25504 24556 25556 24608
rect 27988 24556 28040 24608
rect 29644 24556 29696 24608
rect 31116 24556 31168 24608
rect 46204 24692 46256 24744
rect 47400 24692 47452 24744
rect 47676 24803 47728 24812
rect 47676 24769 47685 24803
rect 47685 24769 47719 24803
rect 47719 24769 47728 24803
rect 47676 24760 47728 24769
rect 45652 24624 45704 24676
rect 35624 24599 35676 24608
rect 35624 24565 35633 24599
rect 35633 24565 35667 24599
rect 35667 24565 35676 24599
rect 35624 24556 35676 24565
rect 40408 24599 40460 24608
rect 40408 24565 40417 24599
rect 40417 24565 40451 24599
rect 40451 24565 40460 24599
rect 40408 24556 40460 24565
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 10140 24352 10192 24404
rect 11980 24352 12032 24404
rect 14188 24395 14240 24404
rect 14188 24361 14197 24395
rect 14197 24361 14231 24395
rect 14231 24361 14240 24395
rect 14188 24352 14240 24361
rect 23480 24352 23532 24404
rect 26608 24352 26660 24404
rect 28632 24352 28684 24404
rect 31484 24352 31536 24404
rect 34796 24395 34848 24404
rect 34796 24361 34805 24395
rect 34805 24361 34839 24395
rect 34839 24361 34848 24395
rect 34796 24352 34848 24361
rect 8576 24284 8628 24336
rect 11520 24284 11572 24336
rect 15844 24284 15896 24336
rect 15660 24216 15712 24268
rect 17592 24216 17644 24268
rect 11428 24148 11480 24200
rect 11520 24148 11572 24200
rect 11704 24148 11756 24200
rect 12072 24191 12124 24200
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 13820 24148 13872 24200
rect 13176 24080 13228 24132
rect 13912 24080 13964 24132
rect 16672 24148 16724 24200
rect 16948 24191 17000 24200
rect 16948 24157 16957 24191
rect 16957 24157 16991 24191
rect 16991 24157 17000 24191
rect 16948 24148 17000 24157
rect 18696 24216 18748 24268
rect 27988 24216 28040 24268
rect 28356 24259 28408 24268
rect 28356 24225 28365 24259
rect 28365 24225 28399 24259
rect 28399 24225 28408 24259
rect 28356 24216 28408 24225
rect 16856 24080 16908 24132
rect 17224 24123 17276 24132
rect 17224 24089 17233 24123
rect 17233 24089 17267 24123
rect 17267 24089 17276 24123
rect 17224 24080 17276 24089
rect 20628 24080 20680 24132
rect 22100 24080 22152 24132
rect 25136 24080 25188 24132
rect 26424 24148 26476 24200
rect 26608 24191 26660 24200
rect 26608 24157 26617 24191
rect 26617 24157 26651 24191
rect 26651 24157 26660 24191
rect 26608 24148 26660 24157
rect 27620 24148 27672 24200
rect 28080 24148 28132 24200
rect 28540 24191 28592 24200
rect 28540 24157 28542 24191
rect 28542 24157 28576 24191
rect 28576 24157 28592 24191
rect 33232 24284 33284 24336
rect 34060 24284 34112 24336
rect 31024 24216 31076 24268
rect 35624 24216 35676 24268
rect 40408 24259 40460 24268
rect 40408 24225 40417 24259
rect 40417 24225 40451 24259
rect 40451 24225 40460 24259
rect 40408 24216 40460 24225
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48228 24216 48280 24268
rect 28540 24148 28592 24157
rect 34704 24191 34756 24200
rect 11152 24012 11204 24064
rect 11796 24012 11848 24064
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 12716 24055 12768 24064
rect 12716 24021 12741 24055
rect 12741 24021 12768 24055
rect 12716 24012 12768 24021
rect 14096 24012 14148 24064
rect 15384 24012 15436 24064
rect 18512 24012 18564 24064
rect 25780 24012 25832 24064
rect 26148 24012 26200 24064
rect 26424 24012 26476 24064
rect 28448 24012 28500 24064
rect 28724 24055 28776 24064
rect 28724 24021 28733 24055
rect 28733 24021 28767 24055
rect 28767 24021 28776 24055
rect 28724 24012 28776 24021
rect 30564 24080 30616 24132
rect 34704 24157 34713 24191
rect 34713 24157 34747 24191
rect 34747 24157 34756 24191
rect 34704 24148 34756 24157
rect 40224 24191 40276 24200
rect 40224 24157 40233 24191
rect 40233 24157 40267 24191
rect 40267 24157 40276 24191
rect 40224 24148 40276 24157
rect 43352 24191 43404 24200
rect 43352 24157 43361 24191
rect 43361 24157 43395 24191
rect 43395 24157 43404 24191
rect 43352 24148 43404 24157
rect 43536 24191 43588 24200
rect 43536 24157 43545 24191
rect 43545 24157 43579 24191
rect 43579 24157 43588 24191
rect 43536 24148 43588 24157
rect 45468 24148 45520 24200
rect 45560 24148 45612 24200
rect 31760 24080 31812 24132
rect 32956 24080 33008 24132
rect 44272 24123 44324 24132
rect 44272 24089 44281 24123
rect 44281 24089 44315 24123
rect 44315 24089 44324 24123
rect 44272 24080 44324 24089
rect 45100 24080 45152 24132
rect 46020 24080 46072 24132
rect 46480 24080 46532 24132
rect 37280 24012 37332 24064
rect 43812 24012 43864 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 8944 23851 8996 23860
rect 8944 23817 8953 23851
rect 8953 23817 8987 23851
rect 8987 23817 8996 23851
rect 8944 23808 8996 23817
rect 11152 23808 11204 23860
rect 12072 23808 12124 23860
rect 17224 23808 17276 23860
rect 19340 23808 19392 23860
rect 19984 23851 20036 23860
rect 19984 23817 19993 23851
rect 19993 23817 20027 23851
rect 20027 23817 20036 23851
rect 19984 23808 20036 23817
rect 20628 23851 20680 23860
rect 20628 23817 20637 23851
rect 20637 23817 20671 23851
rect 20671 23817 20680 23851
rect 20628 23808 20680 23817
rect 27804 23808 27856 23860
rect 27988 23808 28040 23860
rect 28448 23851 28500 23860
rect 28448 23817 28457 23851
rect 28457 23817 28491 23851
rect 28491 23817 28500 23851
rect 28448 23808 28500 23817
rect 11520 23783 11572 23792
rect 11520 23749 11529 23783
rect 11529 23749 11563 23783
rect 11563 23749 11572 23783
rect 11520 23740 11572 23749
rect 14096 23783 14148 23792
rect 14096 23749 14105 23783
rect 14105 23749 14139 23783
rect 14139 23749 14148 23783
rect 14096 23740 14148 23749
rect 18420 23783 18472 23792
rect 18420 23749 18429 23783
rect 18429 23749 18463 23783
rect 18463 23749 18472 23783
rect 18420 23740 18472 23749
rect 28080 23783 28132 23792
rect 28080 23749 28089 23783
rect 28089 23749 28123 23783
rect 28123 23749 28132 23783
rect 28080 23740 28132 23749
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 8944 23672 8996 23724
rect 13912 23715 13964 23724
rect 13912 23681 13921 23715
rect 13921 23681 13955 23715
rect 13955 23681 13964 23715
rect 13912 23672 13964 23681
rect 17408 23672 17460 23724
rect 17776 23715 17828 23724
rect 17776 23681 17785 23715
rect 17785 23681 17819 23715
rect 17819 23681 17828 23715
rect 17776 23672 17828 23681
rect 18788 23672 18840 23724
rect 20720 23672 20772 23724
rect 22100 23672 22152 23724
rect 26148 23715 26200 23724
rect 26148 23681 26157 23715
rect 26157 23681 26191 23715
rect 26191 23681 26200 23715
rect 26148 23672 26200 23681
rect 26424 23715 26476 23724
rect 26424 23681 26433 23715
rect 26433 23681 26467 23715
rect 26467 23681 26476 23715
rect 26424 23672 26476 23681
rect 28356 23672 28408 23724
rect 28724 23672 28776 23724
rect 30196 23808 30248 23860
rect 30564 23851 30616 23860
rect 30564 23817 30573 23851
rect 30573 23817 30607 23851
rect 30607 23817 30616 23851
rect 30564 23808 30616 23817
rect 29736 23715 29788 23724
rect 29736 23681 29745 23715
rect 29745 23681 29779 23715
rect 29779 23681 29788 23715
rect 29736 23672 29788 23681
rect 11796 23579 11848 23588
rect 11796 23545 11805 23579
rect 11805 23545 11839 23579
rect 11839 23545 11848 23579
rect 11796 23536 11848 23545
rect 14188 23604 14240 23656
rect 30472 23740 30524 23792
rect 30196 23715 30248 23724
rect 30196 23681 30205 23715
rect 30205 23681 30239 23715
rect 30239 23681 30248 23715
rect 30196 23672 30248 23681
rect 30932 23672 30984 23724
rect 32772 23740 32824 23792
rect 33416 23740 33468 23792
rect 34704 23808 34756 23860
rect 40224 23808 40276 23860
rect 43352 23808 43404 23860
rect 45560 23808 45612 23860
rect 42800 23783 42852 23792
rect 42800 23749 42809 23783
rect 42809 23749 42843 23783
rect 42843 23749 42852 23783
rect 42800 23740 42852 23749
rect 44364 23740 44416 23792
rect 45008 23740 45060 23792
rect 45376 23740 45428 23792
rect 34428 23672 34480 23724
rect 38384 23672 38436 23724
rect 42616 23672 42668 23724
rect 43812 23715 43864 23724
rect 43812 23681 43821 23715
rect 43821 23681 43855 23715
rect 43855 23681 43864 23715
rect 43812 23672 43864 23681
rect 45468 23672 45520 23724
rect 33600 23536 33652 23588
rect 11704 23468 11756 23520
rect 16764 23511 16816 23520
rect 16764 23477 16773 23511
rect 16773 23477 16807 23511
rect 16807 23477 16816 23511
rect 16764 23468 16816 23477
rect 16856 23468 16908 23520
rect 18328 23468 18380 23520
rect 18788 23511 18840 23520
rect 18788 23477 18797 23511
rect 18797 23477 18831 23511
rect 18831 23477 18840 23511
rect 18788 23468 18840 23477
rect 21916 23511 21968 23520
rect 21916 23477 21925 23511
rect 21925 23477 21959 23511
rect 21959 23477 21968 23511
rect 21916 23468 21968 23477
rect 25320 23468 25372 23520
rect 26976 23468 27028 23520
rect 28080 23468 28132 23520
rect 30932 23468 30984 23520
rect 31208 23468 31260 23520
rect 32772 23511 32824 23520
rect 32772 23477 32781 23511
rect 32781 23477 32815 23511
rect 32815 23477 32824 23511
rect 32772 23468 32824 23477
rect 43720 23647 43772 23656
rect 43720 23613 43729 23647
rect 43729 23613 43763 23647
rect 43763 23613 43772 23647
rect 43720 23604 43772 23613
rect 46296 23647 46348 23656
rect 46296 23613 46305 23647
rect 46305 23613 46339 23647
rect 46339 23613 46348 23647
rect 46296 23604 46348 23613
rect 48044 23536 48096 23588
rect 47676 23511 47728 23520
rect 47676 23477 47685 23511
rect 47685 23477 47719 23511
rect 47719 23477 47728 23511
rect 47676 23468 47728 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 16948 23264 17000 23316
rect 26608 23264 26660 23316
rect 32956 23307 33008 23316
rect 32956 23273 32965 23307
rect 32965 23273 32999 23307
rect 32999 23273 33008 23307
rect 32956 23264 33008 23273
rect 42616 23264 42668 23316
rect 16856 23196 16908 23248
rect 28816 23196 28868 23248
rect 42800 23196 42852 23248
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 15384 23171 15436 23180
rect 15384 23137 15393 23171
rect 15393 23137 15427 23171
rect 15427 23137 15436 23171
rect 15384 23128 15436 23137
rect 15660 23171 15712 23180
rect 15660 23137 15669 23171
rect 15669 23137 15703 23171
rect 15703 23137 15712 23171
rect 15660 23128 15712 23137
rect 16672 23128 16724 23180
rect 11428 23103 11480 23112
rect 11428 23069 11437 23103
rect 11437 23069 11471 23103
rect 11471 23069 11480 23103
rect 11428 23060 11480 23069
rect 14648 23060 14700 23112
rect 15016 23060 15068 23112
rect 16764 23060 16816 23112
rect 20904 23128 20956 23180
rect 22744 23128 22796 23180
rect 24952 23128 25004 23180
rect 25412 23128 25464 23180
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 19340 23060 19392 23112
rect 11336 22992 11388 23044
rect 12440 22992 12492 23044
rect 23204 23060 23256 23112
rect 27620 23103 27672 23112
rect 27620 23069 27629 23103
rect 27629 23069 27663 23103
rect 27663 23069 27672 23103
rect 27620 23060 27672 23069
rect 28356 23060 28408 23112
rect 30380 23128 30432 23180
rect 32036 23128 32088 23180
rect 40224 23128 40276 23180
rect 41420 23171 41472 23180
rect 41420 23137 41429 23171
rect 41429 23137 41463 23171
rect 41463 23137 41472 23171
rect 41420 23128 41472 23137
rect 43352 23128 43404 23180
rect 29736 23060 29788 23112
rect 30196 23103 30248 23112
rect 30196 23069 30205 23103
rect 30205 23069 30239 23103
rect 30239 23069 30248 23103
rect 30196 23060 30248 23069
rect 30748 23060 30800 23112
rect 33416 23103 33468 23112
rect 33416 23069 33425 23103
rect 33425 23069 33459 23103
rect 33459 23069 33468 23103
rect 33416 23060 33468 23069
rect 40684 23060 40736 23112
rect 43076 23060 43128 23112
rect 43720 23060 43772 23112
rect 46664 23196 46716 23248
rect 47676 23128 47728 23180
rect 48136 23171 48188 23180
rect 48136 23137 48145 23171
rect 48145 23137 48179 23171
rect 48179 23137 48188 23171
rect 48136 23128 48188 23137
rect 44364 23103 44416 23112
rect 44364 23069 44373 23103
rect 44373 23069 44407 23103
rect 44407 23069 44416 23103
rect 44364 23060 44416 23069
rect 45468 23060 45520 23112
rect 10232 22924 10284 22976
rect 13176 22967 13228 22976
rect 13176 22933 13185 22967
rect 13185 22933 13219 22967
rect 13219 22933 13228 22967
rect 13176 22924 13228 22933
rect 13912 22924 13964 22976
rect 20168 22924 20220 22976
rect 21916 22992 21968 23044
rect 25320 23035 25372 23044
rect 25320 23001 25329 23035
rect 25329 23001 25363 23035
rect 25363 23001 25372 23035
rect 25320 22992 25372 23001
rect 27712 22992 27764 23044
rect 28080 22992 28132 23044
rect 28724 22992 28776 23044
rect 30288 22992 30340 23044
rect 30656 22992 30708 23044
rect 32772 22992 32824 23044
rect 20628 22924 20680 22976
rect 21824 22967 21876 22976
rect 21824 22933 21833 22967
rect 21833 22933 21867 22967
rect 21867 22933 21876 22967
rect 21824 22924 21876 22933
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 28448 22967 28500 22976
rect 28448 22933 28457 22967
rect 28457 22933 28491 22967
rect 28491 22933 28500 22967
rect 28448 22924 28500 22933
rect 31024 22924 31076 22976
rect 33508 22967 33560 22976
rect 33508 22933 33517 22967
rect 33517 22933 33551 22967
rect 33551 22933 33560 22967
rect 33508 22924 33560 22933
rect 45836 22992 45888 23044
rect 43536 22924 43588 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 11428 22720 11480 22772
rect 12440 22720 12492 22772
rect 18420 22720 18472 22772
rect 19248 22763 19300 22772
rect 19248 22729 19257 22763
rect 19257 22729 19291 22763
rect 19291 22729 19300 22763
rect 19248 22720 19300 22729
rect 27712 22763 27764 22772
rect 27712 22729 27721 22763
rect 27721 22729 27755 22763
rect 27755 22729 27764 22763
rect 27712 22720 27764 22729
rect 30196 22720 30248 22772
rect 30472 22720 30524 22772
rect 31852 22720 31904 22772
rect 39764 22720 39816 22772
rect 40684 22763 40736 22772
rect 40684 22729 40693 22763
rect 40693 22729 40727 22763
rect 40727 22729 40736 22763
rect 40684 22720 40736 22729
rect 45652 22720 45704 22772
rect 47584 22720 47636 22772
rect 3516 22652 3568 22704
rect 9956 22627 10008 22636
rect 9956 22593 9965 22627
rect 9965 22593 9999 22627
rect 9999 22593 10008 22627
rect 9956 22584 10008 22593
rect 11152 22516 11204 22568
rect 11336 22584 11388 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 13176 22584 13228 22636
rect 17408 22627 17460 22636
rect 17408 22593 17417 22627
rect 17417 22593 17451 22627
rect 17451 22593 17460 22627
rect 17408 22584 17460 22593
rect 18420 22584 18472 22636
rect 12808 22516 12860 22568
rect 13820 22559 13872 22568
rect 13820 22525 13829 22559
rect 13829 22525 13863 22559
rect 13863 22525 13872 22559
rect 13820 22516 13872 22525
rect 15568 22516 15620 22568
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 12440 22448 12492 22500
rect 18328 22448 18380 22500
rect 27896 22652 27948 22704
rect 29552 22652 29604 22704
rect 30288 22652 30340 22704
rect 31024 22695 31076 22704
rect 31024 22661 31033 22695
rect 31033 22661 31067 22695
rect 31067 22661 31076 22695
rect 31024 22652 31076 22661
rect 31208 22695 31260 22704
rect 31208 22661 31217 22695
rect 31217 22661 31251 22695
rect 31251 22661 31260 22695
rect 31208 22652 31260 22661
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 27436 22584 27488 22636
rect 28724 22627 28776 22636
rect 28724 22593 28733 22627
rect 28733 22593 28767 22627
rect 28767 22593 28776 22627
rect 28724 22584 28776 22593
rect 22008 22516 22060 22568
rect 24124 22559 24176 22568
rect 24124 22525 24133 22559
rect 24133 22525 24167 22559
rect 24167 22525 24176 22559
rect 24124 22516 24176 22525
rect 24308 22559 24360 22568
rect 24308 22525 24317 22559
rect 24317 22525 24351 22559
rect 24351 22525 24360 22559
rect 24308 22516 24360 22525
rect 29092 22627 29144 22636
rect 29092 22593 29101 22627
rect 29101 22593 29135 22627
rect 29135 22593 29144 22627
rect 29092 22584 29144 22593
rect 30380 22584 30432 22636
rect 32036 22584 32088 22636
rect 33508 22584 33560 22636
rect 40132 22584 40184 22636
rect 29736 22559 29788 22568
rect 29736 22525 29745 22559
rect 29745 22525 29779 22559
rect 29779 22525 29788 22559
rect 29736 22516 29788 22525
rect 31760 22516 31812 22568
rect 45284 22584 45336 22636
rect 45652 22584 45704 22636
rect 47860 22627 47912 22636
rect 47860 22593 47869 22627
rect 47869 22593 47903 22627
rect 47903 22593 47912 22627
rect 47860 22584 47912 22593
rect 48044 22584 48096 22636
rect 46020 22516 46072 22568
rect 46204 22559 46256 22568
rect 46204 22525 46213 22559
rect 46213 22525 46247 22559
rect 46247 22525 46256 22559
rect 46204 22516 46256 22525
rect 44272 22448 44324 22500
rect 47768 22516 47820 22568
rect 10324 22423 10376 22432
rect 10324 22389 10333 22423
rect 10333 22389 10367 22423
rect 10367 22389 10376 22423
rect 10324 22380 10376 22389
rect 11060 22380 11112 22432
rect 17960 22380 18012 22432
rect 27068 22423 27120 22432
rect 27068 22389 27077 22423
rect 27077 22389 27111 22423
rect 27111 22389 27120 22423
rect 27068 22380 27120 22389
rect 29276 22423 29328 22432
rect 29276 22389 29285 22423
rect 29285 22389 29319 22423
rect 29319 22389 29328 22423
rect 29276 22380 29328 22389
rect 31944 22380 31996 22432
rect 39764 22380 39816 22432
rect 40316 22423 40368 22432
rect 40316 22389 40325 22423
rect 40325 22389 40359 22423
rect 40359 22389 40368 22423
rect 40316 22380 40368 22389
rect 45652 22380 45704 22432
rect 45744 22423 45796 22432
rect 45744 22389 45753 22423
rect 45753 22389 45787 22423
rect 45787 22389 45796 22423
rect 45744 22380 45796 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 10324 22176 10376 22228
rect 18052 22176 18104 22228
rect 25872 22176 25924 22228
rect 43076 22219 43128 22228
rect 9956 22108 10008 22160
rect 10232 22083 10284 22092
rect 10232 22049 10241 22083
rect 10241 22049 10275 22083
rect 10275 22049 10284 22083
rect 10232 22040 10284 22049
rect 12808 22108 12860 22160
rect 29092 22108 29144 22160
rect 43076 22185 43085 22219
rect 43085 22185 43119 22219
rect 43119 22185 43128 22219
rect 43076 22176 43128 22185
rect 42892 22108 42944 22160
rect 11980 22083 12032 22092
rect 11980 22049 11989 22083
rect 11989 22049 12023 22083
rect 12023 22049 12032 22083
rect 11980 22040 12032 22049
rect 13820 22040 13872 22092
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 18420 22040 18472 22092
rect 20904 22083 20956 22092
rect 8944 22015 8996 22024
rect 8944 21981 8953 22015
rect 8953 21981 8987 22015
rect 8987 21981 8996 22015
rect 8944 21972 8996 21981
rect 12532 22015 12584 22024
rect 8852 21836 8904 21888
rect 9128 21836 9180 21888
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 11060 21904 11112 21956
rect 13912 21972 13964 22024
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 16580 22015 16632 22024
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 17960 21972 18012 22024
rect 18328 21972 18380 22024
rect 18788 21972 18840 22024
rect 14648 21904 14700 21956
rect 18696 21904 18748 21956
rect 19248 21947 19300 21956
rect 19248 21913 19257 21947
rect 19257 21913 19291 21947
rect 19291 21913 19300 21947
rect 19248 21904 19300 21913
rect 20904 22049 20913 22083
rect 20913 22049 20947 22083
rect 20947 22049 20956 22083
rect 20904 22040 20956 22049
rect 24308 22040 24360 22092
rect 27620 22040 27672 22092
rect 21456 21972 21508 22024
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23204 21972 23256 21981
rect 25504 22015 25556 22024
rect 25504 21981 25513 22015
rect 25513 21981 25547 22015
rect 25547 21981 25556 22015
rect 25504 21972 25556 21981
rect 45560 22040 45612 22092
rect 46940 22083 46992 22092
rect 46940 22049 46949 22083
rect 46949 22049 46983 22083
rect 46983 22049 46992 22083
rect 46940 22040 46992 22049
rect 29276 21972 29328 22024
rect 31944 22015 31996 22024
rect 31944 21981 31953 22015
rect 31953 21981 31987 22015
rect 31987 21981 31996 22015
rect 31944 21972 31996 21981
rect 33876 21972 33928 22024
rect 40132 22015 40184 22024
rect 40132 21981 40141 22015
rect 40141 21981 40175 22015
rect 40175 21981 40184 22015
rect 40132 21972 40184 21981
rect 40316 22015 40368 22024
rect 40316 21981 40325 22015
rect 40325 21981 40359 22015
rect 40359 21981 40368 22015
rect 40316 21972 40368 21981
rect 43444 21972 43496 22024
rect 45192 21972 45244 22024
rect 27068 21904 27120 21956
rect 28816 21947 28868 21956
rect 28816 21913 28825 21947
rect 28825 21913 28859 21947
rect 28859 21913 28868 21947
rect 28816 21904 28868 21913
rect 40592 21904 40644 21956
rect 43076 21947 43128 21956
rect 43076 21913 43085 21947
rect 43085 21913 43119 21947
rect 43119 21913 43128 21947
rect 43076 21904 43128 21913
rect 18420 21836 18472 21888
rect 18512 21836 18564 21888
rect 27712 21836 27764 21888
rect 31760 21879 31812 21888
rect 31760 21845 31769 21879
rect 31769 21845 31803 21879
rect 31803 21845 31812 21879
rect 31760 21836 31812 21845
rect 34520 21836 34572 21888
rect 43352 21836 43404 21888
rect 45284 21879 45336 21888
rect 45284 21845 45293 21879
rect 45293 21845 45327 21879
rect 45327 21845 45336 21879
rect 45284 21836 45336 21845
rect 45468 21836 45520 21888
rect 45652 21904 45704 21956
rect 47768 21836 47820 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 20 21564 72 21616
rect 10968 21632 11020 21684
rect 14648 21675 14700 21684
rect 14648 21641 14657 21675
rect 14657 21641 14691 21675
rect 14691 21641 14700 21675
rect 14648 21632 14700 21641
rect 16672 21632 16724 21684
rect 8852 21607 8904 21616
rect 8852 21573 8861 21607
rect 8861 21573 8895 21607
rect 8895 21573 8904 21607
rect 8852 21564 8904 21573
rect 12532 21564 12584 21616
rect 13728 21564 13780 21616
rect 13912 21496 13964 21548
rect 18420 21564 18472 21616
rect 28724 21632 28776 21684
rect 33876 21675 33928 21684
rect 33876 21641 33885 21675
rect 33885 21641 33919 21675
rect 33919 21641 33928 21675
rect 33876 21632 33928 21641
rect 42892 21632 42944 21684
rect 21824 21564 21876 21616
rect 23480 21564 23532 21616
rect 27712 21607 27764 21616
rect 27712 21573 27721 21607
rect 27721 21573 27755 21607
rect 27755 21573 27764 21607
rect 27712 21564 27764 21573
rect 28172 21564 28224 21616
rect 34428 21607 34480 21616
rect 34428 21573 34437 21607
rect 34437 21573 34471 21607
rect 34471 21573 34480 21607
rect 34428 21564 34480 21573
rect 34520 21607 34572 21616
rect 34520 21573 34529 21607
rect 34529 21573 34563 21607
rect 34563 21573 34572 21607
rect 34520 21564 34572 21573
rect 43076 21607 43128 21616
rect 43076 21573 43085 21607
rect 43085 21573 43119 21607
rect 43119 21573 43128 21607
rect 43076 21564 43128 21573
rect 18328 21496 18380 21548
rect 18512 21539 18564 21548
rect 18512 21505 18521 21539
rect 18521 21505 18555 21539
rect 18555 21505 18564 21539
rect 18512 21496 18564 21505
rect 20168 21496 20220 21548
rect 25504 21496 25556 21548
rect 18052 21428 18104 21480
rect 22284 21471 22336 21480
rect 22284 21437 22293 21471
rect 22293 21437 22327 21471
rect 22327 21437 22336 21471
rect 22284 21428 22336 21437
rect 23020 21471 23072 21480
rect 23020 21437 23029 21471
rect 23029 21437 23063 21471
rect 23063 21437 23072 21471
rect 23020 21428 23072 21437
rect 42340 21496 42392 21548
rect 42708 21496 42760 21548
rect 44180 21539 44232 21548
rect 44180 21505 44189 21539
rect 44189 21505 44223 21539
rect 44223 21505 44232 21539
rect 45560 21564 45612 21616
rect 46020 21632 46072 21684
rect 44180 21496 44232 21505
rect 45192 21496 45244 21548
rect 46204 21539 46256 21548
rect 46204 21505 46213 21539
rect 46213 21505 46247 21539
rect 46247 21505 46256 21539
rect 46204 21496 46256 21505
rect 47584 21539 47636 21548
rect 47584 21505 47593 21539
rect 47593 21505 47627 21539
rect 47627 21505 47636 21539
rect 47584 21496 47636 21505
rect 48044 21496 48096 21548
rect 47860 21471 47912 21480
rect 47860 21437 47869 21471
rect 47869 21437 47903 21471
rect 47903 21437 47912 21471
rect 47860 21428 47912 21437
rect 3792 21292 3844 21344
rect 18512 21335 18564 21344
rect 18512 21301 18521 21335
rect 18521 21301 18555 21335
rect 18555 21301 18564 21335
rect 18512 21292 18564 21301
rect 20996 21335 21048 21344
rect 20996 21301 21005 21335
rect 21005 21301 21039 21335
rect 21039 21301 21048 21335
rect 20996 21292 21048 21301
rect 22376 21292 22428 21344
rect 34244 21292 34296 21344
rect 35808 21360 35860 21412
rect 42800 21360 42852 21412
rect 43352 21403 43404 21412
rect 43352 21369 43361 21403
rect 43361 21369 43395 21403
rect 43395 21369 43404 21403
rect 43352 21360 43404 21369
rect 45284 21360 45336 21412
rect 35900 21292 35952 21344
rect 43536 21335 43588 21344
rect 43536 21301 43545 21335
rect 43545 21301 43579 21335
rect 43579 21301 43588 21335
rect 43536 21292 43588 21301
rect 44640 21335 44692 21344
rect 44640 21301 44649 21335
rect 44649 21301 44683 21335
rect 44683 21301 44692 21335
rect 44640 21292 44692 21301
rect 45468 21335 45520 21344
rect 45468 21301 45477 21335
rect 45477 21301 45511 21335
rect 45511 21301 45520 21335
rect 45468 21292 45520 21301
rect 45836 21292 45888 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 16580 21131 16632 21140
rect 16580 21097 16589 21131
rect 16589 21097 16623 21131
rect 16623 21097 16632 21131
rect 16580 21088 16632 21097
rect 23020 21088 23072 21140
rect 27436 21088 27488 21140
rect 28172 21088 28224 21140
rect 9956 21020 10008 21072
rect 35808 21063 35860 21072
rect 9128 20995 9180 21004
rect 9128 20961 9137 20995
rect 9137 20961 9171 20995
rect 9171 20961 9180 20995
rect 9128 20952 9180 20961
rect 35808 21029 35817 21063
rect 35817 21029 35851 21063
rect 35851 21029 35860 21063
rect 35808 21020 35860 21029
rect 22376 20995 22428 21004
rect 22376 20961 22385 20995
rect 22385 20961 22419 20995
rect 22419 20961 22428 20995
rect 22376 20952 22428 20961
rect 26792 20952 26844 21004
rect 44272 21020 44324 21072
rect 43444 20995 43496 21004
rect 43444 20961 43453 20995
rect 43453 20961 43487 20995
rect 43487 20961 43496 20995
rect 43444 20952 43496 20961
rect 44088 20995 44140 21004
rect 44088 20961 44097 20995
rect 44097 20961 44131 20995
rect 44131 20961 44140 20995
rect 44088 20952 44140 20961
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 14832 20927 14884 20936
rect 10784 20859 10836 20868
rect 10784 20825 10793 20859
rect 10793 20825 10827 20859
rect 10827 20825 10836 20859
rect 10784 20816 10836 20825
rect 14832 20893 14841 20927
rect 14841 20893 14875 20927
rect 14875 20893 14884 20927
rect 14832 20884 14884 20893
rect 16672 20884 16724 20936
rect 19156 20884 19208 20936
rect 20996 20884 21048 20936
rect 23480 20884 23532 20936
rect 25964 20884 26016 20936
rect 27436 20884 27488 20936
rect 30564 20927 30616 20936
rect 30564 20893 30573 20927
rect 30573 20893 30607 20927
rect 30607 20893 30616 20927
rect 30564 20884 30616 20893
rect 43536 20927 43588 20936
rect 43536 20893 43545 20927
rect 43545 20893 43579 20927
rect 43579 20893 43588 20927
rect 43536 20884 43588 20893
rect 45836 20927 45888 20936
rect 45836 20893 45845 20927
rect 45845 20893 45879 20927
rect 45879 20893 45888 20927
rect 45836 20884 45888 20893
rect 15108 20816 15160 20868
rect 31760 20859 31812 20868
rect 31760 20825 31769 20859
rect 31769 20825 31803 20859
rect 31803 20825 31812 20859
rect 31760 20816 31812 20825
rect 32588 20816 32640 20868
rect 32864 20816 32916 20868
rect 35900 20816 35952 20868
rect 36360 20816 36412 20868
rect 47676 20816 47728 20868
rect 14096 20748 14148 20800
rect 14556 20748 14608 20800
rect 14924 20791 14976 20800
rect 14924 20757 14933 20791
rect 14933 20757 14967 20791
rect 14967 20757 14976 20791
rect 14924 20748 14976 20757
rect 17960 20748 18012 20800
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 30656 20791 30708 20800
rect 30656 20757 30665 20791
rect 30665 20757 30699 20791
rect 30699 20757 30708 20791
rect 30656 20748 30708 20757
rect 45928 20748 45980 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3976 20544 4028 20596
rect 14188 20544 14240 20596
rect 19248 20544 19300 20596
rect 22008 20544 22060 20596
rect 22284 20544 22336 20596
rect 23480 20544 23532 20596
rect 32864 20544 32916 20596
rect 45744 20544 45796 20596
rect 47676 20587 47728 20596
rect 47676 20553 47685 20587
rect 47685 20553 47719 20587
rect 47719 20553 47728 20587
rect 47676 20544 47728 20553
rect 10968 20476 11020 20528
rect 11152 20408 11204 20460
rect 18512 20476 18564 20528
rect 24124 20476 24176 20528
rect 32220 20519 32272 20528
rect 32220 20485 32229 20519
rect 32229 20485 32263 20519
rect 32263 20485 32272 20519
rect 32220 20476 32272 20485
rect 32312 20519 32364 20528
rect 32312 20485 32321 20519
rect 32321 20485 32355 20519
rect 32355 20485 32364 20519
rect 32312 20476 32364 20485
rect 12716 20408 12768 20460
rect 12808 20451 12860 20460
rect 12808 20417 12817 20451
rect 12817 20417 12851 20451
rect 12851 20417 12860 20451
rect 12808 20408 12860 20417
rect 14924 20408 14976 20460
rect 15108 20408 15160 20460
rect 17960 20451 18012 20460
rect 17960 20417 17969 20451
rect 17969 20417 18003 20451
rect 18003 20417 18012 20451
rect 17960 20408 18012 20417
rect 19340 20408 19392 20460
rect 20996 20451 21048 20460
rect 20996 20417 21005 20451
rect 21005 20417 21039 20451
rect 21039 20417 21048 20451
rect 20996 20408 21048 20417
rect 21916 20408 21968 20460
rect 12992 20340 13044 20392
rect 15660 20340 15712 20392
rect 20168 20340 20220 20392
rect 19248 20272 19300 20324
rect 22192 20272 22244 20324
rect 22744 20272 22796 20324
rect 25412 20408 25464 20460
rect 27436 20408 27488 20460
rect 30012 20408 30064 20460
rect 44088 20476 44140 20528
rect 44640 20476 44692 20528
rect 42800 20451 42852 20460
rect 28540 20383 28592 20392
rect 28540 20349 28549 20383
rect 28549 20349 28583 20383
rect 28583 20349 28592 20383
rect 28540 20340 28592 20349
rect 28816 20383 28868 20392
rect 28816 20349 28825 20383
rect 28825 20349 28859 20383
rect 28859 20349 28868 20383
rect 28816 20340 28868 20349
rect 32312 20340 32364 20392
rect 32588 20383 32640 20392
rect 32588 20349 32597 20383
rect 32597 20349 32631 20383
rect 32631 20349 32640 20383
rect 32588 20340 32640 20349
rect 40408 20340 40460 20392
rect 41880 20383 41932 20392
rect 41880 20349 41889 20383
rect 41889 20349 41923 20383
rect 41923 20349 41932 20383
rect 41880 20340 41932 20349
rect 42800 20417 42809 20451
rect 42809 20417 42843 20451
rect 42843 20417 42852 20451
rect 42800 20408 42852 20417
rect 43720 20451 43772 20460
rect 43720 20417 43729 20451
rect 43729 20417 43763 20451
rect 43763 20417 43772 20451
rect 43720 20408 43772 20417
rect 46756 20408 46808 20460
rect 43076 20340 43128 20392
rect 43812 20383 43864 20392
rect 43812 20349 43821 20383
rect 43821 20349 43855 20383
rect 43855 20349 43864 20383
rect 43812 20340 43864 20349
rect 45836 20383 45888 20392
rect 45836 20349 45845 20383
rect 45845 20349 45879 20383
rect 45879 20349 45888 20383
rect 45836 20340 45888 20349
rect 46940 20340 46992 20392
rect 28724 20272 28776 20324
rect 11428 20204 11480 20256
rect 15108 20204 15160 20256
rect 18236 20204 18288 20256
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 21916 20204 21968 20256
rect 23020 20204 23072 20256
rect 25044 20204 25096 20256
rect 26332 20247 26384 20256
rect 26332 20213 26341 20247
rect 26341 20213 26375 20247
rect 26375 20213 26384 20247
rect 26332 20204 26384 20213
rect 27068 20247 27120 20256
rect 27068 20213 27077 20247
rect 27077 20213 27111 20247
rect 27111 20213 27120 20247
rect 27068 20204 27120 20213
rect 28172 20204 28224 20256
rect 40684 20272 40736 20324
rect 46296 20272 46348 20324
rect 31300 20247 31352 20256
rect 31300 20213 31309 20247
rect 31309 20213 31343 20247
rect 31343 20213 31352 20247
rect 31300 20204 31352 20213
rect 32312 20204 32364 20256
rect 42616 20247 42668 20256
rect 42616 20213 42625 20247
rect 42625 20213 42659 20247
rect 42659 20213 42668 20247
rect 42616 20204 42668 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3424 20000 3476 20052
rect 28816 20000 28868 20052
rect 40408 20043 40460 20052
rect 40408 20009 40417 20043
rect 40417 20009 40451 20043
rect 40451 20009 40460 20043
rect 40408 20000 40460 20009
rect 42156 20000 42208 20052
rect 12716 19932 12768 19984
rect 14372 19932 14424 19984
rect 15660 19975 15712 19984
rect 15660 19941 15669 19975
rect 15669 19941 15703 19975
rect 15703 19941 15712 19975
rect 15660 19932 15712 19941
rect 11428 19907 11480 19916
rect 11428 19873 11437 19907
rect 11437 19873 11471 19907
rect 11471 19873 11480 19907
rect 11428 19864 11480 19873
rect 1768 19796 1820 19848
rect 14832 19864 14884 19916
rect 15016 19864 15068 19916
rect 21088 19907 21140 19916
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 15108 19796 15160 19848
rect 16672 19796 16724 19848
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 19156 19796 19208 19848
rect 14188 19728 14240 19780
rect 12808 19660 12860 19712
rect 14372 19703 14424 19712
rect 14372 19669 14381 19703
rect 14381 19669 14415 19703
rect 14415 19669 14424 19703
rect 14372 19660 14424 19669
rect 14648 19660 14700 19712
rect 17224 19660 17276 19712
rect 18236 19660 18288 19712
rect 21088 19873 21097 19907
rect 21097 19873 21131 19907
rect 21131 19873 21140 19907
rect 21088 19864 21140 19873
rect 21456 19864 21508 19916
rect 22744 19864 22796 19916
rect 21088 19728 21140 19780
rect 22376 19728 22428 19780
rect 24124 19932 24176 19984
rect 43444 19975 43496 19984
rect 25044 19907 25096 19916
rect 25044 19873 25053 19907
rect 25053 19873 25087 19907
rect 25087 19873 25096 19907
rect 25044 19864 25096 19873
rect 26884 19864 26936 19916
rect 27160 19864 27212 19916
rect 28264 19864 28316 19916
rect 28816 19864 28868 19916
rect 30656 19907 30708 19916
rect 30656 19873 30665 19907
rect 30665 19873 30699 19907
rect 30699 19873 30708 19907
rect 30656 19864 30708 19873
rect 33048 19864 33100 19916
rect 43444 19941 43453 19975
rect 43453 19941 43487 19975
rect 43487 19941 43496 19975
rect 43444 19932 43496 19941
rect 43720 20000 43772 20052
rect 45836 19932 45888 19984
rect 40684 19864 40736 19916
rect 42616 19864 42668 19916
rect 45744 19907 45796 19916
rect 24860 19796 24912 19848
rect 28356 19839 28408 19848
rect 28356 19805 28365 19839
rect 28365 19805 28399 19839
rect 28399 19805 28408 19839
rect 28356 19796 28408 19805
rect 26332 19728 26384 19780
rect 27160 19728 27212 19780
rect 28908 19660 28960 19712
rect 42248 19796 42300 19848
rect 43260 19839 43312 19848
rect 43260 19805 43269 19839
rect 43269 19805 43303 19839
rect 43303 19805 43312 19839
rect 43260 19796 43312 19805
rect 43444 19839 43496 19848
rect 43444 19805 43453 19839
rect 43453 19805 43487 19839
rect 43487 19805 43496 19839
rect 45744 19873 45753 19907
rect 45753 19873 45787 19907
rect 45787 19873 45796 19907
rect 45744 19864 45796 19873
rect 45928 19907 45980 19916
rect 45928 19873 45937 19907
rect 45937 19873 45971 19907
rect 45971 19873 45980 19907
rect 45928 19864 45980 19873
rect 43444 19796 43496 19805
rect 45560 19796 45612 19848
rect 43720 19728 43772 19780
rect 41144 19660 41196 19712
rect 46480 19728 46532 19780
rect 45008 19660 45060 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 13912 19456 13964 19508
rect 15016 19456 15068 19508
rect 20168 19456 20220 19508
rect 14372 19388 14424 19440
rect 14740 19388 14792 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 12808 19320 12860 19372
rect 14004 19320 14056 19372
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14556 19320 14608 19372
rect 18236 19388 18288 19440
rect 21088 19456 21140 19508
rect 22376 19456 22428 19508
rect 28356 19499 28408 19508
rect 17224 19363 17276 19372
rect 17224 19329 17233 19363
rect 17233 19329 17267 19363
rect 17267 19329 17276 19363
rect 17224 19320 17276 19329
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 1584 19184 1636 19236
rect 14280 19184 14332 19236
rect 12992 19116 13044 19168
rect 14648 19116 14700 19168
rect 18512 19252 18564 19304
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 23020 19388 23072 19440
rect 22192 19363 22244 19372
rect 20168 19320 20220 19329
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 26240 19388 26292 19440
rect 27160 19388 27212 19440
rect 27988 19431 28040 19440
rect 27988 19397 27997 19431
rect 27997 19397 28031 19431
rect 28031 19397 28040 19431
rect 27988 19388 28040 19397
rect 28356 19465 28365 19499
rect 28365 19465 28399 19499
rect 28399 19465 28408 19499
rect 28356 19456 28408 19465
rect 28540 19456 28592 19508
rect 31760 19456 31812 19508
rect 43444 19456 43496 19508
rect 43812 19499 43864 19508
rect 43812 19465 43821 19499
rect 43821 19465 43855 19499
rect 43855 19465 43864 19499
rect 43812 19456 43864 19465
rect 20812 19252 20864 19304
rect 20904 19252 20956 19304
rect 25412 19363 25464 19372
rect 25412 19329 25421 19363
rect 25421 19329 25455 19363
rect 25455 19329 25464 19363
rect 25412 19320 25464 19329
rect 28172 19363 28224 19372
rect 28172 19329 28181 19363
rect 28181 19329 28215 19363
rect 28215 19329 28224 19363
rect 28172 19320 28224 19329
rect 24676 19295 24728 19304
rect 24676 19261 24685 19295
rect 24685 19261 24719 19295
rect 24719 19261 24728 19295
rect 24676 19252 24728 19261
rect 28724 19388 28776 19440
rect 28816 19363 28868 19372
rect 28816 19329 28825 19363
rect 28825 19329 28859 19363
rect 28859 19329 28868 19363
rect 28816 19320 28868 19329
rect 30380 19388 30432 19440
rect 25504 19184 25556 19236
rect 30472 19252 30524 19304
rect 41420 19388 41472 19440
rect 42156 19388 42208 19440
rect 42248 19388 42300 19440
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 42800 19320 42852 19372
rect 43076 19363 43128 19372
rect 43076 19329 43085 19363
rect 43085 19329 43119 19363
rect 43119 19329 43128 19363
rect 43076 19320 43128 19329
rect 44180 19388 44232 19440
rect 43904 19363 43956 19372
rect 43904 19329 43913 19363
rect 43913 19329 43947 19363
rect 43947 19329 43956 19363
rect 43904 19320 43956 19329
rect 44088 19320 44140 19372
rect 43168 19252 43220 19304
rect 43260 19252 43312 19304
rect 45376 19295 45428 19304
rect 45376 19261 45385 19295
rect 45385 19261 45419 19295
rect 45419 19261 45428 19295
rect 45376 19252 45428 19261
rect 45836 19295 45888 19304
rect 45836 19261 45845 19295
rect 45845 19261 45879 19295
rect 45879 19261 45888 19295
rect 45836 19252 45888 19261
rect 20536 19116 20588 19168
rect 20812 19159 20864 19168
rect 20812 19125 20821 19159
rect 20821 19125 20855 19159
rect 20855 19125 20864 19159
rect 20812 19116 20864 19125
rect 22008 19116 22060 19168
rect 25228 19116 25280 19168
rect 25688 19116 25740 19168
rect 46848 19184 46900 19236
rect 47584 19227 47636 19236
rect 47584 19193 47593 19227
rect 47593 19193 47627 19227
rect 47627 19193 47636 19227
rect 47584 19184 47636 19193
rect 43168 19116 43220 19168
rect 43996 19116 44048 19168
rect 47952 19363 48004 19372
rect 47952 19329 47961 19363
rect 47961 19329 47995 19363
rect 47995 19329 48004 19363
rect 47952 19320 48004 19329
rect 48044 19252 48096 19304
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 3240 18912 3292 18964
rect 18512 18887 18564 18896
rect 18512 18853 18521 18887
rect 18521 18853 18555 18887
rect 18555 18853 18564 18887
rect 18512 18844 18564 18853
rect 20904 18844 20956 18896
rect 21180 18844 21232 18896
rect 27160 18844 27212 18896
rect 28724 18887 28776 18896
rect 28724 18853 28733 18887
rect 28733 18853 28767 18887
rect 28767 18853 28776 18887
rect 28724 18844 28776 18853
rect 14004 18776 14056 18828
rect 14924 18776 14976 18828
rect 2320 18708 2372 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 13912 18708 13964 18760
rect 20168 18776 20220 18828
rect 16764 18708 16816 18760
rect 18972 18708 19024 18760
rect 20536 18751 20588 18760
rect 20536 18717 20545 18751
rect 20545 18717 20579 18751
rect 20579 18717 20588 18751
rect 20536 18708 20588 18717
rect 21088 18776 21140 18828
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 25504 18819 25556 18828
rect 25504 18785 25513 18819
rect 25513 18785 25547 18819
rect 25547 18785 25556 18819
rect 25504 18776 25556 18785
rect 30472 18819 30524 18828
rect 30472 18785 30481 18819
rect 30481 18785 30515 18819
rect 30515 18785 30524 18819
rect 30472 18776 30524 18785
rect 45376 18912 45428 18964
rect 47584 18912 47636 18964
rect 48044 18912 48096 18964
rect 21180 18751 21232 18760
rect 21180 18717 21189 18751
rect 21189 18717 21223 18751
rect 21223 18717 21232 18751
rect 21180 18708 21232 18717
rect 23664 18751 23716 18760
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 23664 18708 23716 18717
rect 24308 18708 24360 18760
rect 27988 18751 28040 18760
rect 27988 18717 27997 18751
rect 27997 18717 28031 18751
rect 28031 18717 28040 18751
rect 27988 18708 28040 18717
rect 28172 18751 28224 18760
rect 28172 18717 28181 18751
rect 28181 18717 28215 18751
rect 28215 18717 28224 18751
rect 28172 18708 28224 18717
rect 28908 18751 28960 18760
rect 28908 18717 28917 18751
rect 28917 18717 28951 18751
rect 28951 18717 28960 18751
rect 28908 18708 28960 18717
rect 29644 18751 29696 18760
rect 29644 18717 29653 18751
rect 29653 18717 29687 18751
rect 29687 18717 29696 18751
rect 29644 18708 29696 18717
rect 40500 18751 40552 18760
rect 40500 18717 40509 18751
rect 40509 18717 40543 18751
rect 40543 18717 40552 18751
rect 40500 18708 40552 18717
rect 40684 18751 40736 18760
rect 40684 18717 40693 18751
rect 40693 18717 40727 18751
rect 40727 18717 40736 18751
rect 40684 18708 40736 18717
rect 41696 18708 41748 18760
rect 48136 18819 48188 18828
rect 43260 18708 43312 18760
rect 15108 18640 15160 18692
rect 16028 18640 16080 18692
rect 22100 18640 22152 18692
rect 24400 18683 24452 18692
rect 24400 18649 24409 18683
rect 24409 18649 24443 18683
rect 24443 18649 24452 18683
rect 24400 18640 24452 18649
rect 27068 18640 27120 18692
rect 28264 18683 28316 18692
rect 28264 18649 28273 18683
rect 28273 18649 28307 18683
rect 28307 18649 28316 18683
rect 28264 18640 28316 18649
rect 29828 18683 29880 18692
rect 29828 18649 29837 18683
rect 29837 18649 29871 18683
rect 29871 18649 29880 18683
rect 29828 18640 29880 18649
rect 13728 18572 13780 18624
rect 14280 18572 14332 18624
rect 14740 18572 14792 18624
rect 16396 18572 16448 18624
rect 23020 18572 23072 18624
rect 24676 18572 24728 18624
rect 24952 18572 25004 18624
rect 41052 18572 41104 18624
rect 42708 18572 42760 18624
rect 43812 18708 43864 18760
rect 43996 18751 44048 18760
rect 43996 18717 44005 18751
rect 44005 18717 44039 18751
rect 44039 18717 44048 18751
rect 43996 18708 44048 18717
rect 44180 18751 44232 18760
rect 44180 18717 44189 18751
rect 44189 18717 44223 18751
rect 44223 18717 44232 18751
rect 44180 18708 44232 18717
rect 45008 18751 45060 18760
rect 43720 18640 43772 18692
rect 45008 18717 45017 18751
rect 45017 18717 45051 18751
rect 45051 18717 45060 18751
rect 45008 18708 45060 18717
rect 45284 18708 45336 18760
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 47676 18640 47728 18692
rect 47216 18572 47268 18624
rect 47952 18572 48004 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 29460 18368 29512 18420
rect 29828 18368 29880 18420
rect 14280 18343 14332 18352
rect 14280 18309 14289 18343
rect 14289 18309 14323 18343
rect 14323 18309 14332 18343
rect 14280 18300 14332 18309
rect 15108 18343 15160 18352
rect 15108 18309 15117 18343
rect 15117 18309 15151 18343
rect 15151 18309 15160 18343
rect 15108 18300 15160 18309
rect 21180 18300 21232 18352
rect 22100 18300 22152 18352
rect 24860 18300 24912 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 14464 18275 14516 18284
rect 14464 18241 14473 18275
rect 14473 18241 14507 18275
rect 14507 18241 14516 18275
rect 14464 18232 14516 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 14924 18232 14976 18284
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 2872 18164 2924 18216
rect 2964 18207 3016 18216
rect 2964 18173 2973 18207
rect 2973 18173 3007 18207
rect 3007 18173 3016 18207
rect 2964 18164 3016 18173
rect 14832 18164 14884 18216
rect 15108 18164 15160 18216
rect 16028 18164 16080 18216
rect 18420 18232 18472 18284
rect 20904 18232 20956 18284
rect 20996 18232 21048 18284
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 24676 18232 24728 18284
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 20444 18207 20496 18216
rect 20444 18173 20453 18207
rect 20453 18173 20487 18207
rect 20487 18173 20496 18207
rect 20444 18164 20496 18173
rect 21180 18164 21232 18216
rect 23204 18164 23256 18216
rect 27620 18275 27672 18284
rect 27620 18241 27629 18275
rect 27629 18241 27663 18275
rect 27663 18241 27672 18275
rect 27620 18232 27672 18241
rect 28264 18275 28316 18284
rect 28264 18241 28273 18275
rect 28273 18241 28307 18275
rect 28307 18241 28316 18275
rect 28264 18232 28316 18241
rect 30380 18300 30432 18352
rect 44180 18368 44232 18420
rect 47676 18411 47728 18420
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 32404 18232 32456 18284
rect 45652 18300 45704 18352
rect 45836 18343 45888 18352
rect 45836 18309 45845 18343
rect 45845 18309 45879 18343
rect 45879 18309 45888 18343
rect 45836 18300 45888 18309
rect 40500 18232 40552 18284
rect 40684 18232 40736 18284
rect 40960 18232 41012 18284
rect 42708 18275 42760 18284
rect 42708 18241 42717 18275
rect 42717 18241 42751 18275
rect 42751 18241 42760 18275
rect 42708 18232 42760 18241
rect 41052 18164 41104 18216
rect 43720 18232 43772 18284
rect 46848 18275 46900 18284
rect 46848 18241 46857 18275
rect 46857 18241 46891 18275
rect 46891 18241 46900 18275
rect 46848 18232 46900 18241
rect 47216 18232 47268 18284
rect 43444 18207 43496 18216
rect 29644 18096 29696 18148
rect 43444 18173 43453 18207
rect 43453 18173 43487 18207
rect 43487 18173 43496 18207
rect 43444 18164 43496 18173
rect 43996 18207 44048 18216
rect 43996 18173 44005 18207
rect 44005 18173 44039 18207
rect 44039 18173 44048 18207
rect 43996 18164 44048 18173
rect 44180 18207 44232 18216
rect 44180 18173 44189 18207
rect 44189 18173 44223 18207
rect 44223 18173 44232 18207
rect 44180 18164 44232 18173
rect 13360 18028 13412 18080
rect 16672 18028 16724 18080
rect 30748 18028 30800 18080
rect 32404 18028 32456 18080
rect 41328 18028 41380 18080
rect 44088 18096 44140 18148
rect 46940 18071 46992 18080
rect 46940 18037 46949 18071
rect 46949 18037 46983 18071
rect 46983 18037 46992 18071
rect 46940 18028 46992 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 14096 17824 14148 17876
rect 14832 17824 14884 17876
rect 21456 17867 21508 17876
rect 21456 17833 21465 17867
rect 21465 17833 21499 17867
rect 21499 17833 21508 17867
rect 21456 17824 21508 17833
rect 24308 17824 24360 17876
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 2872 17620 2924 17672
rect 28816 17688 28868 17740
rect 30748 17731 30800 17740
rect 30748 17697 30757 17731
rect 30757 17697 30791 17731
rect 30791 17697 30800 17731
rect 30748 17688 30800 17697
rect 41328 17824 41380 17876
rect 41052 17799 41104 17808
rect 41052 17765 41061 17799
rect 41061 17765 41095 17799
rect 41095 17765 41104 17799
rect 41052 17756 41104 17765
rect 41696 17731 41748 17740
rect 41696 17697 41705 17731
rect 41705 17697 41739 17731
rect 41739 17697 41748 17731
rect 41696 17688 41748 17697
rect 14832 17663 14884 17672
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 16396 17663 16448 17672
rect 14832 17620 14884 17629
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 22928 17620 22980 17672
rect 26884 17620 26936 17672
rect 27620 17663 27672 17672
rect 27620 17629 27629 17663
rect 27629 17629 27663 17663
rect 27663 17629 27672 17663
rect 27620 17620 27672 17629
rect 27988 17663 28040 17672
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 28172 17620 28224 17672
rect 28632 17663 28684 17672
rect 28632 17629 28641 17663
rect 28641 17629 28675 17663
rect 28675 17629 28684 17663
rect 28632 17620 28684 17629
rect 43904 17824 43956 17876
rect 42248 17799 42300 17808
rect 42248 17765 42257 17799
rect 42257 17765 42291 17799
rect 42291 17765 42300 17799
rect 44180 17799 44232 17808
rect 42248 17756 42300 17765
rect 44180 17765 44189 17799
rect 44189 17765 44223 17799
rect 44223 17765 44232 17799
rect 44180 17756 44232 17765
rect 43720 17688 43772 17740
rect 15200 17552 15252 17604
rect 16764 17552 16816 17604
rect 18236 17595 18288 17604
rect 18236 17561 18245 17595
rect 18245 17561 18279 17595
rect 18279 17561 18288 17595
rect 18236 17552 18288 17561
rect 21180 17595 21232 17604
rect 21180 17561 21189 17595
rect 21189 17561 21223 17595
rect 21223 17561 21232 17595
rect 21180 17552 21232 17561
rect 23020 17552 23072 17604
rect 43812 17663 43864 17672
rect 43812 17629 43821 17663
rect 43821 17629 43855 17663
rect 43855 17629 43864 17663
rect 43812 17620 43864 17629
rect 46940 17688 46992 17740
rect 44272 17663 44324 17672
rect 44272 17629 44281 17663
rect 44281 17629 44315 17663
rect 44315 17629 44324 17663
rect 44272 17620 44324 17629
rect 45008 17663 45060 17672
rect 45008 17629 45017 17663
rect 45017 17629 45051 17663
rect 45051 17629 45060 17663
rect 45008 17620 45060 17629
rect 46296 17663 46348 17672
rect 46296 17629 46305 17663
rect 46305 17629 46339 17663
rect 46339 17629 46348 17663
rect 46296 17620 46348 17629
rect 32404 17595 32456 17604
rect 1952 17484 2004 17536
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 32404 17561 32413 17595
rect 32413 17561 32447 17595
rect 32447 17561 32456 17595
rect 32404 17552 32456 17561
rect 40960 17484 41012 17536
rect 41236 17527 41288 17536
rect 41236 17493 41245 17527
rect 41245 17493 41279 17527
rect 41279 17493 41288 17527
rect 41236 17484 41288 17493
rect 45284 17552 45336 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 42616 17484 42668 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 16764 17323 16816 17332
rect 16764 17289 16773 17323
rect 16773 17289 16807 17323
rect 16807 17289 16816 17323
rect 16764 17280 16816 17289
rect 1952 17255 2004 17264
rect 1952 17221 1961 17255
rect 1961 17221 1995 17255
rect 1995 17221 2004 17255
rect 1952 17212 2004 17221
rect 15200 17212 15252 17264
rect 24308 17280 24360 17332
rect 24768 17280 24820 17332
rect 27620 17280 27672 17332
rect 32404 17280 32456 17332
rect 41788 17280 41840 17332
rect 22192 17212 22244 17264
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 21180 17144 21232 17196
rect 22928 17187 22980 17196
rect 22928 17153 22937 17187
rect 22937 17153 22971 17187
rect 22971 17153 22980 17187
rect 22928 17144 22980 17153
rect 23296 17144 23348 17196
rect 24308 17144 24360 17196
rect 24952 17144 25004 17196
rect 26240 17212 26292 17264
rect 2044 17076 2096 17128
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 3516 17076 3568 17128
rect 9036 17076 9088 17128
rect 14832 17076 14884 17128
rect 17684 17008 17736 17060
rect 21088 17008 21140 17060
rect 22008 17008 22060 17060
rect 24400 17076 24452 17128
rect 24584 17076 24636 17128
rect 25964 17144 26016 17196
rect 26884 17144 26936 17196
rect 27160 17144 27212 17196
rect 42616 17187 42668 17196
rect 42616 17153 42625 17187
rect 42625 17153 42659 17187
rect 42659 17153 42668 17187
rect 42616 17144 42668 17153
rect 41236 17076 41288 17128
rect 46388 17076 46440 17128
rect 46848 17119 46900 17128
rect 46848 17085 46857 17119
rect 46857 17085 46891 17119
rect 46891 17085 46900 17119
rect 46848 17076 46900 17085
rect 14096 16940 14148 16992
rect 15384 16940 15436 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 25044 17008 25096 17060
rect 42984 17051 43036 17060
rect 42984 17017 42993 17051
rect 42993 17017 43027 17051
rect 43027 17017 43036 17051
rect 42984 17008 43036 17017
rect 44548 17008 44600 17060
rect 45468 17008 45520 17060
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 24676 16940 24728 16992
rect 26056 16983 26108 16992
rect 26056 16949 26065 16983
rect 26065 16949 26099 16983
rect 26099 16949 26108 16983
rect 26056 16940 26108 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 14556 16736 14608 16788
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 17408 16600 17460 16652
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 17960 16643 18012 16652
rect 17960 16609 17969 16643
rect 17969 16609 18003 16643
rect 18003 16609 18012 16643
rect 17960 16600 18012 16609
rect 21088 16736 21140 16788
rect 24400 16736 24452 16788
rect 28632 16736 28684 16788
rect 46296 16736 46348 16788
rect 24676 16668 24728 16720
rect 24768 16668 24820 16720
rect 22100 16600 22152 16652
rect 25044 16643 25096 16652
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 27160 16600 27212 16652
rect 42984 16600 43036 16652
rect 43996 16600 44048 16652
rect 45468 16643 45520 16652
rect 45468 16609 45477 16643
rect 45477 16609 45511 16643
rect 45511 16609 45520 16643
rect 45468 16600 45520 16609
rect 17868 16532 17920 16584
rect 18420 16575 18472 16584
rect 18420 16541 18429 16575
rect 18429 16541 18463 16575
rect 18463 16541 18472 16575
rect 18420 16532 18472 16541
rect 19432 16532 19484 16584
rect 21456 16532 21508 16584
rect 24584 16532 24636 16584
rect 24952 16575 25004 16584
rect 24952 16541 24961 16575
rect 24961 16541 24995 16575
rect 24995 16541 25004 16575
rect 27068 16575 27120 16584
rect 24952 16532 25004 16541
rect 27068 16541 27077 16575
rect 27077 16541 27111 16575
rect 27111 16541 27120 16575
rect 27068 16532 27120 16541
rect 44548 16532 44600 16584
rect 14372 16507 14424 16516
rect 14372 16473 14381 16507
rect 14381 16473 14415 16507
rect 14415 16473 14424 16507
rect 14372 16464 14424 16473
rect 15384 16464 15436 16516
rect 18236 16464 18288 16516
rect 15200 16396 15252 16448
rect 18604 16439 18656 16448
rect 18604 16405 18613 16439
rect 18613 16405 18647 16439
rect 18647 16405 18656 16439
rect 18604 16396 18656 16405
rect 19340 16439 19392 16448
rect 19340 16405 19349 16439
rect 19349 16405 19383 16439
rect 19383 16405 19392 16439
rect 19340 16396 19392 16405
rect 21824 16439 21876 16448
rect 21824 16405 21833 16439
rect 21833 16405 21867 16439
rect 21867 16405 21876 16439
rect 21824 16396 21876 16405
rect 23848 16439 23900 16448
rect 23848 16405 23857 16439
rect 23857 16405 23891 16439
rect 23891 16405 23900 16439
rect 23848 16396 23900 16405
rect 24216 16464 24268 16516
rect 45560 16396 45612 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 18420 16192 18472 16244
rect 15016 16124 15068 16176
rect 15108 16056 15160 16108
rect 17960 16124 18012 16176
rect 19340 16124 19392 16176
rect 14372 15988 14424 16040
rect 16672 16056 16724 16108
rect 20352 16192 20404 16244
rect 23296 16235 23348 16244
rect 21364 16124 21416 16176
rect 23296 16201 23305 16235
rect 23305 16201 23339 16235
rect 23339 16201 23348 16235
rect 23296 16192 23348 16201
rect 25044 16192 25096 16244
rect 20996 16056 21048 16108
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 21916 16056 21968 16108
rect 17592 15988 17644 16040
rect 18604 15988 18656 16040
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 22100 15988 22152 15997
rect 14464 15920 14516 15972
rect 15108 15920 15160 15972
rect 14924 15852 14976 15904
rect 15016 15852 15068 15904
rect 17868 15852 17920 15904
rect 19616 15852 19668 15904
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 22100 15852 22152 15904
rect 25320 16124 25372 16176
rect 23848 16056 23900 16108
rect 41236 16099 41288 16108
rect 41236 16065 41245 16099
rect 41245 16065 41279 16099
rect 41279 16065 41288 16099
rect 41236 16056 41288 16065
rect 46388 16056 46440 16108
rect 24216 15988 24268 16040
rect 24400 16031 24452 16040
rect 24400 15997 24409 16031
rect 24409 15997 24443 16031
rect 24443 15997 24452 16031
rect 24400 15988 24452 15997
rect 23572 15852 23624 15904
rect 41420 15852 41472 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 22284 15648 22336 15700
rect 23572 15691 23624 15700
rect 23572 15657 23581 15691
rect 23581 15657 23615 15691
rect 23615 15657 23624 15691
rect 23572 15648 23624 15657
rect 24400 15691 24452 15700
rect 24400 15657 24409 15691
rect 24409 15657 24443 15691
rect 24443 15657 24452 15691
rect 24400 15648 24452 15657
rect 25320 15691 25372 15700
rect 25320 15657 25329 15691
rect 25329 15657 25363 15691
rect 25363 15657 25372 15691
rect 25320 15648 25372 15657
rect 21364 15623 21416 15632
rect 21364 15589 21373 15623
rect 21373 15589 21407 15623
rect 21407 15589 21416 15623
rect 21364 15580 21416 15589
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 19616 15555 19668 15564
rect 19616 15521 19625 15555
rect 19625 15521 19659 15555
rect 19659 15521 19668 15555
rect 19616 15512 19668 15521
rect 20904 15512 20956 15564
rect 21824 15555 21876 15564
rect 21824 15521 21833 15555
rect 21833 15521 21867 15555
rect 21867 15521 21876 15555
rect 21824 15512 21876 15521
rect 22100 15555 22152 15564
rect 22100 15521 22109 15555
rect 22109 15521 22143 15555
rect 22143 15521 22152 15555
rect 22100 15512 22152 15521
rect 43444 15580 43496 15632
rect 41420 15555 41472 15564
rect 41420 15521 41429 15555
rect 41429 15521 41463 15555
rect 41463 15521 41472 15555
rect 42892 15555 42944 15564
rect 41420 15512 41472 15521
rect 42892 15521 42901 15555
rect 42901 15521 42935 15555
rect 42935 15521 42944 15555
rect 42892 15512 42944 15521
rect 1768 15444 1820 15496
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 14740 15444 14792 15453
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 14924 15376 14976 15428
rect 16672 15308 16724 15360
rect 17868 15376 17920 15428
rect 21180 15376 21232 15428
rect 23112 15376 23164 15428
rect 18052 15308 18104 15360
rect 21456 15308 21508 15360
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 26056 15444 26108 15496
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 14740 15104 14792 15156
rect 17408 15147 17460 15156
rect 17408 15113 17433 15147
rect 17433 15113 17460 15147
rect 17592 15147 17644 15156
rect 17408 15104 17460 15113
rect 17592 15113 17601 15147
rect 17601 15113 17635 15147
rect 17635 15113 17644 15147
rect 17592 15104 17644 15113
rect 21180 15147 21232 15156
rect 21180 15113 21189 15147
rect 21189 15113 21223 15147
rect 21223 15113 21232 15147
rect 21180 15104 21232 15113
rect 23112 15104 23164 15156
rect 17776 15036 17828 15088
rect 21364 15036 21416 15088
rect 21824 15079 21876 15088
rect 21824 15045 21833 15079
rect 21833 15045 21867 15079
rect 21867 15045 21876 15079
rect 21824 15036 21876 15045
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 14556 14968 14608 15020
rect 18052 15011 18104 15020
rect 18052 14977 18061 15011
rect 18061 14977 18095 15011
rect 18095 14977 18104 15011
rect 18052 14968 18104 14977
rect 19432 14968 19484 15020
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 18328 14943 18380 14952
rect 2780 14900 2832 14909
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 19340 14900 19392 14952
rect 21916 14968 21968 15020
rect 22192 14968 22244 15020
rect 25228 14968 25280 15020
rect 17868 14832 17920 14884
rect 20996 14832 21048 14884
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 18328 14560 18380 14612
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 2872 14356 2924 14408
rect 17408 14492 17460 14544
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 19340 14399 19392 14408
rect 19340 14365 19349 14399
rect 19349 14365 19383 14399
rect 19383 14365 19392 14399
rect 19340 14356 19392 14365
rect 22560 14356 22612 14408
rect 30564 14356 30616 14408
rect 17868 14288 17920 14340
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 22928 14263 22980 14272
rect 22928 14229 22937 14263
rect 22937 14229 22971 14263
rect 22971 14229 22980 14263
rect 22928 14220 22980 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 3700 13948 3752 14000
rect 15108 13880 15160 13932
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 3976 13744 4028 13796
rect 14280 13744 14332 13796
rect 21824 13948 21876 14000
rect 22928 13948 22980 14000
rect 45100 13880 45152 13932
rect 46940 13719 46992 13728
rect 46940 13685 46949 13719
rect 46949 13685 46983 13719
rect 46983 13685 46992 13719
rect 46940 13676 46992 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 15844 13472 15896 13524
rect 24860 13472 24912 13524
rect 17776 13404 17828 13456
rect 16948 13379 17000 13388
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 17960 13336 18012 13388
rect 30472 13404 30524 13456
rect 22468 13379 22520 13388
rect 22468 13345 22477 13379
rect 22477 13345 22511 13379
rect 22511 13345 22520 13379
rect 22468 13336 22520 13345
rect 46940 13336 46992 13388
rect 17868 13268 17920 13320
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 46296 13311 46348 13320
rect 46296 13277 46305 13311
rect 46305 13277 46339 13311
rect 46339 13277 46348 13311
rect 46296 13268 46348 13277
rect 22192 13243 22244 13252
rect 22192 13209 22201 13243
rect 22201 13209 22235 13243
rect 22235 13209 22244 13243
rect 22192 13200 22244 13209
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 16764 13132 16816 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3332 12928 3384 12980
rect 22468 12928 22520 12980
rect 15844 12860 15896 12912
rect 22284 12860 22336 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 46296 12792 46348 12844
rect 16580 12724 16632 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 3516 12656 3568 12708
rect 14832 12588 14884 12640
rect 16948 12588 17000 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 16856 12384 16908 12436
rect 17960 12384 18012 12436
rect 22192 12384 22244 12436
rect 16764 12180 16816 12232
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 46940 11024 46992 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 3424 10956 3476 11008
rect 10784 10956 10836 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 46940 10795 46992 10804
rect 46940 10761 46949 10795
rect 46949 10761 46983 10795
rect 46983 10761 46992 10795
rect 46940 10752 46992 10761
rect 45652 10616 45704 10668
rect 46664 10616 46716 10668
rect 47584 10659 47636 10668
rect 47584 10625 47593 10659
rect 47593 10625 47627 10659
rect 47627 10625 47636 10659
rect 47584 10616 47636 10625
rect 46296 10412 46348 10464
rect 46480 10412 46532 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 46480 10115 46532 10124
rect 46480 10081 46489 10115
rect 46489 10081 46523 10115
rect 46523 10081 46532 10115
rect 46480 10072 46532 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 46112 9392 46164 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47768 8891 47820 8900
rect 47768 8857 47777 8891
rect 47777 8857 47811 8891
rect 47811 8857 47820 8891
rect 47768 8848 47820 8857
rect 29736 8780 29788 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 45100 8483 45152 8492
rect 45100 8449 45109 8483
rect 45109 8449 45143 8483
rect 45143 8449 45152 8483
rect 45100 8440 45152 8449
rect 3424 8236 3476 8288
rect 18052 8236 18104 8288
rect 18512 8236 18564 8288
rect 45284 8236 45336 8288
rect 45560 8236 45612 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1860 8032 1912 8084
rect 45100 8032 45152 8084
rect 45376 7896 45428 7948
rect 47676 7896 47728 7948
rect 44824 7828 44876 7880
rect 47308 7871 47360 7880
rect 47308 7837 47317 7871
rect 47317 7837 47351 7871
rect 47351 7837 47360 7871
rect 47308 7828 47360 7837
rect 45192 7803 45244 7812
rect 45192 7769 45201 7803
rect 45201 7769 45235 7803
rect 45235 7769 45244 7803
rect 45192 7760 45244 7769
rect 45284 7803 45336 7812
rect 45284 7769 45293 7803
rect 45293 7769 45327 7803
rect 45327 7769 45336 7803
rect 45284 7760 45336 7769
rect 16856 7692 16908 7744
rect 32496 7692 32548 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 45192 7488 45244 7540
rect 44824 7463 44876 7472
rect 44824 7429 44833 7463
rect 44833 7429 44867 7463
rect 44867 7429 44876 7463
rect 44824 7420 44876 7429
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 42892 7284 42944 7336
rect 45376 7284 45428 7336
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 43076 6400 43128 6452
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 15568 6196 15620 6248
rect 32220 6196 32272 6248
rect 3240 6128 3292 6180
rect 28448 6128 28500 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 40224 5695 40276 5704
rect 40224 5661 40233 5695
rect 40233 5661 40267 5695
rect 40267 5661 40276 5695
rect 40224 5652 40276 5661
rect 43536 5652 43588 5704
rect 40316 5559 40368 5568
rect 40316 5525 40325 5559
rect 40325 5525 40359 5559
rect 40359 5525 40368 5559
rect 40316 5516 40368 5525
rect 42616 5559 42668 5568
rect 42616 5525 42625 5559
rect 42625 5525 42659 5559
rect 42659 5525 42668 5559
rect 42616 5516 42668 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3976 5312 4028 5364
rect 6644 5244 6696 5296
rect 18696 5219 18748 5228
rect 18696 5185 18705 5219
rect 18705 5185 18739 5219
rect 18739 5185 18748 5219
rect 18696 5176 18748 5185
rect 36544 5244 36596 5296
rect 38476 5244 38528 5296
rect 40224 5312 40276 5364
rect 42616 5287 42668 5296
rect 40316 5176 40368 5228
rect 40776 5176 40828 5228
rect 40960 5219 41012 5228
rect 40960 5185 40969 5219
rect 40969 5185 41003 5219
rect 41003 5185 41012 5219
rect 40960 5176 41012 5185
rect 42616 5253 42625 5287
rect 42625 5253 42659 5287
rect 42659 5253 42668 5287
rect 42616 5244 42668 5253
rect 44364 5244 44416 5296
rect 47860 5219 47912 5228
rect 47860 5185 47869 5219
rect 47869 5185 47903 5219
rect 47903 5185 47912 5219
rect 47860 5176 47912 5185
rect 25596 5040 25648 5092
rect 19248 4972 19300 5024
rect 39764 5015 39816 5024
rect 39764 4981 39773 5015
rect 39773 4981 39807 5015
rect 39807 4981 39816 5015
rect 39764 4972 39816 4981
rect 40500 4972 40552 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 40224 4768 40276 4820
rect 46572 4768 46624 4820
rect 18880 4700 18932 4752
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 19340 4607 19392 4616
rect 19340 4573 19349 4607
rect 19349 4573 19383 4607
rect 19383 4573 19392 4607
rect 19340 4564 19392 4573
rect 20628 4607 20680 4616
rect 20628 4573 20637 4607
rect 20637 4573 20671 4607
rect 20671 4573 20680 4607
rect 20628 4564 20680 4573
rect 22192 4632 22244 4684
rect 25596 4675 25648 4684
rect 25596 4641 25605 4675
rect 25605 4641 25639 4675
rect 25639 4641 25648 4675
rect 25596 4632 25648 4641
rect 27252 4675 27304 4684
rect 27252 4641 27261 4675
rect 27261 4641 27295 4675
rect 27295 4641 27304 4675
rect 27252 4632 27304 4641
rect 39764 4632 39816 4684
rect 40500 4675 40552 4684
rect 40500 4641 40509 4675
rect 40509 4641 40543 4675
rect 40543 4641 40552 4675
rect 40500 4632 40552 4641
rect 42156 4675 42208 4684
rect 42156 4641 42165 4675
rect 42165 4641 42199 4675
rect 42199 4641 42208 4675
rect 42156 4632 42208 4641
rect 42892 4675 42944 4684
rect 42892 4641 42901 4675
rect 42901 4641 42935 4675
rect 42935 4641 42944 4675
rect 42892 4632 42944 4641
rect 44364 4632 44416 4684
rect 44824 4632 44876 4684
rect 22560 4564 22612 4616
rect 23756 4564 23808 4616
rect 46664 4607 46716 4616
rect 22468 4496 22520 4548
rect 18144 4471 18196 4480
rect 18144 4437 18153 4471
rect 18153 4437 18187 4471
rect 18187 4437 18196 4471
rect 18144 4428 18196 4437
rect 20352 4428 20404 4480
rect 20996 4428 21048 4480
rect 22284 4428 22336 4480
rect 22744 4471 22796 4480
rect 22744 4437 22753 4471
rect 22753 4437 22787 4471
rect 22787 4437 22796 4471
rect 22744 4428 22796 4437
rect 25320 4428 25372 4480
rect 46664 4573 46673 4607
rect 46673 4573 46707 4607
rect 46707 4573 46716 4607
rect 46664 4564 46716 4573
rect 46848 4564 46900 4616
rect 39488 4496 39540 4548
rect 42892 4496 42944 4548
rect 43076 4496 43128 4548
rect 32128 4428 32180 4480
rect 46480 4428 46532 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 19340 4224 19392 4276
rect 20628 4224 20680 4276
rect 38384 4224 38436 4276
rect 13728 4131 13780 4140
rect 2964 4020 3016 4072
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 7380 4063 7432 4072
rect 3056 4020 3108 4029
rect 7380 4029 7389 4063
rect 7389 4029 7423 4063
rect 7423 4029 7432 4063
rect 7380 4020 7432 4029
rect 7564 4063 7616 4072
rect 7564 4029 7573 4063
rect 7573 4029 7607 4063
rect 7607 4029 7616 4063
rect 7564 4020 7616 4029
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 17040 4088 17092 4140
rect 17500 4088 17552 4140
rect 17776 4088 17828 4140
rect 3976 3952 4028 4004
rect 7104 3952 7156 4004
rect 16028 4020 16080 4072
rect 18696 4020 18748 4072
rect 19340 4088 19392 4140
rect 19708 4131 19760 4140
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 21548 4088 21600 4140
rect 22468 4131 22520 4140
rect 22468 4097 22477 4131
rect 22477 4097 22511 4131
rect 22511 4097 22520 4131
rect 22468 4088 22520 4097
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 22560 4088 22612 4097
rect 20536 4020 20588 4072
rect 20720 4020 20772 4072
rect 12072 3952 12124 4004
rect 18604 3952 18656 4004
rect 18788 3952 18840 4004
rect 26700 4088 26752 4140
rect 27344 4088 27396 4140
rect 31668 4088 31720 4140
rect 36636 4088 36688 4140
rect 36912 4088 36964 4140
rect 37648 4156 37700 4208
rect 38476 4199 38528 4208
rect 38476 4165 38485 4199
rect 38485 4165 38519 4199
rect 38519 4165 38528 4199
rect 38476 4156 38528 4165
rect 40592 4199 40644 4208
rect 40592 4165 40601 4199
rect 40601 4165 40635 4199
rect 40635 4165 40644 4199
rect 40592 4156 40644 4165
rect 40776 4224 40828 4276
rect 41236 4156 41288 4208
rect 47768 4199 47820 4208
rect 47768 4165 47777 4199
rect 47777 4165 47811 4199
rect 47811 4165 47820 4199
rect 47768 4156 47820 4165
rect 40868 4088 40920 4140
rect 46756 4131 46808 4140
rect 46756 4097 46765 4131
rect 46765 4097 46799 4131
rect 46799 4097 46808 4131
rect 46756 4088 46808 4097
rect 32128 3952 32180 4004
rect 36176 3952 36228 4004
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 11520 3884 11572 3936
rect 14004 3884 14056 3936
rect 17960 3927 18012 3936
rect 17960 3893 17969 3927
rect 17969 3893 18003 3927
rect 18003 3893 18012 3927
rect 17960 3884 18012 3893
rect 18512 3884 18564 3936
rect 20812 3884 20864 3936
rect 22100 3884 22152 3936
rect 23112 3884 23164 3936
rect 26240 3884 26292 3936
rect 27528 3884 27580 3936
rect 32772 3884 32824 3936
rect 36268 3884 36320 3936
rect 38384 4020 38436 4072
rect 39488 4063 39540 4072
rect 39488 4029 39497 4063
rect 39497 4029 39531 4063
rect 39531 4029 39540 4063
rect 39488 4020 39540 4029
rect 39672 4063 39724 4072
rect 39672 4029 39681 4063
rect 39681 4029 39715 4063
rect 39715 4029 39724 4063
rect 39672 4020 39724 4029
rect 39948 4020 40000 4072
rect 47216 4020 47268 4072
rect 36544 3995 36596 4004
rect 36544 3961 36553 3995
rect 36553 3961 36587 3995
rect 36587 3961 36596 3995
rect 36544 3952 36596 3961
rect 40132 3927 40184 3936
rect 40132 3893 40141 3927
rect 40141 3893 40175 3927
rect 40175 3893 40184 3927
rect 40132 3884 40184 3893
rect 40408 3884 40460 3936
rect 42800 3884 42852 3936
rect 42984 3884 43036 3936
rect 43812 3927 43864 3936
rect 43812 3893 43821 3927
rect 43821 3893 43855 3927
rect 43855 3893 43864 3927
rect 43812 3884 43864 3893
rect 46296 3927 46348 3936
rect 46296 3893 46305 3927
rect 46305 3893 46339 3927
rect 46339 3893 46348 3927
rect 46296 3884 46348 3893
rect 46940 3927 46992 3936
rect 46940 3893 46949 3927
rect 46949 3893 46983 3927
rect 46983 3893 46992 3927
rect 46940 3884 46992 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 19708 3680 19760 3732
rect 20260 3680 20312 3732
rect 21548 3723 21600 3732
rect 21548 3689 21557 3723
rect 21557 3689 21591 3723
rect 21591 3689 21600 3723
rect 21548 3680 21600 3689
rect 22192 3723 22244 3732
rect 22192 3689 22201 3723
rect 22201 3689 22235 3723
rect 22235 3689 22244 3723
rect 22192 3680 22244 3689
rect 23664 3680 23716 3732
rect 25136 3680 25188 3732
rect 6460 3587 6512 3596
rect 1768 3476 1820 3528
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 9496 3544 9548 3596
rect 9588 3544 9640 3596
rect 13728 3612 13780 3664
rect 18420 3612 18472 3664
rect 18696 3612 18748 3664
rect 27344 3680 27396 3732
rect 32680 3680 32732 3732
rect 32772 3680 32824 3732
rect 39304 3612 39356 3664
rect 40960 3680 41012 3732
rect 41420 3680 41472 3732
rect 43536 3723 43588 3732
rect 43536 3689 43545 3723
rect 43545 3689 43579 3723
rect 43579 3689 43588 3723
rect 43536 3680 43588 3689
rect 40408 3612 40460 3664
rect 40500 3612 40552 3664
rect 46940 3612 46992 3664
rect 26608 3544 26660 3596
rect 26884 3544 26936 3596
rect 33692 3544 33744 3596
rect 33876 3544 33928 3596
rect 40224 3544 40276 3596
rect 42156 3587 42208 3596
rect 42156 3553 42165 3587
rect 42165 3553 42199 3587
rect 42199 3553 42208 3587
rect 42156 3544 42208 3553
rect 46296 3587 46348 3596
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 13820 3476 13872 3528
rect 10232 3408 10284 3460
rect 17224 3476 17276 3528
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 18604 3476 18656 3528
rect 20352 3519 20404 3528
rect 18236 3408 18288 3460
rect 18880 3408 18932 3460
rect 19708 3408 19760 3460
rect 1952 3340 2004 3392
rect 8208 3340 8260 3392
rect 11704 3340 11756 3392
rect 17684 3383 17736 3392
rect 17684 3349 17693 3383
rect 17693 3349 17727 3383
rect 17727 3349 17736 3383
rect 17684 3340 17736 3349
rect 19432 3340 19484 3392
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 22100 3519 22152 3528
rect 22100 3485 22109 3519
rect 22109 3485 22143 3519
rect 22143 3485 22152 3519
rect 22100 3476 22152 3485
rect 22928 3476 22980 3528
rect 25412 3519 25464 3528
rect 19892 3408 19944 3460
rect 25412 3485 25421 3519
rect 25421 3485 25455 3519
rect 25455 3485 25464 3519
rect 25412 3476 25464 3485
rect 27252 3519 27304 3528
rect 27252 3485 27261 3519
rect 27261 3485 27295 3519
rect 27295 3485 27304 3519
rect 27252 3476 27304 3485
rect 32680 3476 32732 3528
rect 32956 3519 33008 3528
rect 32956 3485 32965 3519
rect 32965 3485 32999 3519
rect 32999 3485 33008 3519
rect 32956 3476 33008 3485
rect 33140 3476 33192 3528
rect 37832 3476 37884 3528
rect 39948 3476 40000 3528
rect 40132 3519 40184 3528
rect 40132 3485 40141 3519
rect 40141 3485 40175 3519
rect 40175 3485 40184 3519
rect 40776 3519 40828 3528
rect 40132 3476 40184 3485
rect 40776 3485 40785 3519
rect 40785 3485 40819 3519
rect 40819 3485 40828 3519
rect 40776 3476 40828 3485
rect 43076 3519 43128 3528
rect 43076 3485 43085 3519
rect 43085 3485 43119 3519
rect 43119 3485 43128 3519
rect 43076 3476 43128 3485
rect 44548 3476 44600 3528
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 26976 3408 27028 3460
rect 33048 3451 33100 3460
rect 33048 3417 33057 3451
rect 33057 3417 33091 3451
rect 33091 3417 33100 3451
rect 33048 3408 33100 3417
rect 33876 3408 33928 3460
rect 41328 3408 41380 3460
rect 48964 3408 49016 3460
rect 26240 3340 26292 3392
rect 26332 3340 26384 3392
rect 36544 3340 36596 3392
rect 38016 3340 38068 3392
rect 40868 3340 40920 3392
rect 44088 3383 44140 3392
rect 44088 3349 44097 3383
rect 44097 3349 44131 3383
rect 44131 3349 44140 3383
rect 44088 3340 44140 3349
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3884 3136 3936 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 8208 3111 8260 3120
rect 8208 3077 8217 3111
rect 8217 3077 8251 3111
rect 8251 3077 8260 3111
rect 8208 3068 8260 3077
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 14004 3111 14056 3120
rect 14004 3077 14013 3111
rect 14013 3077 14047 3111
rect 14047 3077 14056 3111
rect 14004 3068 14056 3077
rect 17776 3111 17828 3120
rect 17776 3077 17785 3111
rect 17785 3077 17819 3111
rect 17819 3077 17828 3111
rect 17776 3068 17828 3077
rect 18880 3111 18932 3120
rect 18880 3077 18889 3111
rect 18889 3077 18923 3111
rect 18923 3077 18932 3111
rect 18880 3068 18932 3077
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 5908 3000 5960 3052
rect 7380 3000 7432 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 17500 3000 17552 3052
rect 17684 3043 17736 3052
rect 17684 3009 17693 3043
rect 17693 3009 17727 3043
rect 17727 3009 17736 3043
rect 17684 3000 17736 3009
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 32772 3068 32824 3120
rect 33048 3111 33100 3120
rect 33048 3077 33057 3111
rect 33057 3077 33091 3111
rect 33091 3077 33100 3111
rect 33048 3068 33100 3077
rect 664 2932 716 2984
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 7748 2864 7800 2916
rect 10968 2932 11020 2984
rect 14188 2932 14240 2984
rect 15200 2932 15252 2984
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 17408 2932 17460 2984
rect 21916 3000 21968 3052
rect 22928 3043 22980 3052
rect 22928 3009 22937 3043
rect 22937 3009 22971 3043
rect 22971 3009 22980 3043
rect 22928 3000 22980 3009
rect 25596 3043 25648 3052
rect 25596 3009 25605 3043
rect 25605 3009 25639 3043
rect 25639 3009 25648 3043
rect 25596 3000 25648 3009
rect 26056 3000 26108 3052
rect 19616 2975 19668 2984
rect 19616 2941 19625 2975
rect 19625 2941 19659 2975
rect 19659 2941 19668 2975
rect 19984 2975 20036 2984
rect 19616 2932 19668 2941
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 23112 2975 23164 2984
rect 23112 2941 23121 2975
rect 23121 2941 23155 2975
rect 23155 2941 23164 2975
rect 23112 2932 23164 2941
rect 7564 2796 7616 2848
rect 9036 2796 9088 2848
rect 9588 2796 9640 2848
rect 20352 2864 20404 2916
rect 22468 2907 22520 2916
rect 22468 2873 22477 2907
rect 22477 2873 22511 2907
rect 22511 2873 22520 2907
rect 22468 2864 22520 2873
rect 22560 2864 22612 2916
rect 33140 2932 33192 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 36636 3136 36688 3188
rect 37648 3136 37700 3188
rect 38016 3111 38068 3120
rect 38016 3077 38025 3111
rect 38025 3077 38059 3111
rect 38059 3077 38068 3111
rect 38016 3068 38068 3077
rect 40776 3136 40828 3188
rect 41328 3179 41380 3188
rect 41328 3145 41337 3179
rect 41337 3145 41371 3179
rect 41371 3145 41380 3179
rect 41328 3136 41380 3145
rect 41604 3068 41656 3120
rect 37832 3043 37884 3052
rect 37832 3009 37841 3043
rect 37841 3009 37875 3043
rect 37875 3009 37884 3043
rect 37832 3000 37884 3009
rect 39304 2975 39356 2984
rect 39304 2941 39313 2975
rect 39313 2941 39347 2975
rect 39347 2941 39356 2975
rect 39304 2932 39356 2941
rect 39488 2932 39540 2984
rect 40408 2975 40460 2984
rect 40408 2941 40417 2975
rect 40417 2941 40451 2975
rect 40451 2941 40460 2975
rect 40408 2932 40460 2941
rect 41512 3043 41564 3052
rect 41512 3009 41521 3043
rect 41521 3009 41555 3043
rect 41555 3009 41564 3043
rect 43812 3136 43864 3188
rect 48044 3179 48096 3188
rect 48044 3145 48053 3179
rect 48053 3145 48087 3179
rect 48087 3145 48096 3179
rect 48044 3136 48096 3145
rect 42984 3111 43036 3120
rect 42984 3077 42993 3111
rect 42993 3077 43027 3111
rect 43027 3077 43036 3111
rect 42984 3068 43036 3077
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 41512 3000 41564 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 48320 3000 48372 3052
rect 41880 2932 41932 2984
rect 43168 2932 43220 2984
rect 47676 2932 47728 2984
rect 26056 2839 26108 2848
rect 26056 2805 26065 2839
rect 26065 2805 26099 2839
rect 26099 2805 26108 2839
rect 26056 2796 26108 2805
rect 26976 2839 27028 2848
rect 26976 2805 26985 2839
rect 26985 2805 27019 2839
rect 27019 2805 27028 2839
rect 26976 2796 27028 2805
rect 44088 2864 44140 2916
rect 35532 2796 35584 2848
rect 36176 2796 36228 2848
rect 36544 2796 36596 2848
rect 47584 2796 47636 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3240 2592 3292 2644
rect 8024 2592 8076 2644
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 18052 2592 18104 2644
rect 18236 2635 18288 2644
rect 18236 2601 18245 2635
rect 18245 2601 18279 2635
rect 18279 2601 18288 2635
rect 18236 2592 18288 2601
rect 19340 2635 19392 2644
rect 19340 2601 19349 2635
rect 19349 2601 19383 2635
rect 19383 2601 19392 2635
rect 19340 2592 19392 2601
rect 20720 2592 20772 2644
rect 21456 2592 21508 2644
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 23940 2592 23992 2644
rect 25412 2592 25464 2644
rect 28172 2592 28224 2644
rect 5172 2388 5224 2440
rect 8392 2388 8444 2440
rect 15200 2388 15252 2440
rect 1308 2320 1360 2372
rect 2596 2320 2648 2372
rect 27068 2524 27120 2576
rect 31116 2592 31168 2644
rect 35532 2635 35584 2644
rect 35532 2601 35541 2635
rect 35541 2601 35575 2635
rect 35575 2601 35584 2635
rect 35532 2592 35584 2601
rect 16120 2388 16172 2440
rect 15476 2320 15528 2372
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 17960 2388 18012 2440
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 22284 2456 22336 2508
rect 25320 2456 25372 2508
rect 33784 2524 33836 2576
rect 40592 2592 40644 2644
rect 40776 2592 40828 2644
rect 41512 2592 41564 2644
rect 35624 2456 35676 2508
rect 22468 2388 22520 2440
rect 22744 2431 22796 2440
rect 22744 2397 22753 2431
rect 22753 2397 22787 2431
rect 22787 2397 22796 2431
rect 22744 2388 22796 2397
rect 23664 2431 23716 2440
rect 23664 2397 23673 2431
rect 23673 2397 23707 2431
rect 23707 2397 23716 2431
rect 23664 2388 23716 2397
rect 20628 2320 20680 2372
rect 23204 2320 23256 2372
rect 29644 2388 29696 2440
rect 35440 2388 35492 2440
rect 24492 2320 24544 2372
rect 26424 2320 26476 2372
rect 27068 2320 27120 2372
rect 28356 2320 28408 2372
rect 31300 2320 31352 2372
rect 36360 2456 36412 2508
rect 39948 2456 40000 2508
rect 44180 2524 44232 2576
rect 42340 2456 42392 2508
rect 43076 2456 43128 2508
rect 36084 2320 36136 2372
rect 24400 2252 24452 2304
rect 26332 2295 26384 2304
rect 26332 2261 26341 2295
rect 26341 2261 26375 2295
rect 26375 2261 26384 2295
rect 26332 2252 26384 2261
rect 39672 2388 39724 2440
rect 40408 2431 40460 2440
rect 40408 2397 40417 2431
rect 40417 2397 40451 2431
rect 40451 2397 40460 2431
rect 40408 2388 40460 2397
rect 40592 2388 40644 2440
rect 41236 2388 41288 2440
rect 43812 2388 43864 2440
rect 38016 2320 38068 2372
rect 39304 2320 39356 2372
rect 40684 2320 40736 2372
rect 41420 2320 41472 2372
rect 41604 2320 41656 2372
rect 47032 2388 47084 2440
rect 48044 2388 48096 2440
rect 46388 2320 46440 2372
rect 40776 2252 40828 2304
rect 45468 2295 45520 2304
rect 45468 2261 45477 2295
rect 45477 2261 45511 2295
rect 45511 2261 45520 2295
rect 45468 2252 45520 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 35624 2048 35676 2100
rect 40684 2048 40736 2100
rect 23388 1980 23440 2032
rect 45468 1980 45520 2032
rect 26332 1912 26384 1964
rect 40316 1912 40368 1964
rect 15752 1844 15804 1896
rect 36176 1844 36228 1896
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 32 21622 60 49200
rect 1858 47696 1914 47705
rect 1858 47631 1914 47640
rect 1872 46646 1900 47631
rect 1964 47054 1992 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2608 46918 2636 49200
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3514 47016 3570 47025
rect 3514 46951 3570 46960
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 1860 46640 1912 46646
rect 1860 46582 1912 46588
rect 2320 46368 2372 46374
rect 2320 46310 2372 46316
rect 2780 46368 2832 46374
rect 2780 46310 2832 46316
rect 2962 46336 3018 46345
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1676 43240 1728 43246
rect 1676 43182 1728 43188
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 40225 1440 40462
rect 1398 40216 1454 40225
rect 1398 40151 1454 40160
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1412 35698 1440 36110
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1596 35086 1624 35391
rect 1584 35080 1636 35086
rect 1584 35022 1636 35028
rect 1492 34944 1544 34950
rect 1492 34886 1544 34892
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1504 33046 1532 34886
rect 1492 33040 1544 33046
rect 1492 32982 1544 32988
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1596 31822 1624 32671
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1688 26234 1716 43182
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 2136 41132 2188 41138
rect 2136 41074 2188 41080
rect 1768 40384 1820 40390
rect 1768 40326 1820 40332
rect 1780 29238 1808 40326
rect 1952 32224 2004 32230
rect 1952 32166 2004 32172
rect 1964 31346 1992 32166
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1768 29232 1820 29238
rect 1768 29174 1820 29180
rect 1596 26206 1716 26234
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23225 1440 23666
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 20 21616 72 21622
rect 20 21558 72 21564
rect 1596 19242 1624 26206
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 1964 20890 1992 25094
rect 1872 20862 1992 20890
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1584 19236 1636 19242
rect 1584 19178 1636 19184
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1872 8090 1900 20862
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2148 17678 2176 41074
rect 2228 36100 2280 36106
rect 2228 36042 2280 36048
rect 2240 35290 2268 36042
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 2228 35080 2280 35086
rect 2228 35022 2280 35028
rect 2240 19394 2268 35022
rect 2332 26042 2360 46310
rect 2792 45422 2820 46310
rect 2962 46271 3018 46280
rect 2872 45824 2924 45830
rect 2872 45766 2924 45772
rect 2884 45558 2912 45766
rect 2872 45552 2924 45558
rect 2872 45494 2924 45500
rect 2976 45422 3004 46271
rect 3056 45960 3108 45966
rect 3056 45902 3108 45908
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 2964 45416 3016 45422
rect 2964 45358 3016 45364
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36242 2820 36751
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 2688 33516 2740 33522
rect 2688 33458 2740 33464
rect 2700 32502 2728 33458
rect 2780 33312 2832 33318
rect 2780 33254 2832 33260
rect 2688 32496 2740 32502
rect 2688 32438 2740 32444
rect 2792 32026 2820 33254
rect 2962 32056 3018 32065
rect 2780 32020 2832 32026
rect 2962 31991 3018 32000
rect 2780 31962 2832 31968
rect 2872 31680 2924 31686
rect 2872 31622 2924 31628
rect 2884 31414 2912 31622
rect 2872 31408 2924 31414
rect 2872 31350 2924 31356
rect 2976 31278 3004 31991
rect 3068 31958 3096 45902
rect 3422 44976 3478 44985
rect 3422 44911 3478 44920
rect 3330 39536 3386 39545
rect 3330 39471 3386 39480
rect 3344 39098 3372 39471
rect 3332 39092 3384 39098
rect 3332 39034 3384 39040
rect 3240 32836 3292 32842
rect 3240 32778 3292 32784
rect 3252 32366 3280 32778
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 3056 31952 3108 31958
rect 3056 31894 3108 31900
rect 3068 31822 3096 31894
rect 3056 31816 3108 31822
rect 3056 31758 3108 31764
rect 2964 31272 3016 31278
rect 2964 31214 3016 31220
rect 2320 26036 2372 26042
rect 2320 25978 2372 25984
rect 2240 19366 2360 19394
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2332 18766 2360 19366
rect 3252 18970 3280 32302
rect 3330 28656 3386 28665
rect 3330 28591 3386 28600
rect 3344 27674 3372 28591
rect 3332 27668 3384 27674
rect 3332 27610 3384 27616
rect 3436 20058 3464 44911
rect 3528 22710 3556 46951
rect 3896 46594 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 47054 4752 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7328 49314
rect 7074 49200 7186 49286
rect 5828 47054 5856 49200
rect 7300 47054 7328 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49200 13626 50000
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 4712 47048 4764 47054
rect 4712 46990 4764 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7288 47048 7340 47054
rect 7288 46990 7340 46996
rect 8206 47016 8262 47025
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 4988 46980 5040 46986
rect 4988 46922 5040 46928
rect 6644 46980 6696 46986
rect 8206 46951 8208 46960
rect 6644 46922 6696 46928
rect 8260 46951 8262 46960
rect 8208 46922 8260 46928
rect 3896 46566 4016 46594
rect 3988 46510 4016 46566
rect 3884 46504 3936 46510
rect 3884 46446 3936 46452
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3896 46170 3924 46446
rect 3884 46164 3936 46170
rect 3884 46106 3936 46112
rect 3606 43616 3662 43625
rect 3606 43551 3662 43560
rect 3620 24614 3648 43551
rect 3976 33312 4028 33318
rect 3976 33254 4028 33260
rect 3988 32910 4016 33254
rect 3976 32904 4028 32910
rect 3976 32846 4028 32852
rect 3790 31376 3846 31385
rect 3790 31311 3846 31320
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3804 21350 3832 31311
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3988 19825 4016 20538
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2962 18456 3018 18465
rect 2962 18391 3018 18400
rect 2976 18222 3004 18391
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2884 17882 2912 18158
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17270 1992 17478
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2056 16794 2084 17070
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2792 16425 2820 17070
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2884 14414 2912 17614
rect 3516 17128 3568 17134
rect 3514 17096 3516 17105
rect 3568 17096 3570 17105
rect 3514 17031 3570 17040
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 2148 3534 2176 14350
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3344 6914 3372 12922
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10305 3464 10950
rect 3422 10296 3478 10305
rect 3422 10231 3478 10240
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7585 3464 8230
rect 3422 7576 3478 7585
rect 3422 7511 3478 7520
rect 3344 6886 3464 6914
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2976 3738 3004 4014
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1780 3058 1808 3470
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3126 1992 3334
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 1320 800 1348 2314
rect 2608 800 2636 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3068 785 3096 4014
rect 3252 2650 3280 6122
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3436 1465 3464 6886
rect 3528 3505 3556 12650
rect 3712 6905 3740 13942
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3988 13705 4016 13738
rect 3974 13696 4030 13705
rect 3974 13631 4030 13640
rect 4080 6914 4108 46922
rect 4620 46436 4672 46442
rect 4620 46378 4672 46384
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4632 46170 4660 46378
rect 4620 46164 4672 46170
rect 4620 46106 4672 46112
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 5000 19961 5028 46922
rect 4986 19952 5042 19961
rect 4986 19887 5042 19896
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3698 6896 3754 6905
rect 3698 6831 3754 6840
rect 3988 6886 4108 6914
rect 3988 5370 4016 6886
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 6656 5302 6684 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 46034 10456 46310
rect 10980 46034 11008 49200
rect 11624 47054 11652 49200
rect 12268 47054 12296 49200
rect 12912 47054 12940 49200
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 12256 47048 12308 47054
rect 12256 46990 12308 46996
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 11704 46980 11756 46986
rect 11704 46922 11756 46928
rect 12440 46980 12492 46986
rect 12440 46922 12492 46928
rect 13360 46980 13412 46986
rect 13360 46922 13412 46928
rect 10416 46028 10468 46034
rect 10416 45970 10468 45976
rect 10968 46028 11020 46034
rect 10968 45970 11020 45976
rect 10600 45892 10652 45898
rect 10600 45834 10652 45840
rect 10508 45824 10560 45830
rect 10508 45766 10560 45772
rect 8312 45526 8432 45554
rect 7564 39092 7616 39098
rect 7564 39034 7616 39040
rect 7576 27334 7604 39034
rect 8208 38888 8260 38894
rect 8208 38830 8260 38836
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 3988 3738 4016 3946
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5908 3528 5960 3534
rect 3514 3496 3570 3505
rect 5908 3470 5960 3476
rect 3514 3431 3570 3440
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 3896 800 3924 3130
rect 5920 3058 5948 3470
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5184 800 5212 2382
rect 6472 800 6500 3538
rect 7116 800 7144 3946
rect 7392 3058 7420 4014
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7576 2854 7604 4014
rect 8220 3534 8248 38830
rect 8312 32026 8340 45526
rect 10520 45490 10548 45766
rect 10612 45626 10640 45834
rect 10600 45620 10652 45626
rect 10600 45562 10652 45568
rect 10508 45484 10560 45490
rect 10508 45426 10560 45432
rect 11716 33114 11744 46922
rect 12452 36786 12480 46922
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 11704 32972 11756 32978
rect 11704 32914 11756 32920
rect 9680 32836 9732 32842
rect 9680 32778 9732 32784
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 9416 31890 9444 32234
rect 9404 31884 9456 31890
rect 9404 31826 9456 31832
rect 9692 31346 9720 32778
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 9876 31890 9904 31962
rect 9772 31884 9824 31890
rect 9772 31826 9824 31832
rect 9864 31884 9916 31890
rect 9864 31826 9916 31832
rect 9784 31482 9812 31826
rect 11532 31482 11560 32302
rect 11716 32026 11744 32914
rect 13268 32904 13320 32910
rect 13268 32846 13320 32852
rect 11796 32768 11848 32774
rect 11796 32710 11848 32716
rect 11808 32502 11836 32710
rect 11796 32496 11848 32502
rect 11796 32438 11848 32444
rect 12808 32496 12860 32502
rect 12808 32438 12860 32444
rect 12820 32026 12848 32438
rect 13280 32230 13308 32846
rect 13268 32224 13320 32230
rect 13268 32166 13320 32172
rect 11704 32020 11756 32026
rect 11704 31962 11756 31968
rect 12808 32020 12860 32026
rect 12808 31962 12860 31968
rect 12900 31884 12952 31890
rect 12900 31826 12952 31832
rect 12624 31816 12676 31822
rect 12624 31758 12676 31764
rect 12532 31748 12584 31754
rect 12532 31690 12584 31696
rect 9772 31476 9824 31482
rect 9772 31418 9824 31424
rect 11520 31476 11572 31482
rect 11520 31418 11572 31424
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 9128 29572 9180 29578
rect 9128 29514 9180 29520
rect 9036 29232 9088 29238
rect 9036 29174 9088 29180
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8944 24744 8996 24750
rect 8944 24686 8996 24692
rect 8588 24342 8616 24686
rect 8576 24336 8628 24342
rect 8576 24278 8628 24284
rect 8956 23866 8984 24686
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 8956 22030 8984 23666
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8864 21622 8892 21830
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 9048 17134 9076 29174
rect 9140 29170 9168 29514
rect 9128 29164 9180 29170
rect 9128 29106 9180 29112
rect 9692 28558 9720 31282
rect 10980 30734 11008 31282
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 11704 30728 11756 30734
rect 11704 30670 11756 30676
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9784 28762 9812 29038
rect 9772 28756 9824 28762
rect 9772 28698 9824 28704
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9692 26994 9720 28494
rect 10980 28150 11008 30670
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 11072 30258 11100 30602
rect 11060 30252 11112 30258
rect 11060 30194 11112 30200
rect 11716 29850 11744 30670
rect 12544 30598 12572 31690
rect 11796 30592 11848 30598
rect 11796 30534 11848 30540
rect 12532 30592 12584 30598
rect 12532 30534 12584 30540
rect 11808 30326 11836 30534
rect 11796 30320 11848 30326
rect 11796 30262 11848 30268
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 12452 29850 12480 30262
rect 11704 29844 11756 29850
rect 11704 29786 11756 29792
rect 12440 29844 12492 29850
rect 12440 29786 12492 29792
rect 12544 29730 12572 30534
rect 12452 29702 12572 29730
rect 11244 29640 11296 29646
rect 11244 29582 11296 29588
rect 11256 28694 11284 29582
rect 12452 29510 12480 29702
rect 12636 29646 12664 31758
rect 12912 30870 12940 31826
rect 12900 30864 12952 30870
rect 12900 30806 12952 30812
rect 12716 30660 12768 30666
rect 12716 30602 12768 30608
rect 12728 29714 12756 30602
rect 12912 30598 12940 30806
rect 13268 30796 13320 30802
rect 13268 30738 13320 30744
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 13096 30598 13124 30670
rect 13280 30598 13308 30738
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 13268 30592 13320 30598
rect 13268 30534 13320 30540
rect 12716 29708 12768 29714
rect 12716 29650 12768 29656
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12440 29504 12492 29510
rect 12440 29446 12492 29452
rect 11244 28688 11296 28694
rect 11244 28630 11296 28636
rect 10968 28144 11020 28150
rect 10968 28086 11020 28092
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9784 27130 9812 27338
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 10980 26994 11008 28086
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 9692 25770 9720 26930
rect 10796 25838 10824 26930
rect 11060 26852 11112 26858
rect 11060 26794 11112 26800
rect 11072 26586 11100 26794
rect 11060 26580 11112 26586
rect 11060 26522 11112 26528
rect 11256 26382 11284 28630
rect 11796 28620 11848 28626
rect 11796 28562 11848 28568
rect 11808 28150 11836 28562
rect 12452 28558 12480 29446
rect 12636 28966 12664 29582
rect 12912 29238 12940 30534
rect 13096 30190 13124 30534
rect 13280 30394 13308 30534
rect 13268 30388 13320 30394
rect 13268 30330 13320 30336
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13280 29578 13308 30330
rect 13268 29572 13320 29578
rect 13268 29514 13320 29520
rect 12900 29232 12952 29238
rect 12900 29174 12952 29180
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 13372 28762 13400 46922
rect 13556 46918 13584 49200
rect 13544 46912 13596 46918
rect 13544 46854 13596 46860
rect 14200 46510 14228 49200
rect 14648 46980 14700 46986
rect 14648 46922 14700 46928
rect 13728 46504 13780 46510
rect 13728 46446 13780 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 13740 45626 13768 46446
rect 13728 45620 13780 45626
rect 13728 45562 13780 45568
rect 14660 35894 14688 46922
rect 15488 45554 15516 49200
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49200 27150 50000
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49200 31014 50000
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49200 41318 50000
rect 41850 49314 41962 50000
rect 41850 49286 42288 49314
rect 41850 49200 41962 49286
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 16948 47048 17000 47054
rect 16948 46990 17000 46996
rect 16120 45620 16172 45626
rect 16120 45562 16172 45568
rect 15488 45526 16068 45554
rect 14568 35866 14688 35894
rect 13636 33448 13688 33454
rect 13636 33390 13688 33396
rect 14372 33448 14424 33454
rect 14372 33390 14424 33396
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13556 32434 13584 32846
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 13648 31754 13676 33390
rect 14384 32570 14412 33390
rect 14372 32564 14424 32570
rect 14372 32506 14424 32512
rect 14096 32360 14148 32366
rect 14096 32302 14148 32308
rect 13728 32224 13780 32230
rect 13728 32166 13780 32172
rect 13556 31726 13676 31754
rect 13556 30666 13584 31726
rect 13740 30734 13768 32166
rect 14108 31482 14136 32302
rect 14096 31476 14148 31482
rect 14096 31418 14148 31424
rect 13912 31272 13964 31278
rect 13912 31214 13964 31220
rect 13728 30728 13780 30734
rect 13728 30670 13780 30676
rect 13544 30660 13596 30666
rect 13544 30602 13596 30608
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 13372 28490 13400 28698
rect 13360 28484 13412 28490
rect 13360 28426 13412 28432
rect 13464 28422 13492 29106
rect 13556 28558 13584 30602
rect 13924 30394 13952 31214
rect 14108 30870 14136 31418
rect 14096 30864 14148 30870
rect 14096 30806 14148 30812
rect 13912 30388 13964 30394
rect 13912 30330 13964 30336
rect 14108 30122 14136 30806
rect 14096 30116 14148 30122
rect 14096 30058 14148 30064
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13910 28520 13966 28529
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 11796 28144 11848 28150
rect 11796 28086 11848 28092
rect 12440 28144 12492 28150
rect 12440 28086 12492 28092
rect 12452 27606 12480 28086
rect 12440 27600 12492 27606
rect 12440 27542 12492 27548
rect 11520 27532 11572 27538
rect 11520 27474 11572 27480
rect 11060 26376 11112 26382
rect 11060 26318 11112 26324
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 10784 25832 10836 25838
rect 10784 25774 10836 25780
rect 11072 25770 11100 26318
rect 11532 25974 11560 27474
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11900 26586 11928 26998
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 12544 26382 12572 27406
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 11520 25968 11572 25974
rect 11520 25910 11572 25916
rect 11428 25900 11480 25906
rect 11428 25842 11480 25848
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 9680 25764 9732 25770
rect 9680 25706 9732 25712
rect 11060 25764 11112 25770
rect 11060 25706 11112 25712
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9876 25362 9904 25638
rect 11440 25498 11468 25842
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 10152 24410 10180 25162
rect 11440 24682 11468 25434
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11532 24886 11560 25094
rect 11520 24880 11572 24886
rect 11520 24822 11572 24828
rect 11428 24676 11480 24682
rect 11428 24618 11480 24624
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 11440 24206 11468 24618
rect 11532 24342 11560 24822
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 11716 24206 11744 24550
rect 11992 24410 12020 24754
rect 12084 24614 12112 25842
rect 12544 25294 12572 26318
rect 13096 25974 13124 26726
rect 13464 26382 13492 28358
rect 13556 28150 13584 28494
rect 13910 28455 13912 28464
rect 13964 28455 13966 28464
rect 13912 28426 13964 28432
rect 13544 28144 13596 28150
rect 13544 28086 13596 28092
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13832 26858 13860 27406
rect 13820 26852 13872 26858
rect 13820 26794 13872 26800
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13084 25968 13136 25974
rect 13084 25910 13136 25916
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11164 23866 11192 24006
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9968 22166 9996 22578
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9140 21010 9168 21830
rect 9968 21078 9996 22102
rect 10244 22098 10272 22918
rect 11164 22574 11192 23802
rect 11532 23798 11560 24142
rect 11992 24070 12020 24346
rect 12084 24206 12112 24550
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11520 23792 11572 23798
rect 11520 23734 11572 23740
rect 11808 23594 11836 24006
rect 11796 23588 11848 23594
rect 11796 23530 11848 23536
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11716 23186 11744 23462
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11348 22642 11376 22986
rect 11440 22778 11468 23054
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10336 22234 10364 22374
rect 10324 22228 10376 22234
rect 10324 22170 10376 22176
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 11072 21962 11100 22374
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 10796 11014 10824 20810
rect 10980 20534 11008 21626
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 11164 20466 11192 22510
rect 11992 22098 12020 24006
rect 12084 23866 12112 24142
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 12452 22778 12480 22986
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12544 22658 12572 25230
rect 13188 25158 13216 25842
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13280 25498 13308 25638
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12728 24070 12756 24754
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 13188 22982 13216 24074
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 12452 22642 12572 22658
rect 13188 22642 13216 22918
rect 12440 22636 12572 22642
rect 12492 22630 12572 22636
rect 13176 22636 13228 22642
rect 12440 22578 12492 22584
rect 13176 22578 13228 22584
rect 12452 22506 12480 22578
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 12820 22166 12848 22510
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12544 21622 12572 21966
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12820 20466 12848 22102
rect 13740 21622 13768 25094
rect 13832 24206 13860 26794
rect 13924 24682 13952 28426
rect 14292 28422 14320 29038
rect 14476 28422 14504 29106
rect 14568 28626 14596 35866
rect 16040 33590 16068 45526
rect 16028 33584 16080 33590
rect 16028 33526 16080 33532
rect 16132 32978 16160 45562
rect 16960 34066 16988 46990
rect 17420 45626 17448 49200
rect 18708 47054 18736 49200
rect 19996 47054 20024 49200
rect 18696 47048 18748 47054
rect 18696 46990 18748 46996
rect 19984 47048 20036 47054
rect 19984 46990 20036 46996
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 18880 46980 18932 46986
rect 18880 46922 18932 46928
rect 17408 45620 17460 45626
rect 17408 45562 17460 45568
rect 16948 34060 17000 34066
rect 16948 34002 17000 34008
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14660 30326 14688 31078
rect 15212 30938 15240 31826
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 15384 31680 15436 31686
rect 15384 31622 15436 31628
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 14740 30592 14792 30598
rect 14740 30534 14792 30540
rect 14648 30320 14700 30326
rect 14648 30262 14700 30268
rect 14648 28960 14700 28966
rect 14648 28902 14700 28908
rect 14660 28694 14688 28902
rect 14648 28688 14700 28694
rect 14648 28630 14700 28636
rect 14556 28620 14608 28626
rect 14556 28562 14608 28568
rect 14280 28416 14332 28422
rect 14464 28416 14516 28422
rect 14332 28376 14412 28404
rect 14280 28358 14332 28364
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14108 27062 14136 27406
rect 14384 27334 14412 28376
rect 14464 28358 14516 28364
rect 14660 28370 14688 28630
rect 14752 28490 14780 30534
rect 15212 30190 15240 30874
rect 15396 30802 15424 31622
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15384 30796 15436 30802
rect 15384 30738 15436 30744
rect 15200 30184 15252 30190
rect 15200 30126 15252 30132
rect 15580 29646 15608 31282
rect 15752 30728 15804 30734
rect 15752 30670 15804 30676
rect 16592 30682 16620 31758
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 15764 30394 15792 30670
rect 16592 30654 16712 30682
rect 16776 30666 16804 31078
rect 16684 30598 16712 30654
rect 16764 30660 16816 30666
rect 16764 30602 16816 30608
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 17500 30592 17552 30598
rect 17500 30534 17552 30540
rect 15752 30388 15804 30394
rect 15752 30330 15804 30336
rect 16120 30252 16172 30258
rect 16120 30194 16172 30200
rect 16132 29714 16160 30194
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 15568 29640 15620 29646
rect 15620 29600 15792 29628
rect 15568 29582 15620 29588
rect 15764 29170 15792 29600
rect 15936 29572 15988 29578
rect 15936 29514 15988 29520
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15200 29096 15252 29102
rect 15200 29038 15252 29044
rect 15212 28558 15240 29038
rect 15200 28552 15252 28558
rect 15384 28552 15436 28558
rect 15200 28494 15252 28500
rect 15382 28520 15384 28529
rect 15436 28520 15438 28529
rect 14740 28484 14792 28490
rect 14740 28426 14792 28432
rect 15016 28484 15068 28490
rect 15382 28455 15438 28464
rect 15016 28426 15068 28432
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14476 27130 14504 28358
rect 14660 28342 14780 28370
rect 14752 28082 14780 28342
rect 15028 28082 15056 28426
rect 15292 28416 15344 28422
rect 15488 28404 15516 29106
rect 15948 29102 15976 29514
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15936 29096 15988 29102
rect 15936 29038 15988 29044
rect 15344 28376 15516 28404
rect 15292 28358 15344 28364
rect 15488 28082 15516 28376
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15580 28218 15608 28358
rect 15568 28212 15620 28218
rect 15568 28154 15620 28160
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 15476 28076 15528 28082
rect 15476 28018 15528 28024
rect 14752 27130 14780 28018
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14096 27056 14148 27062
rect 14096 26998 14148 27004
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 14568 26246 14596 26930
rect 14832 26920 14884 26926
rect 14832 26862 14884 26868
rect 14844 26314 14872 26862
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 14924 26376 14976 26382
rect 14976 26336 15056 26364
rect 14924 26318 14976 26324
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14384 25498 14412 25774
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 13912 24676 13964 24682
rect 13912 24618 13964 24624
rect 14200 24410 14228 24686
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 13912 24132 13964 24138
rect 13912 24074 13964 24080
rect 13924 23730 13952 24074
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14108 23798 14136 24006
rect 14096 23792 14148 23798
rect 14096 23734 14148 23740
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 13912 22976 13964 22982
rect 13912 22918 13964 22924
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13832 22098 13860 22510
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 13924 22030 13952 22918
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13924 21554 13952 21966
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11440 19922 11468 20198
rect 12728 19990 12756 20402
rect 12716 19984 12768 19990
rect 12716 19926 12768 19932
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 12820 19718 12848 20402
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12820 19378 12848 19654
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 13004 19174 13032 20334
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13924 18766 13952 19450
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14016 18834 14044 19314
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13372 18086 13400 18702
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9508 3602 9536 4558
rect 13740 4146 13768 18566
rect 14108 17882 14136 20742
rect 14200 20602 14228 23598
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14292 19854 14320 21966
rect 14384 19990 14412 25434
rect 14568 25226 14596 26182
rect 14844 26042 14872 26250
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14660 25226 14688 25842
rect 15028 25770 15056 26336
rect 15200 26036 15252 26042
rect 15200 25978 15252 25984
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15016 25764 15068 25770
rect 15016 25706 15068 25712
rect 15028 25242 15056 25706
rect 15120 25362 15148 25842
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 14556 25220 14608 25226
rect 14556 25162 14608 25168
rect 14648 25220 14700 25226
rect 15028 25214 15148 25242
rect 14648 25162 14700 25168
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14476 24886 14504 25094
rect 14464 24880 14516 24886
rect 14464 24822 14516 24828
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14200 19378 14228 19722
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14292 19242 14320 19790
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14384 19446 14412 19654
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 18358 14320 18566
rect 14476 18442 14504 24686
rect 14568 20806 14596 25162
rect 14660 23118 14688 25162
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14660 21690 14688 21898
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14844 19922 14872 20878
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14936 20466 14964 20742
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 15028 20074 15056 23054
rect 15120 20874 15148 25214
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15120 20466 15148 20810
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 14936 20046 15056 20074
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14384 18414 14504 18442
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16658 14136 16934
rect 14096 16652 14148 16658
rect 14384 16640 14412 18414
rect 14568 18290 14596 19314
rect 14660 19174 14688 19654
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14096 16594 14148 16600
rect 14292 16612 14412 16640
rect 14476 18170 14504 18226
rect 14660 18170 14688 19110
rect 14752 18630 14780 19382
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14844 18222 14872 19858
rect 14936 18834 14964 20046
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 15028 19514 15056 19858
rect 15120 19854 15148 20198
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15120 18358 15148 18634
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 14924 18284 14976 18290
rect 14976 18244 15056 18272
rect 14924 18226 14976 18232
rect 14476 18142 14688 18170
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14292 13802 14320 16612
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14384 16046 14412 16458
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14476 15978 14504 18142
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14844 17678 14872 17818
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14568 16794 14596 17138
rect 14844 17134 14872 17614
rect 15028 17542 15056 18244
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14568 15026 14596 16730
rect 15028 16182 15056 17478
rect 15120 17202 15148 18158
rect 15212 17610 15240 25978
rect 15304 25294 15332 26726
rect 15396 26586 15424 26930
rect 15384 26580 15436 26586
rect 15384 26522 15436 26528
rect 15488 26042 15516 27270
rect 15580 27130 15608 28154
rect 15672 28082 15700 29038
rect 16132 28558 16160 29650
rect 17040 29572 17092 29578
rect 17040 29514 17092 29520
rect 17052 29306 17080 29514
rect 17040 29300 17092 29306
rect 17040 29242 17092 29248
rect 16120 28552 16172 28558
rect 17512 28529 17540 30534
rect 18052 29504 18104 29510
rect 18052 29446 18104 29452
rect 18064 29238 18092 29446
rect 18052 29232 18104 29238
rect 18052 29174 18104 29180
rect 16120 28494 16172 28500
rect 17498 28520 17554 28529
rect 15660 28076 15712 28082
rect 15660 28018 15712 28024
rect 15568 27124 15620 27130
rect 15568 27066 15620 27072
rect 15580 26314 15608 27066
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15568 26308 15620 26314
rect 15568 26250 15620 26256
rect 15672 26042 15700 26318
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 15476 26036 15528 26042
rect 15476 25978 15528 25984
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15580 25498 15608 25842
rect 15948 25498 15976 26250
rect 16132 25906 16160 28494
rect 17498 28455 17554 28464
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16684 28082 16712 28358
rect 17960 28144 18012 28150
rect 17960 28086 18012 28092
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17420 26042 17448 26930
rect 17604 26858 17632 27406
rect 17972 27130 18000 28086
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 17960 26988 18012 26994
rect 18064 26976 18092 29174
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 18328 29096 18380 29102
rect 18328 29038 18380 29044
rect 18156 28234 18184 29038
rect 18156 28218 18276 28234
rect 18156 28212 18288 28218
rect 18156 28206 18236 28212
rect 18156 28014 18184 28206
rect 18236 28154 18288 28160
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18340 27606 18368 29038
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 18012 26948 18092 26976
rect 17960 26930 18012 26936
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17604 26382 17632 26794
rect 18156 26586 18184 26862
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17408 26036 17460 26042
rect 17408 25978 17460 25984
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 17420 25702 17448 25978
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15936 25492 15988 25498
rect 15936 25434 15988 25440
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15856 24818 15884 25230
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15856 24342 15884 24754
rect 16120 24676 16172 24682
rect 16120 24618 16172 24624
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15660 24268 15712 24274
rect 15660 24210 15712 24216
rect 15384 24064 15436 24070
rect 15384 24006 15436 24012
rect 15396 23186 15424 24006
rect 15672 23186 15700 24210
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15212 17270 15240 17546
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 15120 16114 15148 17138
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15396 16522 15424 16934
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15212 15994 15240 16390
rect 15120 15978 15240 15994
rect 15108 15972 15240 15978
rect 15160 15966 15240 15972
rect 15108 15914 15160 15920
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14752 15162 14780 15438
rect 14936 15434 14964 15846
rect 15028 15570 15056 15846
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 15120 13938 15148 15914
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8220 3126 8248 3334
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7760 800 7788 2858
rect 8036 2650 8064 2926
rect 9600 2854 9628 3538
rect 10244 3466 10272 3878
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 11532 3058 11560 3878
rect 12084 3534 12112 3946
rect 13740 3670 13768 4082
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 3126 11744 3334
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 13832 3058 13860 3470
rect 14016 3126 14044 3878
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8404 800 8432 2382
rect 9048 800 9076 2790
rect 10980 800 11008 2926
rect 14200 800 14228 2926
rect 14844 800 14872 12582
rect 15580 6254 15608 22510
rect 16132 22098 16160 24618
rect 17420 24290 17448 25638
rect 17604 25498 17632 26318
rect 18788 26308 18840 26314
rect 18788 26250 18840 26256
rect 18800 26042 18828 26250
rect 18788 26036 18840 26042
rect 18788 25978 18840 25984
rect 18144 25696 18196 25702
rect 18144 25638 18196 25644
rect 17592 25492 17644 25498
rect 17592 25434 17644 25440
rect 18156 25294 18184 25638
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17420 24274 17632 24290
rect 17420 24268 17644 24274
rect 17420 24262 17592 24268
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16684 23186 16712 24142
rect 16856 24132 16908 24138
rect 16856 24074 16908 24080
rect 16868 23526 16896 24074
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16592 21146 16620 21966
rect 16684 21690 16712 23122
rect 16776 23118 16804 23462
rect 16868 23254 16896 23462
rect 16960 23322 16988 24142
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17236 23866 17264 24074
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17420 23730 17448 24262
rect 17592 24210 17644 24216
rect 17788 23730 17816 24550
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16856 23248 16908 23254
rect 16856 23190 16908 23196
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 17420 22642 17448 23666
rect 18340 23526 18368 24754
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18524 24070 18552 24686
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18512 24064 18564 24070
rect 18432 24024 18512 24052
rect 18432 23798 18460 24024
rect 18512 24006 18564 24012
rect 18420 23792 18472 23798
rect 18420 23734 18472 23740
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 18340 22506 18368 23462
rect 18432 22778 18460 23734
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18328 22500 18380 22506
rect 18328 22442 18380 22448
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 22030 18000 22374
rect 18052 22228 18104 22234
rect 18052 22170 18104 22176
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16684 20942 16712 21626
rect 18064 21486 18092 22170
rect 18432 22098 18460 22578
rect 18708 22574 18736 24210
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18800 23526 18828 23666
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18340 21554 18368 21966
rect 18432 21894 18460 22034
rect 18708 21962 18736 22510
rect 18800 22030 18828 23462
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18420 21888 18472 21894
rect 18420 21830 18472 21836
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18432 21622 18460 21830
rect 18420 21616 18472 21622
rect 18420 21558 18472 21564
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15672 19990 15700 20334
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 16684 19854 16712 20878
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17972 20466 18000 20742
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18248 19854 18276 20198
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17236 19378 17264 19654
rect 18248 19446 18276 19654
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 16040 18222 16068 18634
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15856 12918 15884 13466
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 16040 4078 16068 18158
rect 16408 17678 16436 18566
rect 16776 18290 16804 18702
rect 18432 18290 18460 21558
rect 18524 21554 18552 21830
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18524 20534 18552 21286
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18524 18902 18552 19246
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16684 17202 16712 18022
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 16776 17338 16804 17546
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16684 16266 16712 17138
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17696 16658 17724 17002
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 16684 16238 16804 16266
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 15366 16712 16050
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 12850 16712 15302
rect 16776 13190 16804 16238
rect 17420 15162 17448 16594
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 15162 17632 15982
rect 17880 15910 17908 16526
rect 17972 16182 18000 16594
rect 18248 16522 18276 17546
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18432 16250 18460 16526
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17420 14550 17448 15098
rect 17788 15094 17816 15642
rect 17880 15434 17908 15846
rect 18432 15502 18460 16186
rect 18616 16046 18644 16390
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17788 14414 17816 15030
rect 17880 14890 17908 15370
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18064 15026 18092 15302
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16580 12776 16632 12782
rect 16776 12730 16804 13126
rect 16632 12724 16804 12730
rect 16580 12718 16804 12724
rect 16592 12702 16804 12718
rect 16776 12238 16804 12702
rect 16868 12442 16896 13806
rect 17788 13462 17816 14350
rect 17880 14346 17908 14826
rect 18340 14618 18368 14894
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16960 12646 16988 13330
rect 17880 13326 17908 14282
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 17972 12442 18000 13330
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 18064 8294 18092 12718
rect 18524 8294 18552 13806
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2446 15240 2926
rect 16868 2650 16896 7686
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17052 3738 17080 4082
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17236 2990 17264 3470
rect 17512 3058 17540 4082
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17696 3058 17724 3334
rect 17788 3126 17816 4082
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 800 15516 2314
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 1902 15792 2246
rect 15752 1896 15804 1902
rect 15752 1838 15804 1844
rect 16132 800 16160 2382
rect 17420 800 17448 2926
rect 17972 2446 18000 3878
rect 18064 2650 18092 4558
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18156 2446 18184 4422
rect 18708 4078 18736 5170
rect 18892 4758 18920 46922
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19432 46504 19484 46510
rect 19432 46446 19484 46452
rect 20168 46504 20220 46510
rect 20168 46446 20220 46452
rect 19444 46170 19472 46446
rect 20180 46170 20208 46446
rect 19432 46164 19484 46170
rect 19432 46106 19484 46112
rect 20168 46164 20220 46170
rect 20168 46106 20220 46112
rect 20076 45960 20128 45966
rect 20076 45902 20128 45908
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 20088 44402 20116 45902
rect 20076 44396 20128 44402
rect 20076 44338 20128 44344
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 20088 41138 20116 44338
rect 20076 41132 20128 41138
rect 20076 41074 20128 41080
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 20364 32910 20392 46990
rect 20640 46510 20668 49200
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20720 46368 20772 46374
rect 20720 46310 20772 46316
rect 20732 46034 20760 46310
rect 21284 46034 21312 49200
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 24872 46646 24900 46990
rect 24860 46640 24912 46646
rect 24860 46582 24912 46588
rect 25148 46510 25176 49200
rect 25504 47048 25556 47054
rect 25504 46990 25556 46996
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25516 46034 25544 46990
rect 25792 46034 25820 49200
rect 27080 46646 27108 49200
rect 28368 47054 28396 49200
rect 29656 47054 29684 49200
rect 30944 47138 30972 49200
rect 30944 47110 31064 47138
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 30932 47048 30984 47054
rect 30932 46990 30984 46996
rect 30196 46980 30248 46986
rect 30196 46922 30248 46928
rect 29920 46912 29972 46918
rect 29920 46854 29972 46860
rect 27068 46640 27120 46646
rect 27068 46582 27120 46588
rect 20720 46028 20772 46034
rect 20720 45970 20772 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 25504 46028 25556 46034
rect 25504 45970 25556 45976
rect 25780 46028 25832 46034
rect 25780 45970 25832 45976
rect 24860 45960 24912 45966
rect 24860 45902 24912 45908
rect 20904 45892 20956 45898
rect 20904 45834 20956 45840
rect 20916 45626 20944 45834
rect 20904 45620 20956 45626
rect 20904 45562 20956 45568
rect 24872 45558 24900 45902
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25424 45626 25452 45834
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 24860 45552 24912 45558
rect 24860 45494 24912 45500
rect 26056 45484 26108 45490
rect 26056 45426 26108 45432
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 25964 38956 26016 38962
rect 25964 38898 26016 38904
rect 23480 36032 23532 36038
rect 23480 35974 23532 35980
rect 22836 35760 22888 35766
rect 22836 35702 22888 35708
rect 22848 35290 22876 35702
rect 23492 35630 23520 35974
rect 23480 35624 23532 35630
rect 23480 35566 23532 35572
rect 24676 35624 24728 35630
rect 24676 35566 24728 35572
rect 24952 35624 25004 35630
rect 24952 35566 25004 35572
rect 24688 35494 24716 35566
rect 23480 35488 23532 35494
rect 23480 35430 23532 35436
rect 24676 35488 24728 35494
rect 24676 35430 24728 35436
rect 22836 35284 22888 35290
rect 22836 35226 22888 35232
rect 22008 35080 22060 35086
rect 22008 35022 22060 35028
rect 20812 34400 20864 34406
rect 20812 34342 20864 34348
rect 20824 34134 20852 34342
rect 22020 34134 22048 35022
rect 23492 34746 23520 35430
rect 24688 35222 24716 35430
rect 24964 35290 24992 35566
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 24676 35216 24728 35222
rect 24676 35158 24728 35164
rect 24492 35080 24544 35086
rect 24492 35022 24544 35028
rect 23480 34740 23532 34746
rect 23480 34682 23532 34688
rect 23204 34604 23256 34610
rect 23204 34546 23256 34552
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22836 34400 22888 34406
rect 22836 34342 22888 34348
rect 22664 34202 22692 34342
rect 22652 34196 22704 34202
rect 22652 34138 22704 34144
rect 20812 34128 20864 34134
rect 20812 34070 20864 34076
rect 22008 34128 22060 34134
rect 22008 34070 22060 34076
rect 20824 33998 20852 34070
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 20352 32904 20404 32910
rect 20352 32846 20404 32852
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 20824 31890 20852 33934
rect 20904 33856 20956 33862
rect 20904 33798 20956 33804
rect 20916 33522 20944 33798
rect 20904 33516 20956 33522
rect 20904 33458 20956 33464
rect 21928 33318 21956 33934
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22008 33448 22060 33454
rect 22008 33390 22060 33396
rect 21732 33312 21784 33318
rect 21732 33254 21784 33260
rect 21916 33312 21968 33318
rect 21916 33254 21968 33260
rect 21744 32434 21772 33254
rect 22020 33114 22048 33390
rect 22008 33108 22060 33114
rect 22008 33050 22060 33056
rect 22008 32836 22060 32842
rect 22008 32778 22060 32784
rect 22020 32434 22048 32778
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 21732 32428 21784 32434
rect 21732 32370 21784 32376
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 20812 31884 20864 31890
rect 20812 31826 20864 31832
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 20456 31414 20484 31758
rect 20812 31680 20864 31686
rect 20812 31622 20864 31628
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 19156 31272 19208 31278
rect 19156 31214 19208 31220
rect 20720 31272 20772 31278
rect 20720 31214 20772 31220
rect 19168 30802 19196 31214
rect 20732 30938 20760 31214
rect 20720 30932 20772 30938
rect 20720 30874 20772 30880
rect 19156 30796 19208 30802
rect 19156 30738 19208 30744
rect 20824 30666 20852 31622
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20812 30660 20864 30666
rect 20812 30602 20864 30608
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 20916 30258 20944 31078
rect 21744 30666 21772 32370
rect 22008 32292 22060 32298
rect 22008 32234 22060 32240
rect 22020 32201 22048 32234
rect 22006 32192 22062 32201
rect 22006 32127 22062 32136
rect 22204 31686 22232 32710
rect 21916 31680 21968 31686
rect 21916 31622 21968 31628
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 21824 31408 21876 31414
rect 21824 31350 21876 31356
rect 21836 31142 21864 31350
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21836 30734 21864 31078
rect 21928 30734 21956 31622
rect 22020 31278 22048 31622
rect 22008 31272 22060 31278
rect 22008 31214 22060 31220
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 21088 30660 21140 30666
rect 21088 30602 21140 30608
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 21008 30190 21036 30534
rect 21100 30326 21128 30602
rect 21456 30592 21508 30598
rect 21456 30534 21508 30540
rect 21088 30320 21140 30326
rect 21088 30262 21140 30268
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 21272 30048 21324 30054
rect 21272 29990 21324 29996
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 21284 29170 21312 29990
rect 21468 29850 21496 30534
rect 21744 30122 21772 30602
rect 21732 30116 21784 30122
rect 21732 30058 21784 30064
rect 21456 29844 21508 29850
rect 21456 29786 21508 29792
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21272 29164 21324 29170
rect 21272 29106 21324 29112
rect 21086 28656 21142 28665
rect 21086 28591 21142 28600
rect 21100 28558 21128 28591
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 21088 28552 21140 28558
rect 21088 28494 21140 28500
rect 19248 27600 19300 27606
rect 19248 27542 19300 27548
rect 19260 25362 19288 27542
rect 19352 26450 19380 28494
rect 20628 28484 20680 28490
rect 20628 28426 20680 28432
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 20640 28218 20668 28426
rect 20996 28416 21048 28422
rect 20996 28358 21048 28364
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 21008 28014 21036 28358
rect 20996 28008 21048 28014
rect 20996 27950 21048 27956
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19340 24812 19392 24818
rect 19444 24800 19472 26726
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 20088 25294 20116 26386
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19392 24772 19472 24800
rect 19340 24754 19392 24760
rect 19352 23866 19380 24754
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19996 23866 20024 24686
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 19352 23118 19380 23802
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19260 22778 19288 23054
rect 20168 22976 20220 22982
rect 20168 22918 20220 22924
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 19168 20312 19196 20878
rect 19260 20602 19288 21898
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 20180 21554 20208 22918
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19352 20466 19380 20742
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 20180 20398 20208 21490
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 19248 20324 19300 20330
rect 19168 20284 19248 20312
rect 19168 19854 19196 20284
rect 19248 20266 19300 20272
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 20180 19514 20208 20334
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20180 19378 20208 19450
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18984 18766 19012 19246
rect 20180 18834 20208 19314
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19352 16182 19380 16390
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19444 15178 19472 16526
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15570 19656 15846
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19352 15150 19472 15178
rect 19352 14958 19380 15150
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19352 14414 19380 14894
rect 19444 14618 19472 14962
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 18880 4752 18932 4758
rect 18880 4694 18932 4700
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18420 3664 18472 3670
rect 18418 3632 18420 3641
rect 18472 3632 18474 3641
rect 18418 3567 18474 3576
rect 18524 3534 18552 3878
rect 18616 3534 18644 3946
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18248 2650 18276 3402
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18708 800 18736 3606
rect 18800 3058 18828 3946
rect 18880 3460 18932 3466
rect 18880 3402 18932 3408
rect 18892 3126 18920 3402
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19260 2446 19288 4966
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19352 4282 19380 4558
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19352 2650 19380 4082
rect 19720 3738 19748 4082
rect 20272 3738 20300 26862
rect 20640 25906 20668 27814
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20824 26874 20852 27338
rect 21100 26994 21128 28494
rect 21180 28484 21232 28490
rect 21180 28426 21232 28432
rect 21192 28218 21220 28426
rect 21272 28416 21324 28422
rect 21272 28358 21324 28364
rect 21180 28212 21232 28218
rect 21180 28154 21232 28160
rect 21192 27062 21220 28154
rect 21284 28082 21312 28358
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21284 27946 21312 28018
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21284 27470 21312 27882
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21454 27296 21510 27305
rect 21454 27231 21510 27240
rect 21180 27056 21232 27062
rect 21180 26998 21232 27004
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21468 26926 21496 27231
rect 21456 26920 21508 26926
rect 20824 26858 21128 26874
rect 21456 26862 21508 26868
rect 20824 26852 21140 26858
rect 20824 26846 21088 26852
rect 21088 26794 21140 26800
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 20732 26518 20760 26726
rect 21008 26586 21036 26726
rect 21100 26586 21128 26794
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 20720 26512 20772 26518
rect 20720 26454 20772 26460
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20732 26042 20760 26250
rect 21468 26246 21496 26522
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 21270 24848 21326 24857
rect 21270 24783 21272 24792
rect 21324 24783 21326 24792
rect 21272 24754 21324 24760
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 23866 20668 24074
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18766 20576 19110
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20640 18578 20668 22918
rect 20732 22642 20760 23666
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20732 21434 20760 22578
rect 20916 22098 20944 23122
rect 20904 22092 20956 22098
rect 20904 22034 20956 22040
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 20732 21406 21220 21434
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21008 20942 21036 21286
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21008 20466 21036 20878
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20824 19174 20852 19246
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20916 18986 20944 19246
rect 20824 18958 20944 18986
rect 20824 18578 20852 18958
rect 20904 18896 20956 18902
rect 20904 18838 20956 18844
rect 20640 18550 20852 18578
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 16250 20392 16934
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20364 4146 20392 4422
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20456 3618 20484 18158
rect 20640 12434 20668 18550
rect 20916 18290 20944 18838
rect 21008 18290 21036 20402
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19922 21128 20198
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 21100 19514 21128 19722
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21100 18834 21128 19450
rect 21192 18902 21220 21406
rect 21468 19922 21496 21966
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21192 18358 21220 18702
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21192 17610 21220 18158
rect 21468 17882 21496 19858
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21192 17202 21220 17546
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 21100 16794 21128 17002
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21100 16114 21128 16730
rect 21468 16590 21496 17818
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20916 15570 20944 15846
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 21008 14890 21036 16050
rect 21376 15638 21404 16118
rect 21364 15632 21416 15638
rect 21364 15574 21416 15580
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21192 15162 21220 15370
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21376 15094 21404 15574
rect 21468 15366 21496 16526
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21364 15088 21416 15094
rect 21364 15030 21416 15036
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 21560 12434 21588 29446
rect 22020 29322 22048 31214
rect 22296 30258 22324 33798
rect 22376 33380 22428 33386
rect 22376 33322 22428 33328
rect 22388 32910 22416 33322
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22468 32904 22520 32910
rect 22468 32846 22520 32852
rect 22652 32904 22704 32910
rect 22652 32846 22704 32852
rect 22480 32570 22508 32846
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22664 32502 22692 32846
rect 22652 32496 22704 32502
rect 22652 32438 22704 32444
rect 22376 32428 22428 32434
rect 22376 32370 22428 32376
rect 22388 31822 22416 32370
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22388 31278 22416 31758
rect 22376 31272 22428 31278
rect 22376 31214 22428 31220
rect 22480 31142 22508 32302
rect 22652 32292 22704 32298
rect 22652 32234 22704 32240
rect 22664 31822 22692 32234
rect 22652 31816 22704 31822
rect 22652 31758 22704 31764
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22468 31136 22520 31142
rect 22468 31078 22520 31084
rect 22480 30938 22508 31078
rect 22468 30932 22520 30938
rect 22468 30874 22520 30880
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 22112 29782 22140 30194
rect 22100 29776 22152 29782
rect 22100 29718 22152 29724
rect 22192 29640 22244 29646
rect 21928 29294 22048 29322
rect 22112 29600 22192 29628
rect 21640 29164 21692 29170
rect 21640 29106 21692 29112
rect 21652 27674 21680 29106
rect 21824 28484 21876 28490
rect 21824 28426 21876 28432
rect 21836 28218 21864 28426
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 21640 27668 21692 27674
rect 21640 27610 21692 27616
rect 21928 27470 21956 29294
rect 22112 28966 22140 29600
rect 22192 29582 22244 29588
rect 22296 28994 22324 30194
rect 22388 30190 22416 30670
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22480 29850 22508 30874
rect 22468 29844 22520 29850
rect 22468 29786 22520 29792
rect 22572 29170 22600 31214
rect 22652 30592 22704 30598
rect 22652 30534 22704 30540
rect 22664 29850 22692 30534
rect 22756 30258 22784 33934
rect 22848 33930 22876 34342
rect 23216 34202 23244 34546
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 22836 33924 22888 33930
rect 22836 33866 22888 33872
rect 23492 33658 23520 34682
rect 24504 34542 24532 35022
rect 23572 34536 23624 34542
rect 23572 34478 23624 34484
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 23480 33652 23532 33658
rect 23480 33594 23532 33600
rect 23584 33538 23612 34478
rect 24688 34066 24716 35158
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 24964 34610 24992 34886
rect 24952 34604 25004 34610
rect 24952 34546 25004 34552
rect 25136 34536 25188 34542
rect 25136 34478 25188 34484
rect 24952 34400 25004 34406
rect 24952 34342 25004 34348
rect 24216 34060 24268 34066
rect 24216 34002 24268 34008
rect 24676 34060 24728 34066
rect 24676 34002 24728 34008
rect 23492 33510 23612 33538
rect 23388 33312 23440 33318
rect 23388 33254 23440 33260
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 23112 32360 23164 32366
rect 23112 32302 23164 32308
rect 22744 30252 22796 30258
rect 22744 30194 22796 30200
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 22652 29844 22704 29850
rect 22652 29786 22704 29792
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22204 28966 22324 28994
rect 22100 28960 22152 28966
rect 22100 28902 22152 28908
rect 22112 28626 22140 28902
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 22020 28082 22048 28358
rect 22112 28150 22140 28562
rect 22100 28144 22152 28150
rect 22100 28086 22152 28092
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22204 27656 22232 28966
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22296 28082 22324 28358
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22020 27628 22232 27656
rect 22284 27668 22336 27674
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 21652 26314 21680 27406
rect 21928 26330 21956 27406
rect 22020 26994 22048 27628
rect 22284 27610 22336 27616
rect 22190 27024 22246 27033
rect 22008 26988 22060 26994
rect 22190 26959 22192 26968
rect 22008 26930 22060 26936
rect 22244 26959 22246 26968
rect 22192 26930 22244 26936
rect 22100 26512 22152 26518
rect 22100 26454 22152 26460
rect 22112 26330 22140 26454
rect 22296 26450 22324 27610
rect 22572 27538 22600 29106
rect 22560 27532 22612 27538
rect 22560 27474 22612 27480
rect 22468 27464 22520 27470
rect 22468 27406 22520 27412
rect 22480 26586 22508 27406
rect 22756 26926 22784 30194
rect 23032 29578 23060 30194
rect 23124 29646 23152 32302
rect 23216 32230 23244 32710
rect 23400 32570 23428 33254
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23204 32224 23256 32230
rect 23204 32166 23256 32172
rect 23388 30184 23440 30190
rect 23388 30126 23440 30132
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23020 29572 23072 29578
rect 23020 29514 23072 29520
rect 23124 28994 23152 29582
rect 23032 28966 23152 28994
rect 23032 28694 23060 28966
rect 23020 28688 23072 28694
rect 23020 28630 23072 28636
rect 22836 27328 22888 27334
rect 22834 27296 22836 27305
rect 22888 27296 22890 27305
rect 22834 27231 22890 27240
rect 22744 26920 22796 26926
rect 22744 26862 22796 26868
rect 22848 26858 22876 27231
rect 22836 26852 22888 26858
rect 22836 26794 22888 26800
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 21640 26308 21692 26314
rect 21928 26302 22140 26330
rect 21640 26250 21692 26256
rect 23296 26240 23348 26246
rect 23296 26182 23348 26188
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22204 24834 22232 25842
rect 23308 25770 23336 26182
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22388 25362 22416 25638
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22112 24818 22232 24834
rect 22100 24812 22232 24818
rect 22152 24806 22232 24812
rect 22100 24754 22152 24760
rect 22112 24138 22140 24754
rect 22664 24682 22692 25162
rect 22744 25152 22796 25158
rect 22744 25094 22796 25100
rect 22756 24750 22784 25094
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22112 23730 22140 24074
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 23050 21956 23462
rect 22756 23186 22784 24686
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21836 21622 21864 22918
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 22020 20602 22048 22510
rect 23216 22030 23244 23054
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 23020 21480 23072 21486
rect 23020 21422 23072 21428
rect 22296 20602 22324 21422
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 21010 22416 21286
rect 23032 21146 23060 21422
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21928 20262 21956 20402
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 22020 19174 22048 20538
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22204 19378 22232 20266
rect 22756 19922 22784 20266
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22388 19514 22416 19722
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 23032 19446 23060 20198
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 22112 18358 22140 18634
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22204 18290 22232 19314
rect 23032 18630 23060 19382
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21836 15570 21864 16390
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21836 14006 21864 15030
rect 21928 15026 21956 16050
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21928 13818 21956 14962
rect 21836 13790 21956 13818
rect 21836 12850 21864 13790
rect 22020 13326 22048 17002
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22112 16046 22140 16594
rect 22204 16574 22232 17206
rect 22940 17202 22968 17614
rect 23032 17610 23060 18566
rect 23216 18222 23244 21966
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 22928 17196 22980 17202
rect 22928 17138 22980 17144
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 22204 16546 22324 16574
rect 22100 16040 22152 16046
rect 22152 15988 22232 15994
rect 22100 15982 22232 15988
rect 22112 15966 22232 15982
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22112 15570 22140 15846
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22204 15026 22232 15966
rect 22296 15706 22324 16546
rect 23308 16250 23336 17138
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 23112 15428 23164 15434
rect 23112 15370 23164 15376
rect 23124 15162 23152 15370
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 22204 12442 22232 13194
rect 22296 12918 22324 14214
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22480 12986 22508 13330
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 20548 12406 20668 12434
rect 21468 12406 21588 12434
rect 22192 12436 22244 12442
rect 20548 4078 20576 12406
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20640 4282 20668 4558
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 21008 4146 21036 4422
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 19996 3590 20484 3618
rect 19720 3466 19932 3482
rect 19708 3460 19944 3466
rect 19760 3454 19892 3460
rect 19708 3402 19760 3408
rect 19892 3402 19944 3408
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3074 19472 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 3074 20024 3590
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 19444 3046 19656 3074
rect 19628 2990 19656 3046
rect 19904 3046 20024 3074
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19904 2530 19932 3046
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19352 2502 19932 2530
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19352 800 19380 2502
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2926
rect 20364 2922 20392 3470
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20732 2650 20760 4014
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20824 3534 20852 3878
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 21468 2650 21496 12406
rect 22192 12378 22244 12384
rect 22572 12238 22600 14350
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 14006 22968 14214
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21560 3738 21588 4082
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 22112 3534 22140 3878
rect 22204 3738 22232 4626
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22468 4548 22520 4554
rect 22468 4490 22520 4496
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20640 800 20668 2314
rect 21928 800 21956 2994
rect 22296 2514 22324 4422
rect 22480 4146 22508 4490
rect 22572 4146 22600 4558
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22480 2446 22508 2858
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22572 800 22600 2858
rect 22756 2446 22784 4422
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22940 3058 22968 3470
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 23124 2990 23152 3878
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 23216 800 23244 2314
rect 23400 2038 23428 30126
rect 23492 28762 23520 33510
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 23584 31958 23612 32982
rect 23572 31952 23624 31958
rect 23572 31894 23624 31900
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 23492 28082 23520 28698
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23480 24880 23532 24886
rect 23480 24822 23532 24828
rect 23492 24410 23520 24822
rect 23480 24404 23532 24410
rect 23480 24346 23532 24352
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 21622 23520 22918
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23492 20602 23520 20878
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23676 18766 23704 31758
rect 24228 31278 24256 34002
rect 24676 33924 24728 33930
rect 24676 33866 24728 33872
rect 24688 33658 24716 33866
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 24308 33448 24360 33454
rect 24308 33390 24360 33396
rect 24216 31272 24268 31278
rect 24216 31214 24268 31220
rect 24228 30802 24256 31214
rect 24216 30796 24268 30802
rect 24216 30738 24268 30744
rect 24228 30598 24256 30738
rect 24216 30592 24268 30598
rect 24216 30534 24268 30540
rect 24320 30122 24348 33390
rect 24964 32910 24992 34342
rect 25148 33930 25176 34478
rect 25136 33924 25188 33930
rect 25136 33866 25188 33872
rect 25136 33312 25188 33318
rect 25136 33254 25188 33260
rect 25148 33114 25176 33254
rect 25136 33108 25188 33114
rect 25136 33050 25188 33056
rect 24952 32904 25004 32910
rect 24952 32846 25004 32852
rect 24584 32496 24636 32502
rect 24584 32438 24636 32444
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 24412 31260 24440 31622
rect 24504 31414 24532 31622
rect 24492 31408 24544 31414
rect 24492 31350 24544 31356
rect 24492 31272 24544 31278
rect 24412 31232 24492 31260
rect 24492 31214 24544 31220
rect 24492 30388 24544 30394
rect 24492 30330 24544 30336
rect 24308 30116 24360 30122
rect 24308 30058 24360 30064
rect 24308 29776 24360 29782
rect 24308 29718 24360 29724
rect 24320 29238 24348 29718
rect 24308 29232 24360 29238
rect 24308 29174 24360 29180
rect 24400 28552 24452 28558
rect 24400 28494 24452 28500
rect 24412 28150 24440 28494
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24228 26586 24256 26930
rect 24216 26580 24268 26586
rect 24216 26522 24268 26528
rect 23756 26308 23808 26314
rect 23756 26250 23808 26256
rect 23768 25974 23796 26250
rect 23756 25968 23808 25974
rect 23756 25910 23808 25916
rect 23768 25498 23796 25910
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23860 16574 23888 25842
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24136 20534 24164 22510
rect 24320 22098 24348 22510
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24136 19990 24164 20470
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24320 17882 24348 18702
rect 24400 18692 24452 18698
rect 24400 18634 24452 18640
rect 24308 17876 24360 17882
rect 24308 17818 24360 17824
rect 24320 17338 24348 17818
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24320 17202 24348 17274
rect 24308 17196 24360 17202
rect 24308 17138 24360 17144
rect 24412 17134 24440 18634
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16794 24440 16934
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 23860 16546 23980 16574
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23860 16114 23888 16390
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23584 15706 23612 15846
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23676 2446 23704 3674
rect 23768 2650 23796 4558
rect 23952 2650 23980 16546
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 24228 16046 24256 16458
rect 24216 16040 24268 16046
rect 24216 15982 24268 15988
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24412 15706 24440 15982
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 24504 2496 24532 30330
rect 24596 29170 24624 32438
rect 24964 32434 24992 32846
rect 25148 32502 25176 33050
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25240 32609 25268 32846
rect 25226 32600 25282 32609
rect 25226 32535 25282 32544
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 24674 31920 24730 31929
rect 24674 31855 24730 31864
rect 24768 31884 24820 31890
rect 24688 31822 24716 31855
rect 24768 31826 24820 31832
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 24780 30054 24808 31826
rect 25332 31754 25360 38898
rect 25976 38826 26004 38898
rect 25964 38820 26016 38826
rect 25964 38762 26016 38768
rect 26068 37806 26096 45426
rect 27344 45416 27396 45422
rect 27344 45358 27396 45364
rect 26148 39092 26200 39098
rect 26148 39034 26200 39040
rect 26160 38350 26188 39034
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 26160 37874 26188 38286
rect 26332 38208 26384 38214
rect 26332 38150 26384 38156
rect 26148 37868 26200 37874
rect 26148 37810 26200 37816
rect 25412 37800 25464 37806
rect 25412 37742 25464 37748
rect 26056 37800 26108 37806
rect 26056 37742 26108 37748
rect 25240 31726 25360 31754
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 24688 29170 24716 29514
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24768 28960 24820 28966
rect 24768 28902 24820 28908
rect 24780 28490 24808 28902
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24872 28218 24900 30602
rect 25044 30592 25096 30598
rect 25044 30534 25096 30540
rect 25056 30258 25084 30534
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24964 29850 24992 30126
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 24964 29714 24992 29786
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 25148 28626 25176 28902
rect 25136 28620 25188 28626
rect 25136 28562 25188 28568
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24860 28212 24912 28218
rect 24860 28154 24912 28160
rect 24780 27674 24808 28154
rect 24768 27668 24820 27674
rect 24768 27610 24820 27616
rect 24872 27470 24900 28154
rect 24952 28144 25004 28150
rect 24952 28086 25004 28092
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 24964 27334 24992 28086
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24688 26382 24716 26794
rect 24872 26382 24900 26862
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24872 25906 24900 26318
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24780 24750 24808 25094
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24872 24682 24900 25842
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24964 23186 24992 27270
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25044 26308 25096 26314
rect 25044 26250 25096 26256
rect 25056 25906 25084 26250
rect 25044 25900 25096 25906
rect 25044 25842 25096 25848
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 25056 24682 25084 25230
rect 25148 24818 25176 26726
rect 25240 26602 25268 31726
rect 25320 30388 25372 30394
rect 25320 30330 25372 30336
rect 25332 26738 25360 30330
rect 25424 26976 25452 37742
rect 26160 37262 26188 37810
rect 26148 37256 26200 37262
rect 26148 37198 26200 37204
rect 25780 36168 25832 36174
rect 25780 36110 25832 36116
rect 25688 36032 25740 36038
rect 25688 35974 25740 35980
rect 25700 35766 25728 35974
rect 25688 35760 25740 35766
rect 25688 35702 25740 35708
rect 25792 34610 25820 36110
rect 26344 35068 26372 38150
rect 27356 37806 27384 45358
rect 28632 44872 28684 44878
rect 28632 44814 28684 44820
rect 26792 37800 26844 37806
rect 26792 37742 26844 37748
rect 27344 37800 27396 37806
rect 27344 37742 27396 37748
rect 26700 37188 26752 37194
rect 26700 37130 26752 37136
rect 26424 36576 26476 36582
rect 26424 36518 26476 36524
rect 26516 36576 26568 36582
rect 26516 36518 26568 36524
rect 26436 35698 26464 36518
rect 26528 36242 26556 36518
rect 26516 36236 26568 36242
rect 26516 36178 26568 36184
rect 26608 36168 26660 36174
rect 26608 36110 26660 36116
rect 26620 35834 26648 36110
rect 26608 35828 26660 35834
rect 26608 35770 26660 35776
rect 26424 35692 26476 35698
rect 26424 35634 26476 35640
rect 26436 35222 26464 35634
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 26424 35216 26476 35222
rect 26424 35158 26476 35164
rect 26344 35040 26464 35068
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25964 34400 26016 34406
rect 25964 34342 26016 34348
rect 25872 33516 25924 33522
rect 25792 33476 25872 33504
rect 25792 32881 25820 33476
rect 25872 33458 25924 33464
rect 25872 32972 25924 32978
rect 25872 32914 25924 32920
rect 25778 32872 25834 32881
rect 25778 32807 25780 32816
rect 25832 32807 25834 32816
rect 25780 32778 25832 32784
rect 25884 32366 25912 32914
rect 25872 32360 25924 32366
rect 25872 32302 25924 32308
rect 25504 32020 25556 32026
rect 25504 31962 25556 31968
rect 25516 31482 25544 31962
rect 25976 31890 26004 34342
rect 26148 33992 26200 33998
rect 26148 33934 26200 33940
rect 26160 33862 26188 33934
rect 26148 33856 26200 33862
rect 26148 33798 26200 33804
rect 26160 33454 26188 33798
rect 26148 33448 26200 33454
rect 26148 33390 26200 33396
rect 26056 33108 26108 33114
rect 26056 33050 26108 33056
rect 26068 32502 26096 33050
rect 26160 32910 26188 33390
rect 26240 32972 26292 32978
rect 26240 32914 26292 32920
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 26252 32774 26280 32914
rect 26240 32768 26292 32774
rect 26240 32710 26292 32716
rect 26056 32496 26108 32502
rect 26056 32438 26108 32444
rect 25964 31884 26016 31890
rect 25964 31826 26016 31832
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25504 31476 25556 31482
rect 25504 31418 25556 31424
rect 25700 30938 25728 31758
rect 25780 31748 25832 31754
rect 25780 31690 25832 31696
rect 25792 31142 25820 31690
rect 25976 31414 26004 31826
rect 25964 31408 26016 31414
rect 25964 31350 26016 31356
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25688 30932 25740 30938
rect 25688 30874 25740 30880
rect 25688 30796 25740 30802
rect 25688 30738 25740 30744
rect 25700 29714 25728 30738
rect 25792 30734 25820 31078
rect 26068 30802 26096 32438
rect 26056 30796 26108 30802
rect 26056 30738 26108 30744
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25688 29708 25740 29714
rect 25688 29650 25740 29656
rect 25792 29646 25820 30670
rect 26252 30122 26280 32710
rect 26436 31668 26464 35040
rect 26528 35018 26556 35430
rect 26516 35012 26568 35018
rect 26516 34954 26568 34960
rect 26528 34678 26556 34954
rect 26516 34672 26568 34678
rect 26516 34614 26568 34620
rect 26528 34202 26556 34614
rect 26516 34196 26568 34202
rect 26516 34138 26568 34144
rect 26620 34082 26648 35770
rect 26528 34066 26648 34082
rect 26516 34060 26648 34066
rect 26568 34054 26648 34060
rect 26516 34002 26568 34008
rect 26712 32178 26740 37130
rect 26804 32298 26832 37742
rect 27528 36848 27580 36854
rect 27528 36790 27580 36796
rect 27540 36718 27568 36790
rect 26976 36712 27028 36718
rect 26976 36654 27028 36660
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 26988 36378 27016 36654
rect 26976 36372 27028 36378
rect 26976 36314 27028 36320
rect 27436 36236 27488 36242
rect 27436 36178 27488 36184
rect 27448 35494 27476 36178
rect 26976 35488 27028 35494
rect 26976 35430 27028 35436
rect 27436 35488 27488 35494
rect 27436 35430 27488 35436
rect 26988 35086 27016 35430
rect 26976 35080 27028 35086
rect 26976 35022 27028 35028
rect 27344 34944 27396 34950
rect 27344 34886 27396 34892
rect 26884 34604 26936 34610
rect 26884 34546 26936 34552
rect 26896 33522 26924 34546
rect 27252 34468 27304 34474
rect 27252 34410 27304 34416
rect 27264 34066 27292 34410
rect 27252 34060 27304 34066
rect 27252 34002 27304 34008
rect 27068 33856 27120 33862
rect 27068 33798 27120 33804
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 27080 33590 27108 33798
rect 27172 33658 27200 33798
rect 27160 33652 27212 33658
rect 27160 33594 27212 33600
rect 27068 33584 27120 33590
rect 27068 33526 27120 33532
rect 27264 33522 27292 34002
rect 27356 33658 27384 34886
rect 27344 33652 27396 33658
rect 27344 33594 27396 33600
rect 26884 33516 26936 33522
rect 26884 33458 26936 33464
rect 27252 33516 27304 33522
rect 27252 33458 27304 33464
rect 26896 32978 26924 33458
rect 26976 33312 27028 33318
rect 26976 33254 27028 33260
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 26792 32292 26844 32298
rect 26792 32234 26844 32240
rect 26712 32150 26924 32178
rect 26792 31816 26844 31822
rect 26792 31758 26844 31764
rect 26436 31640 26740 31668
rect 26436 31482 26464 31640
rect 26424 31476 26476 31482
rect 26424 31418 26476 31424
rect 26608 31408 26660 31414
rect 26608 31350 26660 31356
rect 26424 31340 26476 31346
rect 26424 31282 26476 31288
rect 26436 30938 26464 31282
rect 26424 30932 26476 30938
rect 26424 30874 26476 30880
rect 26424 30320 26476 30326
rect 26424 30262 26476 30268
rect 26240 30116 26292 30122
rect 26240 30058 26292 30064
rect 26240 29844 26292 29850
rect 26240 29786 26292 29792
rect 26056 29708 26108 29714
rect 26056 29650 26108 29656
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29170 25912 29446
rect 25872 29164 25924 29170
rect 25872 29106 25924 29112
rect 25964 29164 26016 29170
rect 25964 29106 26016 29112
rect 25976 29050 26004 29106
rect 25884 29022 26004 29050
rect 25688 28960 25740 28966
rect 25688 28902 25740 28908
rect 25700 28762 25728 28902
rect 25688 28756 25740 28762
rect 25688 28698 25740 28704
rect 25884 27878 25912 29022
rect 26068 28642 26096 29650
rect 26148 29572 26200 29578
rect 26148 29514 26200 29520
rect 26160 28762 26188 29514
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 26252 28642 26280 29786
rect 26068 28614 26188 28642
rect 26252 28614 26372 28642
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 25872 27872 25924 27878
rect 25870 27840 25872 27849
rect 25924 27840 25926 27849
rect 25870 27775 25926 27784
rect 25780 27600 25832 27606
rect 25780 27542 25832 27548
rect 25792 27062 25820 27542
rect 25884 27452 25912 27775
rect 25976 27606 26004 28426
rect 25964 27600 26016 27606
rect 25964 27542 26016 27548
rect 25884 27424 26004 27452
rect 25780 27056 25832 27062
rect 25780 26998 25832 27004
rect 25424 26948 25728 26976
rect 25332 26710 25544 26738
rect 25240 26574 25452 26602
rect 25228 26512 25280 26518
rect 25228 26454 25280 26460
rect 25320 26512 25372 26518
rect 25320 26454 25372 26460
rect 25240 24818 25268 26454
rect 25332 25770 25360 26454
rect 25424 26246 25452 26574
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25320 25764 25372 25770
rect 25320 25706 25372 25712
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25044 24676 25096 24682
rect 25044 24618 25096 24624
rect 25516 24614 25544 26710
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25136 24132 25188 24138
rect 25136 24074 25188 24080
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 25056 19922 25084 20198
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24688 18630 24716 19246
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24688 18290 24716 18566
rect 24872 18358 24900 19790
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24964 18290 24992 18566
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 25148 18170 25176 24074
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25332 23050 25360 23462
rect 25412 23180 25464 23186
rect 25464 23140 25544 23168
rect 25412 23122 25464 23128
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25516 22030 25544 23140
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25516 21554 25544 21966
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25412 20460 25464 20466
rect 25412 20402 25464 20408
rect 25424 19378 25452 20402
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25240 18834 25268 19110
rect 25516 18834 25544 19178
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 24872 18142 25176 18170
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24596 16590 24624 17070
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24688 16726 24716 16934
rect 24780 16726 24808 17274
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24768 16720 24820 16726
rect 24768 16662 24820 16668
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24872 13530 24900 18142
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24964 16590 24992 17138
rect 25044 17060 25096 17066
rect 25044 17002 25096 17008
rect 25056 16658 25084 17002
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 25056 16250 25084 16594
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 25320 16176 25372 16182
rect 25320 16118 25372 16124
rect 25332 15706 25360 16118
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25240 15026 25268 15438
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 25608 5098 25636 25230
rect 25700 19174 25728 26948
rect 25872 25696 25924 25702
rect 25872 25638 25924 25644
rect 25780 25220 25832 25226
rect 25780 25162 25832 25168
rect 25792 24070 25820 25162
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25884 22234 25912 25638
rect 25872 22228 25924 22234
rect 25872 22170 25924 22176
rect 25976 20942 26004 27424
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 26068 26790 26096 26930
rect 26160 26858 26188 28614
rect 26240 28484 26292 28490
rect 26240 28426 26292 28432
rect 26252 28082 26280 28426
rect 26240 28076 26292 28082
rect 26240 28018 26292 28024
rect 26344 27606 26372 28614
rect 26332 27600 26384 27606
rect 26332 27542 26384 27548
rect 26148 26852 26200 26858
rect 26148 26794 26200 26800
rect 26056 26784 26108 26790
rect 26056 26726 26108 26732
rect 26068 26042 26096 26726
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 26436 25294 26464 30262
rect 26516 28688 26568 28694
rect 26620 28665 26648 31350
rect 26516 28630 26568 28636
rect 26606 28656 26662 28665
rect 26528 26586 26556 28630
rect 26606 28591 26662 28600
rect 26516 26580 26568 26586
rect 26516 26522 26568 26528
rect 26528 26246 26556 26522
rect 26516 26240 26568 26246
rect 26516 26182 26568 26188
rect 26608 26036 26660 26042
rect 26608 25978 26660 25984
rect 26620 25770 26648 25978
rect 26608 25764 26660 25770
rect 26608 25706 26660 25712
rect 26620 25498 26648 25706
rect 26608 25492 26660 25498
rect 26608 25434 26660 25440
rect 26424 25288 26476 25294
rect 26424 25230 26476 25236
rect 26436 24886 26464 25230
rect 26424 24880 26476 24886
rect 26424 24822 26476 24828
rect 26436 24206 26464 24822
rect 26608 24404 26660 24410
rect 26608 24346 26660 24352
rect 26620 24206 26648 24346
rect 26424 24200 26476 24206
rect 26424 24142 26476 24148
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 26424 24064 26476 24070
rect 26424 24006 26476 24012
rect 26160 23730 26188 24006
rect 26436 23730 26464 24006
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26620 23322 26648 24142
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25976 17202 26004 20878
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26344 19786 26372 20198
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 26240 19440 26292 19446
rect 26240 19382 26292 19388
rect 26252 17270 26280 19382
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 25964 17196 26016 17202
rect 25964 17138 26016 17144
rect 26056 16992 26108 16998
rect 26056 16934 26108 16940
rect 26068 15502 26096 16934
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 25596 5092 25648 5098
rect 25596 5034 25648 5040
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 24412 2468 24532 2496
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 24412 2310 24440 2468
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 24400 2304 24452 2310
rect 24400 2246 24452 2252
rect 23388 2032 23440 2038
rect 23388 1974 23440 1980
rect 24504 800 24532 2314
rect 25148 800 25176 3674
rect 25332 2514 25360 4422
rect 25412 3528 25464 3534
rect 25412 3470 25464 3476
rect 25424 2650 25452 3470
rect 25608 3058 25636 4626
rect 26712 4146 26740 31640
rect 26804 25906 26832 31758
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 26896 22094 26924 32150
rect 26988 31822 27016 33254
rect 27264 32910 27292 33458
rect 27252 32904 27304 32910
rect 27252 32846 27304 32852
rect 27448 32774 27476 35430
rect 27436 32768 27488 32774
rect 27436 32710 27488 32716
rect 27540 32586 27568 36654
rect 28448 35624 28500 35630
rect 28448 35566 28500 35572
rect 27804 35012 27856 35018
rect 27804 34954 27856 34960
rect 27816 33658 27844 34954
rect 27988 34740 28040 34746
rect 27988 34682 28040 34688
rect 27804 33652 27856 33658
rect 27804 33594 27856 33600
rect 27804 32972 27856 32978
rect 27804 32914 27856 32920
rect 27816 32881 27844 32914
rect 27802 32872 27858 32881
rect 28000 32842 28028 34682
rect 28460 33998 28488 35566
rect 28448 33992 28500 33998
rect 28448 33934 28500 33940
rect 28460 33810 28488 33934
rect 28276 33782 28488 33810
rect 28080 33448 28132 33454
rect 28080 33390 28132 33396
rect 28092 33046 28120 33390
rect 28172 33312 28224 33318
rect 28172 33254 28224 33260
rect 28080 33040 28132 33046
rect 28080 32982 28132 32988
rect 27802 32807 27858 32816
rect 27988 32836 28040 32842
rect 27988 32778 28040 32784
rect 27448 32558 27568 32586
rect 27066 32192 27122 32201
rect 27066 32127 27122 32136
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 27080 31754 27108 32127
rect 27068 31748 27120 31754
rect 27068 31690 27120 31696
rect 27068 30048 27120 30054
rect 27068 29990 27120 29996
rect 27344 30048 27396 30054
rect 27344 29990 27396 29996
rect 27080 29578 27108 29990
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 27252 29640 27304 29646
rect 27252 29582 27304 29588
rect 27068 29572 27120 29578
rect 26988 29532 27068 29560
rect 26988 28422 27016 29532
rect 27068 29514 27120 29520
rect 27068 29096 27120 29102
rect 27068 29038 27120 29044
rect 27080 28626 27108 29038
rect 27068 28620 27120 28626
rect 27068 28562 27120 28568
rect 26976 28416 27028 28422
rect 26976 28358 27028 28364
rect 26988 28098 27016 28358
rect 27172 28218 27200 29582
rect 27264 29510 27292 29582
rect 27252 29504 27304 29510
rect 27252 29446 27304 29452
rect 27264 28558 27292 29446
rect 27356 29306 27384 29990
rect 27344 29300 27396 29306
rect 27344 29242 27396 29248
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27160 28212 27212 28218
rect 27160 28154 27212 28160
rect 26988 28070 27200 28098
rect 26976 27600 27028 27606
rect 26976 27542 27028 27548
rect 26988 23526 27016 27542
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 27080 26518 27108 27406
rect 27172 27334 27200 28070
rect 27264 27606 27292 28358
rect 27252 27600 27304 27606
rect 27252 27542 27304 27548
rect 27356 27538 27384 29242
rect 27448 28218 27476 32558
rect 27988 32496 28040 32502
rect 27988 32438 28040 32444
rect 28000 32298 28028 32438
rect 27528 32292 27580 32298
rect 27528 32234 27580 32240
rect 27988 32292 28040 32298
rect 27988 32234 28040 32240
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 27448 28082 27476 28154
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 27436 27600 27488 27606
rect 27436 27542 27488 27548
rect 27344 27532 27396 27538
rect 27344 27474 27396 27480
rect 27160 27328 27212 27334
rect 27160 27270 27212 27276
rect 27160 27056 27212 27062
rect 27160 26998 27212 27004
rect 27068 26512 27120 26518
rect 27068 26454 27120 26460
rect 27172 26382 27200 26998
rect 27448 26602 27476 27542
rect 27356 26586 27476 26602
rect 27344 26580 27476 26586
rect 27396 26574 27476 26580
rect 27344 26522 27396 26528
rect 27448 26382 27476 26574
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27436 25832 27488 25838
rect 27436 25774 27488 25780
rect 27160 25356 27212 25362
rect 27160 25298 27212 25304
rect 26976 23520 27028 23526
rect 26976 23462 27028 23468
rect 27068 22432 27120 22438
rect 27068 22374 27120 22380
rect 26804 22066 26924 22094
rect 26804 21010 26832 22066
rect 27080 21962 27108 22374
rect 27068 21956 27120 21962
rect 27068 21898 27120 21904
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26896 17678 26924 19858
rect 27080 18698 27108 20198
rect 27172 19922 27200 25298
rect 27448 25226 27476 25774
rect 27436 25220 27488 25226
rect 27436 25162 27488 25168
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27448 21146 27476 22578
rect 27436 21140 27488 21146
rect 27436 21082 27488 21088
rect 27448 20942 27476 21082
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 27448 20466 27476 20878
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27160 19916 27212 19922
rect 27160 19858 27212 19864
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 27172 19446 27200 19722
rect 27160 19440 27212 19446
rect 27160 19382 27212 19388
rect 27172 18902 27200 19382
rect 27160 18896 27212 18902
rect 27160 18838 27212 18844
rect 27068 18692 27120 18698
rect 27068 18634 27120 18640
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 26884 17196 26936 17202
rect 27160 17196 27212 17202
rect 26884 17138 26936 17144
rect 27080 17156 27160 17184
rect 26896 16658 26924 17138
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 27080 16590 27108 17156
rect 27160 17138 27212 17144
rect 27172 16658 27292 16674
rect 27160 16652 27292 16658
rect 27212 16646 27292 16652
rect 27160 16594 27212 16600
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 26700 4140 26752 4146
rect 26700 4082 26752 4088
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 26252 3398 26280 3878
rect 26330 3632 26386 3641
rect 26620 3602 26924 3618
rect 26330 3567 26386 3576
rect 26608 3596 26936 3602
rect 26344 3398 26372 3567
rect 26660 3590 26884 3596
rect 26608 3538 26660 3544
rect 26884 3538 26936 3544
rect 26976 3460 27028 3466
rect 26976 3402 27028 3408
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 26056 3052 26108 3058
rect 26056 2994 26108 3000
rect 26068 2854 26096 2994
rect 26988 2854 27016 3402
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 26976 2848 27028 2854
rect 26976 2790 27028 2796
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 27080 2582 27108 16526
rect 27264 4690 27292 16646
rect 27252 4684 27304 4690
rect 27252 4626 27304 4632
rect 27264 3534 27292 4626
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 27356 3738 27384 4082
rect 27540 3942 27568 32234
rect 27804 32224 27856 32230
rect 27804 32166 27856 32172
rect 27816 31822 27844 32166
rect 28000 31958 28028 32234
rect 27988 31952 28040 31958
rect 28080 31952 28132 31958
rect 27988 31894 28040 31900
rect 28078 31920 28080 31929
rect 28132 31920 28134 31929
rect 28078 31855 28134 31864
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 27620 30184 27672 30190
rect 27620 30126 27672 30132
rect 27632 29850 27660 30126
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 27712 29164 27764 29170
rect 27712 29106 27764 29112
rect 27620 27872 27672 27878
rect 27620 27814 27672 27820
rect 27632 26382 27660 27814
rect 27620 26376 27672 26382
rect 27620 26318 27672 26324
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27632 24206 27660 25774
rect 27724 24682 27752 29106
rect 27816 28762 27844 31758
rect 27896 31272 27948 31278
rect 27896 31214 27948 31220
rect 27804 28756 27856 28762
rect 27804 28698 27856 28704
rect 27804 28008 27856 28014
rect 27908 27962 27936 31214
rect 28080 29572 28132 29578
rect 28080 29514 28132 29520
rect 27856 27956 27936 27962
rect 27804 27950 27936 27956
rect 27816 27934 27936 27950
rect 27908 26790 27936 27934
rect 27988 27872 28040 27878
rect 27986 27840 27988 27849
rect 28040 27840 28042 27849
rect 27986 27775 28042 27784
rect 28092 27674 28120 29514
rect 28080 27668 28132 27674
rect 28080 27610 28132 27616
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27804 26512 27856 26518
rect 27804 26454 27856 26460
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27632 23118 27660 24142
rect 27816 23866 27844 26454
rect 27896 25968 27948 25974
rect 27896 25910 27948 25916
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27632 22098 27660 23054
rect 27712 23044 27764 23050
rect 27712 22986 27764 22992
rect 27724 22778 27752 22986
rect 27712 22772 27764 22778
rect 27712 22714 27764 22720
rect 27908 22710 27936 25910
rect 28092 25498 28120 27610
rect 28080 25492 28132 25498
rect 28080 25434 28132 25440
rect 28092 24750 28120 25434
rect 28080 24744 28132 24750
rect 28080 24686 28132 24692
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 28000 24274 28028 24550
rect 27988 24268 28040 24274
rect 27988 24210 28040 24216
rect 28000 23866 28028 24210
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 28092 23798 28120 24142
rect 28080 23792 28132 23798
rect 28080 23734 28132 23740
rect 28080 23520 28132 23526
rect 28080 23462 28132 23468
rect 28092 23050 28120 23462
rect 28080 23044 28132 23050
rect 28080 22986 28132 22992
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27620 22092 27672 22098
rect 28184 22094 28212 33254
rect 28276 29730 28304 33782
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28460 33318 28488 33458
rect 28540 33448 28592 33454
rect 28540 33390 28592 33396
rect 28448 33312 28500 33318
rect 28448 33254 28500 33260
rect 28460 31414 28488 33254
rect 28552 33046 28580 33390
rect 28540 33040 28592 33046
rect 28540 32982 28592 32988
rect 28540 32768 28592 32774
rect 28540 32710 28592 32716
rect 28552 32570 28580 32710
rect 28540 32564 28592 32570
rect 28540 32506 28592 32512
rect 28552 32230 28580 32506
rect 28540 32224 28592 32230
rect 28540 32166 28592 32172
rect 28644 31958 28672 44814
rect 29932 41414 29960 46854
rect 29932 41386 30052 41414
rect 29920 35624 29972 35630
rect 29920 35566 29972 35572
rect 29932 35290 29960 35566
rect 29920 35284 29972 35290
rect 29920 35226 29972 35232
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 28816 35012 28868 35018
rect 28816 34954 28868 34960
rect 28908 35012 28960 35018
rect 28908 34954 28960 34960
rect 28828 34746 28856 34954
rect 28816 34740 28868 34746
rect 28816 34682 28868 34688
rect 28920 34610 28948 34954
rect 29184 34944 29236 34950
rect 29184 34886 29236 34892
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 29196 34474 29224 34886
rect 29184 34468 29236 34474
rect 29184 34410 29236 34416
rect 29000 34060 29052 34066
rect 29000 34002 29052 34008
rect 29012 33658 29040 34002
rect 29000 33652 29052 33658
rect 29000 33594 29052 33600
rect 29012 33522 29040 33594
rect 29196 33522 29224 34410
rect 29552 34128 29604 34134
rect 29552 34070 29604 34076
rect 29368 33924 29420 33930
rect 29368 33866 29420 33872
rect 29380 33538 29408 33866
rect 29460 33584 29512 33590
rect 29380 33532 29460 33538
rect 29380 33526 29512 33532
rect 29000 33516 29052 33522
rect 29000 33458 29052 33464
rect 29184 33516 29236 33522
rect 29184 33458 29236 33464
rect 29380 33510 29500 33526
rect 29012 32910 29040 33458
rect 29092 33108 29144 33114
rect 29092 33050 29144 33056
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 28814 32600 28870 32609
rect 28814 32535 28870 32544
rect 28828 32502 28856 32535
rect 28816 32496 28868 32502
rect 29000 32496 29052 32502
rect 28816 32438 28868 32444
rect 28998 32464 29000 32473
rect 29052 32464 29054 32473
rect 28908 32428 28960 32434
rect 28998 32399 29054 32408
rect 28908 32370 28960 32376
rect 28920 32212 28948 32370
rect 28920 32184 29040 32212
rect 28632 31952 28684 31958
rect 28632 31894 28684 31900
rect 28448 31408 28500 31414
rect 28448 31350 28500 31356
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28356 30592 28408 30598
rect 28356 30534 28408 30540
rect 28368 30326 28396 30534
rect 28356 30320 28408 30326
rect 28356 30262 28408 30268
rect 28644 30122 28672 30670
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 29012 29850 29040 32184
rect 29104 31890 29132 33050
rect 29184 32836 29236 32842
rect 29184 32778 29236 32784
rect 29196 32366 29224 32778
rect 29380 32774 29408 33510
rect 29368 32768 29420 32774
rect 29368 32710 29420 32716
rect 29276 32564 29328 32570
rect 29276 32506 29328 32512
rect 29184 32360 29236 32366
rect 29184 32302 29236 32308
rect 29092 31884 29144 31890
rect 29092 31826 29144 31832
rect 29104 31142 29132 31826
rect 29196 31414 29224 32302
rect 29184 31408 29236 31414
rect 29184 31350 29236 31356
rect 29092 31136 29144 31142
rect 29092 31078 29144 31084
rect 29104 30138 29132 31078
rect 29104 30110 29224 30138
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 29104 29782 29132 29990
rect 29092 29776 29144 29782
rect 28276 29702 28396 29730
rect 29092 29718 29144 29724
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 27620 22034 27672 22040
rect 28092 22066 28212 22094
rect 28276 22094 28304 29582
rect 28368 29578 28396 29702
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 28644 28558 28672 29650
rect 28816 29640 28868 29646
rect 28816 29582 28868 29588
rect 28828 29306 28856 29582
rect 28816 29300 28868 29306
rect 28816 29242 28868 29248
rect 29000 29164 29052 29170
rect 29000 29106 29052 29112
rect 28908 28960 28960 28966
rect 28908 28902 28960 28908
rect 28722 28656 28778 28665
rect 28722 28591 28778 28600
rect 28632 28552 28684 28558
rect 28632 28494 28684 28500
rect 28448 28484 28500 28490
rect 28448 28426 28500 28432
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 28368 26790 28396 28018
rect 28356 26784 28408 26790
rect 28356 26726 28408 26732
rect 28460 25906 28488 28426
rect 28540 27940 28592 27946
rect 28540 27882 28592 27888
rect 28552 27674 28580 27882
rect 28540 27668 28592 27674
rect 28540 27610 28592 27616
rect 28540 26784 28592 26790
rect 28540 26726 28592 26732
rect 28552 26382 28580 26726
rect 28736 26518 28764 28591
rect 28920 28150 28948 28902
rect 28908 28144 28960 28150
rect 28908 28086 28960 28092
rect 29012 26926 29040 29106
rect 29196 27062 29224 30110
rect 29288 28082 29316 32506
rect 29380 31754 29408 32710
rect 29564 32570 29592 34070
rect 29644 33992 29696 33998
rect 29644 33934 29696 33940
rect 29656 32842 29684 33934
rect 29644 32836 29696 32842
rect 29644 32778 29696 32784
rect 29656 32570 29684 32778
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29644 32564 29696 32570
rect 29644 32506 29696 32512
rect 29460 32496 29512 32502
rect 29460 32438 29512 32444
rect 29642 32464 29698 32473
rect 29472 32298 29500 32438
rect 29642 32399 29698 32408
rect 29656 32366 29684 32399
rect 29644 32360 29696 32366
rect 29644 32302 29696 32308
rect 29460 32292 29512 32298
rect 29460 32234 29512 32240
rect 29380 31726 29500 31754
rect 29368 31408 29420 31414
rect 29368 31350 29420 31356
rect 29276 28076 29328 28082
rect 29276 28018 29328 28024
rect 29380 27470 29408 31350
rect 29472 29186 29500 31726
rect 29472 29158 29684 29186
rect 29748 29170 29776 35090
rect 29828 34944 29880 34950
rect 29828 34886 29880 34892
rect 29840 34202 29868 34886
rect 29828 34196 29880 34202
rect 29828 34138 29880 34144
rect 29828 33924 29880 33930
rect 29828 33866 29880 33872
rect 29840 33658 29868 33866
rect 29828 33652 29880 33658
rect 29828 33594 29880 33600
rect 29828 33040 29880 33046
rect 29828 32982 29880 32988
rect 29840 32298 29868 32982
rect 29828 32292 29880 32298
rect 29828 32234 29880 32240
rect 29840 29238 29868 32234
rect 29828 29232 29880 29238
rect 29828 29174 29880 29180
rect 29460 29096 29512 29102
rect 29460 29038 29512 29044
rect 29368 27464 29420 27470
rect 29368 27406 29420 27412
rect 29184 27056 29236 27062
rect 29184 26998 29236 27004
rect 29196 26926 29224 26998
rect 29380 26994 29408 27406
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29000 26920 29052 26926
rect 29000 26862 29052 26868
rect 29184 26920 29236 26926
rect 29184 26862 29236 26868
rect 28724 26512 28776 26518
rect 28724 26454 28776 26460
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28552 26042 28580 26318
rect 28632 26308 28684 26314
rect 28632 26250 28684 26256
rect 28540 26036 28592 26042
rect 28540 25978 28592 25984
rect 28644 25906 28672 26250
rect 28448 25900 28500 25906
rect 28448 25842 28500 25848
rect 28632 25900 28684 25906
rect 28632 25842 28684 25848
rect 28356 25696 28408 25702
rect 28356 25638 28408 25644
rect 28368 24954 28396 25638
rect 28356 24948 28408 24954
rect 28356 24890 28408 24896
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 28368 23730 28396 24210
rect 28460 24070 28488 25842
rect 29012 25498 29040 26862
rect 29000 25492 29052 25498
rect 29000 25434 29052 25440
rect 29368 25288 29420 25294
rect 29368 25230 29420 25236
rect 29380 24886 29408 25230
rect 29368 24880 29420 24886
rect 29368 24822 29420 24828
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28552 24206 28580 24754
rect 28632 24744 28684 24750
rect 28632 24686 28684 24692
rect 28644 24410 28672 24686
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28448 24064 28500 24070
rect 28448 24006 28500 24012
rect 28724 24064 28776 24070
rect 28724 24006 28776 24012
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28356 23724 28408 23730
rect 28356 23666 28408 23672
rect 28368 23118 28396 23666
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28460 22982 28488 23802
rect 28736 23730 28764 24006
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28816 23248 28868 23254
rect 28816 23190 28868 23196
rect 28724 23044 28776 23050
rect 28724 22986 28776 22992
rect 28448 22976 28500 22982
rect 28448 22918 28500 22924
rect 28736 22642 28764 22986
rect 28724 22636 28776 22642
rect 28724 22578 28776 22584
rect 28276 22066 28488 22094
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27724 21622 27752 21830
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 27986 19952 28042 19961
rect 27986 19887 28042 19896
rect 28000 19446 28028 19887
rect 27988 19440 28040 19446
rect 27988 19382 28040 19388
rect 28000 18766 28028 19382
rect 27988 18760 28040 18766
rect 27988 18702 28040 18708
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27632 17678 27660 18226
rect 28000 17678 28028 18702
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 27632 17338 27660 17614
rect 27620 17332 27672 17338
rect 27620 17274 27672 17280
rect 28092 16574 28120 22066
rect 28172 21616 28224 21622
rect 28172 21558 28224 21564
rect 28184 21146 28212 21558
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28184 19378 28212 20198
rect 28264 19916 28316 19922
rect 28264 19858 28316 19864
rect 28172 19372 28224 19378
rect 28172 19314 28224 19320
rect 28184 18766 28212 19314
rect 28172 18760 28224 18766
rect 28172 18702 28224 18708
rect 28184 17678 28212 18702
rect 28276 18698 28304 19858
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 28368 19514 28396 19790
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28264 18692 28316 18698
rect 28264 18634 28316 18640
rect 28276 18290 28304 18634
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28092 16546 28212 16574
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 28184 2650 28212 16546
rect 28460 6186 28488 22066
rect 28736 21690 28764 22578
rect 28828 21962 28856 23190
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 29104 22166 29132 22578
rect 29276 22432 29328 22438
rect 29276 22374 29328 22380
rect 29092 22160 29144 22166
rect 29092 22102 29144 22108
rect 29288 22030 29316 22374
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 28816 21956 28868 21962
rect 28816 21898 28868 21904
rect 28724 21684 28776 21690
rect 28724 21626 28776 21632
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28552 19514 28580 20334
rect 28724 20324 28776 20330
rect 28724 20266 28776 20272
rect 28540 19508 28592 19514
rect 28540 19450 28592 19456
rect 28736 19446 28764 20266
rect 28828 20058 28856 20334
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28816 19916 28868 19922
rect 28816 19858 28868 19864
rect 28724 19440 28776 19446
rect 28724 19382 28776 19388
rect 28736 18902 28764 19382
rect 28828 19378 28856 19858
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28816 19372 28868 19378
rect 28816 19314 28868 19320
rect 28724 18896 28776 18902
rect 28724 18838 28776 18844
rect 28828 17746 28856 19314
rect 28920 18766 28948 19654
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 29472 18426 29500 29038
rect 29552 27464 29604 27470
rect 29552 27406 29604 27412
rect 29564 26858 29592 27406
rect 29552 26852 29604 26858
rect 29552 26794 29604 26800
rect 29564 25906 29592 26794
rect 29552 25900 29604 25906
rect 29552 25842 29604 25848
rect 29564 22710 29592 25842
rect 29656 24614 29684 29158
rect 29736 29164 29788 29170
rect 29736 29106 29788 29112
rect 29920 29164 29972 29170
rect 29920 29106 29972 29112
rect 29932 28778 29960 29106
rect 29840 28762 29960 28778
rect 29736 28756 29788 28762
rect 29736 28698 29788 28704
rect 29828 28756 29960 28762
rect 29880 28750 29960 28756
rect 29828 28698 29880 28704
rect 29748 28422 29776 28698
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 29748 25430 29776 28358
rect 29920 28076 29972 28082
rect 29840 28036 29920 28064
rect 29840 27538 29868 28036
rect 29920 28018 29972 28024
rect 29828 27532 29880 27538
rect 29828 27474 29880 27480
rect 29840 26926 29868 27474
rect 29828 26920 29880 26926
rect 29828 26862 29880 26868
rect 29840 26586 29868 26862
rect 29828 26580 29880 26586
rect 29828 26522 29880 26528
rect 29736 25424 29788 25430
rect 29736 25366 29788 25372
rect 29644 24608 29696 24614
rect 29644 24550 29696 24556
rect 29736 23724 29788 23730
rect 29736 23666 29788 23672
rect 29748 23118 29776 23666
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29552 22704 29604 22710
rect 29552 22646 29604 22652
rect 29736 22568 29788 22574
rect 29840 22556 29868 26522
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 29932 24954 29960 25230
rect 29920 24948 29972 24954
rect 29920 24890 29972 24896
rect 29788 22528 29868 22556
rect 29736 22510 29788 22516
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 29460 18420 29512 18426
rect 29460 18362 29512 18368
rect 29656 18154 29684 18702
rect 29644 18148 29696 18154
rect 29644 18090 29696 18096
rect 28816 17740 28868 17746
rect 28816 17682 28868 17688
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28644 16794 28672 17614
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 29748 8838 29776 22510
rect 30024 20466 30052 41386
rect 30208 35290 30236 46922
rect 30944 41414 30972 46990
rect 31036 46986 31064 47110
rect 31024 46980 31076 46986
rect 31024 46922 31076 46928
rect 32232 46442 32260 49200
rect 38028 47410 38056 49200
rect 37292 47382 38056 47410
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34244 47252 34296 47258
rect 34244 47194 34296 47200
rect 32404 47116 32456 47122
rect 32404 47058 32456 47064
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 30760 41386 30972 41414
rect 30288 35624 30340 35630
rect 30288 35566 30340 35572
rect 30196 35284 30248 35290
rect 30196 35226 30248 35232
rect 30104 35080 30156 35086
rect 30104 35022 30156 35028
rect 30116 34746 30144 35022
rect 30104 34740 30156 34746
rect 30104 34682 30156 34688
rect 30300 34610 30328 35566
rect 30288 34604 30340 34610
rect 30288 34546 30340 34552
rect 30104 34400 30156 34406
rect 30104 34342 30156 34348
rect 30116 33930 30144 34342
rect 30104 33924 30156 33930
rect 30104 33866 30156 33872
rect 30300 33862 30328 34546
rect 30380 34400 30432 34406
rect 30380 34342 30432 34348
rect 30392 34066 30420 34342
rect 30380 34060 30432 34066
rect 30380 34002 30432 34008
rect 30288 33856 30340 33862
rect 30288 33798 30340 33804
rect 30196 33516 30248 33522
rect 30196 33458 30248 33464
rect 30104 32972 30156 32978
rect 30104 32914 30156 32920
rect 30116 32434 30144 32914
rect 30104 32428 30156 32434
rect 30104 32370 30156 32376
rect 30208 30734 30236 33458
rect 30300 33318 30328 33798
rect 30288 33312 30340 33318
rect 30288 33254 30340 33260
rect 30392 32910 30420 34002
rect 30380 32904 30432 32910
rect 30380 32846 30432 32852
rect 30472 31816 30524 31822
rect 30472 31758 30524 31764
rect 30196 30728 30248 30734
rect 30196 30670 30248 30676
rect 30208 28472 30236 30670
rect 30380 30592 30432 30598
rect 30380 30534 30432 30540
rect 30392 30326 30420 30534
rect 30380 30320 30432 30326
rect 30380 30262 30432 30268
rect 30380 29708 30432 29714
rect 30380 29650 30432 29656
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30300 28694 30328 29582
rect 30392 29306 30420 29650
rect 30380 29300 30432 29306
rect 30380 29242 30432 29248
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30288 28688 30340 28694
rect 30288 28630 30340 28636
rect 30288 28484 30340 28490
rect 30208 28444 30288 28472
rect 30288 28426 30340 28432
rect 30300 27606 30328 28426
rect 30392 27606 30420 29106
rect 30288 27600 30340 27606
rect 30288 27542 30340 27548
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 30300 26518 30328 27542
rect 30484 26858 30512 31758
rect 30564 31408 30616 31414
rect 30564 31350 30616 31356
rect 30576 28014 30604 31350
rect 30656 30184 30708 30190
rect 30656 30126 30708 30132
rect 30668 29306 30696 30126
rect 30656 29300 30708 29306
rect 30656 29242 30708 29248
rect 30564 28008 30616 28014
rect 30564 27950 30616 27956
rect 30576 27674 30604 27950
rect 30564 27668 30616 27674
rect 30564 27610 30616 27616
rect 30472 26852 30524 26858
rect 30472 26794 30524 26800
rect 30288 26512 30340 26518
rect 30288 26454 30340 26460
rect 30484 26450 30512 26794
rect 30472 26444 30524 26450
rect 30472 26386 30524 26392
rect 30104 25832 30156 25838
rect 30104 25774 30156 25780
rect 30116 25294 30144 25774
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30472 25152 30524 25158
rect 30472 25094 30524 25100
rect 30380 24880 30432 24886
rect 30380 24822 30432 24828
rect 30196 23860 30248 23866
rect 30196 23802 30248 23808
rect 30208 23730 30236 23802
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 30392 23186 30420 24822
rect 30484 24818 30512 25094
rect 30472 24812 30524 24818
rect 30472 24754 30524 24760
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30564 24132 30616 24138
rect 30564 24074 30616 24080
rect 30576 23866 30604 24074
rect 30564 23860 30616 23866
rect 30564 23802 30616 23808
rect 30472 23792 30524 23798
rect 30472 23734 30524 23740
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30196 23112 30248 23118
rect 30196 23054 30248 23060
rect 30208 22778 30236 23054
rect 30288 23044 30340 23050
rect 30288 22986 30340 22992
rect 30196 22772 30248 22778
rect 30196 22714 30248 22720
rect 30300 22710 30328 22986
rect 30288 22704 30340 22710
rect 30288 22646 30340 22652
rect 30392 22642 30420 23122
rect 30484 22778 30512 23734
rect 30668 23050 30696 24686
rect 30760 23118 30788 41386
rect 32416 35894 32444 47058
rect 34060 46640 34112 46646
rect 34060 46582 34112 46588
rect 32496 46504 32548 46510
rect 32496 46446 32548 46452
rect 33416 46504 33468 46510
rect 33416 46446 33468 46452
rect 32508 46170 32536 46446
rect 33428 46170 33456 46446
rect 32496 46164 32548 46170
rect 32496 46106 32548 46112
rect 33416 46164 33468 46170
rect 33416 46106 33468 46112
rect 32324 35866 32444 35894
rect 30932 35760 30984 35766
rect 30932 35702 30984 35708
rect 30944 35290 30972 35702
rect 31116 35488 31168 35494
rect 31116 35430 31168 35436
rect 30932 35284 30984 35290
rect 30932 35226 30984 35232
rect 31128 34066 31156 35430
rect 31852 34944 31904 34950
rect 31852 34886 31904 34892
rect 31116 34060 31168 34066
rect 31116 34002 31168 34008
rect 30840 33516 30892 33522
rect 30840 33458 30892 33464
rect 30852 33114 30880 33458
rect 30840 33108 30892 33114
rect 30840 33050 30892 33056
rect 31024 32224 31076 32230
rect 31024 32166 31076 32172
rect 31036 31226 31064 32166
rect 31128 31346 31156 34002
rect 31864 33930 31892 34886
rect 31392 33924 31444 33930
rect 31392 33866 31444 33872
rect 31852 33924 31904 33930
rect 31852 33866 31904 33872
rect 31300 33856 31352 33862
rect 31300 33798 31352 33804
rect 31312 33522 31340 33798
rect 31404 33658 31432 33866
rect 31392 33652 31444 33658
rect 31392 33594 31444 33600
rect 31300 33516 31352 33522
rect 31300 33458 31352 33464
rect 31312 32978 31340 33458
rect 31668 33448 31720 33454
rect 31668 33390 31720 33396
rect 31300 32972 31352 32978
rect 31300 32914 31352 32920
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 31220 32434 31248 32846
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 31220 31822 31248 32370
rect 31208 31816 31260 31822
rect 31208 31758 31260 31764
rect 31116 31340 31168 31346
rect 31116 31282 31168 31288
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31036 31198 31156 31226
rect 31128 30190 31156 31198
rect 31300 30660 31352 30666
rect 31300 30602 31352 30608
rect 31116 30184 31168 30190
rect 31116 30126 31168 30132
rect 30840 29844 30892 29850
rect 30840 29786 30892 29792
rect 31116 29844 31168 29850
rect 31116 29786 31168 29792
rect 30852 29628 30880 29786
rect 31024 29640 31076 29646
rect 30852 29600 31024 29628
rect 30852 29510 30880 29600
rect 31024 29582 31076 29588
rect 30840 29504 30892 29510
rect 30840 29446 30892 29452
rect 30932 29504 30984 29510
rect 31128 29458 31156 29786
rect 30932 29446 30984 29452
rect 30852 29170 30880 29446
rect 30840 29164 30892 29170
rect 30840 29106 30892 29112
rect 30944 27470 30972 29446
rect 31036 29430 31156 29458
rect 31036 29170 31064 29430
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 31036 28694 31064 29106
rect 31208 28960 31260 28966
rect 31208 28902 31260 28908
rect 31024 28688 31076 28694
rect 31024 28630 31076 28636
rect 31220 28626 31248 28902
rect 31208 28620 31260 28626
rect 31208 28562 31260 28568
rect 31220 27470 31248 28562
rect 31312 28150 31340 30602
rect 31404 30598 31432 31282
rect 31392 30592 31444 30598
rect 31392 30534 31444 30540
rect 31576 30048 31628 30054
rect 31576 29990 31628 29996
rect 31588 29714 31616 29990
rect 31392 29708 31444 29714
rect 31392 29650 31444 29656
rect 31576 29708 31628 29714
rect 31576 29650 31628 29656
rect 31404 29170 31432 29650
rect 31484 29504 31536 29510
rect 31484 29446 31536 29452
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31404 28558 31432 29106
rect 31392 28552 31444 28558
rect 31392 28494 31444 28500
rect 31300 28144 31352 28150
rect 31300 28086 31352 28092
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 31208 27464 31260 27470
rect 31208 27406 31260 27412
rect 31496 27402 31524 29446
rect 31576 29164 31628 29170
rect 31576 29106 31628 29112
rect 31588 28966 31616 29106
rect 31576 28960 31628 28966
rect 31576 28902 31628 28908
rect 31484 27396 31536 27402
rect 31484 27338 31536 27344
rect 31024 26988 31076 26994
rect 31024 26930 31076 26936
rect 30840 26784 30892 26790
rect 30840 26726 30892 26732
rect 30852 25906 30880 26726
rect 30932 26240 30984 26246
rect 30932 26182 30984 26188
rect 30944 25906 30972 26182
rect 30840 25900 30892 25906
rect 30840 25842 30892 25848
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 31036 25226 31064 26930
rect 31392 26240 31444 26246
rect 31392 26182 31444 26188
rect 31484 26240 31536 26246
rect 31484 26182 31536 26188
rect 31208 25900 31260 25906
rect 31208 25842 31260 25848
rect 31220 25498 31248 25842
rect 31300 25696 31352 25702
rect 31300 25638 31352 25644
rect 31208 25492 31260 25498
rect 31208 25434 31260 25440
rect 31116 25288 31168 25294
rect 31116 25230 31168 25236
rect 31024 25220 31076 25226
rect 31024 25162 31076 25168
rect 31036 24954 31064 25162
rect 31024 24948 31076 24954
rect 31024 24890 31076 24896
rect 31036 24274 31064 24890
rect 31128 24614 31156 25230
rect 31116 24608 31168 24614
rect 31116 24550 31168 24556
rect 31024 24268 31076 24274
rect 31024 24210 31076 24216
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 30944 23526 30972 23666
rect 30932 23520 30984 23526
rect 30932 23462 30984 23468
rect 31208 23520 31260 23526
rect 31208 23462 31260 23468
rect 30748 23112 30800 23118
rect 30748 23054 30800 23060
rect 30656 23044 30708 23050
rect 30656 22986 30708 22992
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 31036 22710 31064 22918
rect 31220 22710 31248 23462
rect 31024 22704 31076 22710
rect 31024 22646 31076 22652
rect 31208 22704 31260 22710
rect 31208 22646 31260 22652
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 31312 22094 31340 25638
rect 31404 25498 31432 26182
rect 31496 25974 31524 26182
rect 31484 25968 31536 25974
rect 31484 25910 31536 25916
rect 31484 25696 31536 25702
rect 31484 25638 31536 25644
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31496 25362 31524 25638
rect 31484 25356 31536 25362
rect 31484 25298 31536 25304
rect 31484 24812 31536 24818
rect 31484 24754 31536 24760
rect 31496 24410 31524 24754
rect 31484 24404 31536 24410
rect 31484 24346 31536 24352
rect 31312 22066 31432 22094
rect 31404 21162 31432 22066
rect 31128 21134 31432 21162
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 30380 19440 30432 19446
rect 30380 19382 30432 19388
rect 29828 18692 29880 18698
rect 29828 18634 29880 18640
rect 29840 18426 29868 18634
rect 29828 18420 29880 18426
rect 29828 18362 29880 18368
rect 30392 18358 30420 19382
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30484 18834 30512 19246
rect 30472 18828 30524 18834
rect 30472 18770 30524 18776
rect 30380 18352 30432 18358
rect 30380 18294 30432 18300
rect 30576 14414 30604 20878
rect 30656 20800 30708 20806
rect 30656 20742 30708 20748
rect 30668 19922 30696 20742
rect 30656 19916 30708 19922
rect 30656 19858 30708 19864
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30760 17746 30788 18022
rect 30748 17740 30800 17746
rect 30748 17682 30800 17688
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30472 13456 30524 13462
rect 30472 13398 30524 13404
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 28448 6180 28500 6186
rect 28448 6122 28500 6128
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 27068 2576 27120 2582
rect 27068 2518 27120 2524
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 26332 2304 26384 2310
rect 26332 2246 26384 2252
rect 26344 1970 26372 2246
rect 26332 1964 26384 1970
rect 26332 1906 26384 1912
rect 26436 800 26464 2314
rect 27080 800 27108 2314
rect 28368 800 28396 2314
rect 29656 800 29684 2382
rect 3054 776 3110 785
rect 3054 711 3110 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30484 762 30512 13398
rect 31128 2650 31156 21134
rect 31300 20256 31352 20262
rect 31300 20198 31352 20204
rect 31116 2644 31168 2650
rect 31116 2586 31168 2592
rect 31312 2378 31340 20198
rect 31680 4146 31708 33390
rect 31760 32224 31812 32230
rect 31760 32166 31812 32172
rect 31772 31822 31800 32166
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 32220 31748 32272 31754
rect 32220 31690 32272 31696
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 31772 27402 31800 28494
rect 32128 28076 32180 28082
rect 32128 28018 32180 28024
rect 32036 27940 32088 27946
rect 32036 27882 32088 27888
rect 31852 27872 31904 27878
rect 31852 27814 31904 27820
rect 31944 27872 31996 27878
rect 31944 27814 31996 27820
rect 31864 27674 31892 27814
rect 31852 27668 31904 27674
rect 31852 27610 31904 27616
rect 31956 27470 31984 27814
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 31760 27396 31812 27402
rect 31760 27338 31812 27344
rect 31772 27130 31800 27338
rect 31760 27124 31812 27130
rect 31760 27066 31812 27072
rect 31852 26920 31904 26926
rect 31852 26862 31904 26868
rect 31864 26382 31892 26862
rect 31944 26512 31996 26518
rect 31944 26454 31996 26460
rect 31852 26376 31904 26382
rect 31852 26318 31904 26324
rect 31864 25498 31892 26318
rect 31956 26042 31984 26454
rect 32048 26042 32076 27882
rect 32140 26450 32168 28018
rect 32232 27470 32260 31690
rect 32324 29050 32352 35866
rect 33508 34672 33560 34678
rect 33508 34614 33560 34620
rect 33520 33998 33548 34614
rect 33324 33992 33376 33998
rect 33508 33992 33560 33998
rect 33324 33934 33376 33940
rect 33428 33940 33508 33946
rect 33428 33934 33560 33940
rect 32404 33856 32456 33862
rect 32404 33798 32456 33804
rect 32416 33522 32444 33798
rect 33140 33652 33192 33658
rect 33140 33594 33192 33600
rect 32956 33584 33008 33590
rect 32956 33526 33008 33532
rect 32404 33516 32456 33522
rect 32404 33458 32456 33464
rect 32772 33516 32824 33522
rect 32772 33458 32824 33464
rect 32588 33312 32640 33318
rect 32588 33254 32640 33260
rect 32680 33312 32732 33318
rect 32680 33254 32732 33260
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32416 32366 32444 33050
rect 32600 32502 32628 33254
rect 32692 32910 32720 33254
rect 32784 33114 32812 33458
rect 32968 33454 32996 33526
rect 32956 33448 33008 33454
rect 32956 33390 33008 33396
rect 32772 33108 32824 33114
rect 32772 33050 32824 33056
rect 32968 32978 32996 33390
rect 33152 33046 33180 33594
rect 33336 33114 33364 33934
rect 33428 33918 33548 33934
rect 33428 33386 33456 33918
rect 33508 33856 33560 33862
rect 33508 33798 33560 33804
rect 33416 33380 33468 33386
rect 33416 33322 33468 33328
rect 33324 33108 33376 33114
rect 33324 33050 33376 33056
rect 33140 33040 33192 33046
rect 33140 32982 33192 32988
rect 33520 32978 33548 33798
rect 33692 33448 33744 33454
rect 33692 33390 33744 33396
rect 32956 32972 33008 32978
rect 32956 32914 33008 32920
rect 33508 32972 33560 32978
rect 33508 32914 33560 32920
rect 32680 32904 32732 32910
rect 32680 32846 32732 32852
rect 32588 32496 32640 32502
rect 32588 32438 32640 32444
rect 32404 32360 32456 32366
rect 32404 32302 32456 32308
rect 32588 32360 32640 32366
rect 32692 32348 32720 32846
rect 32968 32502 32996 32914
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33600 32904 33652 32910
rect 33600 32846 33652 32852
rect 33428 32570 33456 32846
rect 33416 32564 33468 32570
rect 33416 32506 33468 32512
rect 32956 32496 33008 32502
rect 32956 32438 33008 32444
rect 33232 32428 33284 32434
rect 33232 32370 33284 32376
rect 32640 32320 32720 32348
rect 32588 32302 32640 32308
rect 32600 31822 32628 32302
rect 32680 31884 32732 31890
rect 32680 31826 32732 31832
rect 32588 31816 32640 31822
rect 32588 31758 32640 31764
rect 32600 31482 32628 31758
rect 32588 31476 32640 31482
rect 32588 31418 32640 31424
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 32404 30116 32456 30122
rect 32404 30058 32456 30064
rect 32416 29646 32444 30058
rect 32508 29850 32536 30194
rect 32496 29844 32548 29850
rect 32496 29786 32548 29792
rect 32404 29640 32456 29646
rect 32404 29582 32456 29588
rect 32416 29510 32444 29582
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32588 29164 32640 29170
rect 32588 29106 32640 29112
rect 32324 29022 32444 29050
rect 32312 28960 32364 28966
rect 32312 28902 32364 28908
rect 32324 28694 32352 28902
rect 32312 28688 32364 28694
rect 32312 28630 32364 28636
rect 32416 27946 32444 29022
rect 32600 28762 32628 29106
rect 32588 28756 32640 28762
rect 32588 28698 32640 28704
rect 32496 28416 32548 28422
rect 32496 28358 32548 28364
rect 32508 28082 32536 28358
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 32404 27940 32456 27946
rect 32404 27882 32456 27888
rect 32220 27464 32272 27470
rect 32220 27406 32272 27412
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32312 27396 32364 27402
rect 32312 27338 32364 27344
rect 32128 26444 32180 26450
rect 32128 26386 32180 26392
rect 32324 26330 32352 27338
rect 32140 26302 32352 26330
rect 31944 26036 31996 26042
rect 31944 25978 31996 25984
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 31852 25492 31904 25498
rect 31852 25434 31904 25440
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31772 24750 31800 25298
rect 31852 25220 31904 25226
rect 31852 25162 31904 25168
rect 31760 24744 31812 24750
rect 31760 24686 31812 24692
rect 31772 24138 31800 24686
rect 31760 24132 31812 24138
rect 31760 24074 31812 24080
rect 31864 22778 31892 25162
rect 32048 23186 32076 25978
rect 32140 25770 32168 26302
rect 32128 25764 32180 25770
rect 32128 25706 32180 25712
rect 32220 25152 32272 25158
rect 32220 25094 32272 25100
rect 32232 24954 32260 25094
rect 32220 24948 32272 24954
rect 32220 24890 32272 24896
rect 32036 23180 32088 23186
rect 32036 23122 32088 23128
rect 31852 22772 31904 22778
rect 31852 22714 31904 22720
rect 32048 22642 32076 23122
rect 32036 22636 32088 22642
rect 32036 22578 32088 22584
rect 31760 22568 31812 22574
rect 31760 22510 31812 22516
rect 31772 21894 31800 22510
rect 31944 22432 31996 22438
rect 31944 22374 31996 22380
rect 31956 22030 31984 22374
rect 31944 22024 31996 22030
rect 31944 21966 31996 21972
rect 31760 21888 31812 21894
rect 31760 21830 31812 21836
rect 31760 20868 31812 20874
rect 31760 20810 31812 20816
rect 31772 19514 31800 20810
rect 32220 20528 32272 20534
rect 32220 20470 32272 20476
rect 32312 20528 32364 20534
rect 32312 20470 32364 20476
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 32232 12434 32260 20470
rect 32324 20398 32352 20470
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 32312 20256 32364 20262
rect 32312 20198 32364 20204
rect 32324 19378 32352 20198
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32416 18086 32444 18226
rect 32404 18080 32456 18086
rect 32404 18022 32456 18028
rect 32404 17604 32456 17610
rect 32404 17546 32456 17552
rect 32416 17338 32444 17546
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32140 12406 32260 12434
rect 32140 4486 32168 12406
rect 32508 7750 32536 27406
rect 32588 26376 32640 26382
rect 32588 26318 32640 26324
rect 32600 25362 32628 26318
rect 32588 25356 32640 25362
rect 32588 25298 32640 25304
rect 32588 20868 32640 20874
rect 32588 20810 32640 20816
rect 32600 20398 32628 20810
rect 32588 20392 32640 20398
rect 32588 20334 32640 20340
rect 32692 16574 32720 31826
rect 32772 31748 32824 31754
rect 32772 31690 32824 31696
rect 32784 27402 32812 31690
rect 32956 31680 33008 31686
rect 32956 31622 33008 31628
rect 32772 27396 32824 27402
rect 32772 27338 32824 27344
rect 32864 27056 32916 27062
rect 32864 26998 32916 27004
rect 32772 26852 32824 26858
rect 32772 26794 32824 26800
rect 32784 26382 32812 26794
rect 32876 26382 32904 26998
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 32864 25968 32916 25974
rect 32864 25910 32916 25916
rect 32772 25832 32824 25838
rect 32772 25774 32824 25780
rect 32784 25430 32812 25774
rect 32876 25498 32904 25910
rect 32864 25492 32916 25498
rect 32864 25434 32916 25440
rect 32772 25424 32824 25430
rect 32968 25378 32996 31622
rect 33140 31272 33192 31278
rect 33140 31214 33192 31220
rect 33152 30326 33180 31214
rect 33244 30734 33272 32370
rect 33612 32298 33640 32846
rect 33600 32292 33652 32298
rect 33600 32234 33652 32240
rect 33416 31952 33468 31958
rect 33416 31894 33468 31900
rect 33428 31278 33456 31894
rect 33612 31754 33640 32234
rect 33704 31890 33732 33390
rect 33876 32904 33928 32910
rect 33876 32846 33928 32852
rect 33692 31884 33744 31890
rect 33692 31826 33744 31832
rect 33520 31726 33640 31754
rect 33416 31272 33468 31278
rect 33416 31214 33468 31220
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33324 30592 33376 30598
rect 33324 30534 33376 30540
rect 33140 30320 33192 30326
rect 33140 30262 33192 30268
rect 33336 30258 33364 30534
rect 33520 30258 33548 31726
rect 33704 31414 33732 31826
rect 33692 31408 33744 31414
rect 33692 31350 33744 31356
rect 33692 30660 33744 30666
rect 33692 30602 33744 30608
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33232 30184 33284 30190
rect 33232 30126 33284 30132
rect 33600 30184 33652 30190
rect 33600 30126 33652 30132
rect 33244 29034 33272 30126
rect 33612 29850 33640 30126
rect 33600 29844 33652 29850
rect 33600 29786 33652 29792
rect 33704 29646 33732 30602
rect 33888 30258 33916 32846
rect 33876 30252 33928 30258
rect 33876 30194 33928 30200
rect 33416 29640 33468 29646
rect 33416 29582 33468 29588
rect 33692 29640 33744 29646
rect 33692 29582 33744 29588
rect 33232 29028 33284 29034
rect 33232 28970 33284 28976
rect 33428 28558 33456 29582
rect 33888 29170 33916 30194
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33980 29510 34008 29582
rect 33968 29504 34020 29510
rect 33968 29446 34020 29452
rect 33968 29300 34020 29306
rect 33968 29242 34020 29248
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 33692 29096 33744 29102
rect 33692 29038 33744 29044
rect 33508 29028 33560 29034
rect 33508 28970 33560 28976
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33324 27872 33376 27878
rect 33324 27814 33376 27820
rect 33336 27674 33364 27814
rect 33324 27668 33376 27674
rect 33324 27610 33376 27616
rect 33428 27538 33456 28494
rect 33416 27532 33468 27538
rect 33416 27474 33468 27480
rect 33048 26920 33100 26926
rect 33048 26862 33100 26868
rect 32772 25366 32824 25372
rect 32876 25350 32996 25378
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32784 23798 32812 25230
rect 32772 23792 32824 23798
rect 32772 23734 32824 23740
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 32784 23050 32812 23462
rect 32772 23044 32824 23050
rect 32772 22986 32824 22992
rect 32876 20874 32904 25350
rect 32956 24132 33008 24138
rect 32956 24074 33008 24080
rect 32968 23322 32996 24074
rect 32956 23316 33008 23322
rect 32956 23258 33008 23264
rect 32864 20868 32916 20874
rect 32864 20810 32916 20816
rect 32876 20602 32904 20810
rect 32864 20596 32916 20602
rect 32864 20538 32916 20544
rect 33060 19922 33088 26862
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33232 26308 33284 26314
rect 33232 26250 33284 26256
rect 33244 24342 33272 26250
rect 33336 25294 33364 26386
rect 33520 26382 33548 28970
rect 33600 28960 33652 28966
rect 33600 28902 33652 28908
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 33520 25294 33548 26318
rect 33324 25288 33376 25294
rect 33324 25230 33376 25236
rect 33508 25288 33560 25294
rect 33508 25230 33560 25236
rect 33232 24336 33284 24342
rect 33232 24278 33284 24284
rect 33416 23792 33468 23798
rect 33416 23734 33468 23740
rect 33428 23118 33456 23734
rect 33612 23594 33640 28902
rect 33704 28490 33732 29038
rect 33692 28484 33744 28490
rect 33692 28426 33744 28432
rect 33980 28218 34008 29242
rect 33968 28212 34020 28218
rect 33968 28154 34020 28160
rect 33980 26382 34008 28154
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 33876 25900 33928 25906
rect 33876 25842 33928 25848
rect 33784 25696 33836 25702
rect 33784 25638 33836 25644
rect 33796 25430 33824 25638
rect 33784 25424 33836 25430
rect 33784 25366 33836 25372
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33600 23588 33652 23594
rect 33600 23530 33652 23536
rect 33416 23112 33468 23118
rect 33416 23054 33468 23060
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33520 22642 33548 22918
rect 33508 22636 33560 22642
rect 33508 22578 33560 22584
rect 33048 19916 33100 19922
rect 33048 19858 33100 19864
rect 32692 16546 32812 16574
rect 32496 7744 32548 7750
rect 32496 7686 32548 7692
rect 32220 6248 32272 6254
rect 32220 6190 32272 6196
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 32140 4010 32168 4422
rect 32128 4004 32180 4010
rect 32128 3946 32180 3952
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 30760 870 30972 898
rect 30760 762 30788 870
rect 30944 800 30972 870
rect 32232 800 32260 6190
rect 32784 3942 32812 16546
rect 32772 3936 32824 3942
rect 32772 3878 32824 3884
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 32692 3534 32720 3674
rect 32680 3528 32732 3534
rect 32680 3470 32732 3476
rect 32784 3126 32812 3674
rect 33690 3632 33746 3641
rect 33690 3567 33692 3576
rect 33744 3567 33746 3576
rect 33692 3538 33744 3544
rect 32956 3528 33008 3534
rect 32954 3496 32956 3505
rect 33140 3528 33192 3534
rect 33008 3496 33010 3505
rect 33140 3470 33192 3476
rect 32954 3431 33010 3440
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 33060 3126 33088 3402
rect 32772 3120 32824 3126
rect 32772 3062 32824 3068
rect 33048 3120 33100 3126
rect 33048 3062 33100 3068
rect 33152 2990 33180 3470
rect 33140 2984 33192 2990
rect 33140 2926 33192 2932
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33520 800 33548 2926
rect 33796 2582 33824 25230
rect 33888 24818 33916 25842
rect 33980 25294 34008 26318
rect 33968 25288 34020 25294
rect 33968 25230 34020 25236
rect 33876 24812 33928 24818
rect 33876 24754 33928 24760
rect 34072 24342 34100 46582
rect 34152 26308 34204 26314
rect 34152 26250 34204 26256
rect 34164 24750 34192 26250
rect 34152 24744 34204 24750
rect 34152 24686 34204 24692
rect 34060 24336 34112 24342
rect 34060 24278 34112 24284
rect 33876 22024 33928 22030
rect 33876 21966 33928 21972
rect 33888 21690 33916 21966
rect 33876 21684 33928 21690
rect 33876 21626 33928 21632
rect 34256 21350 34284 47194
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35440 33584 35492 33590
rect 35440 33526 35492 33532
rect 34428 33448 34480 33454
rect 34428 33390 34480 33396
rect 34440 33114 34468 33390
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35452 33114 35480 33526
rect 34428 33108 34480 33114
rect 34428 33050 34480 33056
rect 35440 33108 35492 33114
rect 35440 33050 35492 33056
rect 34704 32904 34756 32910
rect 34704 32846 34756 32852
rect 34520 32292 34572 32298
rect 34520 32234 34572 32240
rect 34428 29708 34480 29714
rect 34428 29650 34480 29656
rect 34440 29578 34468 29650
rect 34428 29572 34480 29578
rect 34428 29514 34480 29520
rect 34440 29170 34468 29514
rect 34428 29164 34480 29170
rect 34428 29106 34480 29112
rect 34440 28626 34468 29106
rect 34428 28620 34480 28626
rect 34428 28562 34480 28568
rect 34532 28150 34560 32234
rect 34716 31822 34744 32846
rect 36176 32224 36228 32230
rect 36176 32166 36228 32172
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 36188 31890 36216 32166
rect 36176 31884 36228 31890
rect 36176 31826 36228 31832
rect 36636 31884 36688 31890
rect 36636 31826 36688 31832
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34796 31816 34848 31822
rect 34796 31758 34848 31764
rect 34716 31346 34744 31758
rect 34808 31414 34836 31758
rect 34796 31408 34848 31414
rect 34796 31350 34848 31356
rect 36648 31346 36676 31826
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 36176 31340 36228 31346
rect 36176 31282 36228 31288
rect 36636 31340 36688 31346
rect 36636 31282 36688 31288
rect 34612 29028 34664 29034
rect 34612 28970 34664 28976
rect 34624 28626 34652 28970
rect 34716 28642 34744 31282
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35348 30320 35400 30326
rect 35348 30262 35400 30268
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35360 29850 35388 30262
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 36084 29708 36136 29714
rect 36084 29650 36136 29656
rect 36096 29170 36124 29650
rect 36188 29646 36216 31282
rect 36268 30048 36320 30054
rect 36268 29990 36320 29996
rect 36176 29640 36228 29646
rect 36176 29582 36228 29588
rect 36280 29578 36308 29990
rect 36452 29844 36504 29850
rect 36452 29786 36504 29792
rect 36268 29572 36320 29578
rect 36268 29514 36320 29520
rect 36084 29164 36136 29170
rect 36084 29106 36136 29112
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 36096 28762 36124 29106
rect 36084 28756 36136 28762
rect 36084 28698 36136 28704
rect 34612 28620 34664 28626
rect 34716 28614 34836 28642
rect 34612 28562 34664 28568
rect 34704 28552 34756 28558
rect 34704 28494 34756 28500
rect 34520 28144 34572 28150
rect 34520 28086 34572 28092
rect 34428 28076 34480 28082
rect 34428 28018 34480 28024
rect 34336 27940 34388 27946
rect 34336 27882 34388 27888
rect 34348 22094 34376 27882
rect 34440 27878 34468 28018
rect 34428 27872 34480 27878
rect 34428 27814 34480 27820
rect 34440 23730 34468 27814
rect 34716 27538 34744 28494
rect 34808 28218 34836 28614
rect 36084 28484 36136 28490
rect 36084 28426 36136 28432
rect 36096 28218 36124 28426
rect 34796 28212 34848 28218
rect 34796 28154 34848 28160
rect 36084 28212 36136 28218
rect 36084 28154 36136 28160
rect 36084 27940 36136 27946
rect 36084 27882 36136 27888
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34704 27532 34756 27538
rect 34704 27474 34756 27480
rect 34716 25974 34744 27474
rect 36096 27470 36124 27882
rect 36464 27606 36492 29786
rect 36452 27600 36504 27606
rect 36452 27542 36504 27548
rect 36084 27464 36136 27470
rect 36084 27406 36136 27412
rect 36464 27130 36492 27542
rect 36452 27124 36504 27130
rect 36452 27066 36504 27072
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 36556 26042 36584 26182
rect 36544 26036 36596 26042
rect 36544 25978 36596 25984
rect 34704 25968 34756 25974
rect 34704 25910 34756 25916
rect 35348 25968 35400 25974
rect 35348 25910 35400 25916
rect 34612 25832 34664 25838
rect 34612 25774 34664 25780
rect 34624 25498 34652 25774
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35360 25498 35388 25910
rect 36084 25696 36136 25702
rect 36084 25638 36136 25644
rect 34612 25492 34664 25498
rect 34612 25434 34664 25440
rect 35348 25492 35400 25498
rect 35348 25434 35400 25440
rect 36096 25362 36124 25638
rect 36084 25356 36136 25362
rect 36084 25298 36136 25304
rect 34704 25288 34756 25294
rect 34704 25230 34756 25236
rect 34716 24206 34744 25230
rect 34796 24880 34848 24886
rect 34796 24822 34848 24828
rect 34808 24410 34836 24822
rect 35624 24608 35676 24614
rect 35624 24550 35676 24556
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34796 24404 34848 24410
rect 34796 24346 34848 24352
rect 35636 24274 35664 24550
rect 35624 24268 35676 24274
rect 35624 24210 35676 24216
rect 34704 24200 34756 24206
rect 34704 24142 34756 24148
rect 34716 23866 34744 24142
rect 37292 24070 37320 47382
rect 37648 47116 37700 47122
rect 37648 47058 37700 47064
rect 37660 32570 37688 47058
rect 38016 47048 38068 47054
rect 38016 46990 38068 46996
rect 38028 46578 38056 46990
rect 38016 46572 38068 46578
rect 38016 46514 38068 46520
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39764 47184 39816 47190
rect 39764 47126 39816 47132
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38200 46504 38252 46510
rect 38200 46446 38252 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38212 46170 38240 46446
rect 38200 46164 38252 46170
rect 38200 46106 38252 46112
rect 38108 45960 38160 45966
rect 38108 45902 38160 45908
rect 38120 38894 38148 45902
rect 38660 45416 38712 45422
rect 38660 45358 38712 45364
rect 38844 45416 38896 45422
rect 38844 45358 38896 45364
rect 38672 44742 38700 45358
rect 38856 45082 38884 45358
rect 38844 45076 38896 45082
rect 38844 45018 38896 45024
rect 38660 44736 38712 44742
rect 38660 44678 38712 44684
rect 38108 38888 38160 38894
rect 38108 38830 38160 38836
rect 37648 32564 37700 32570
rect 37648 32506 37700 32512
rect 37740 32360 37792 32366
rect 37740 32302 37792 32308
rect 37464 31748 37516 31754
rect 37464 31690 37516 31696
rect 37476 31482 37504 31690
rect 37556 31680 37608 31686
rect 37556 31622 37608 31628
rect 37464 31476 37516 31482
rect 37464 31418 37516 31424
rect 37568 31414 37596 31622
rect 37556 31408 37608 31414
rect 37556 31350 37608 31356
rect 37752 31278 37780 32302
rect 37740 31272 37792 31278
rect 37740 31214 37792 31220
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 34704 23860 34756 23866
rect 34704 23802 34756 23808
rect 34428 23724 34480 23730
rect 34428 23666 34480 23672
rect 38384 23724 38436 23730
rect 38384 23666 38436 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34348 22066 34468 22094
rect 34440 21622 34468 22066
rect 34520 21888 34572 21894
rect 34520 21830 34572 21836
rect 34532 21622 34560 21830
rect 34428 21616 34480 21622
rect 34428 21558 34480 21564
rect 34520 21616 34572 21622
rect 34520 21558 34572 21564
rect 35808 21412 35860 21418
rect 35808 21354 35860 21360
rect 34244 21344 34296 21350
rect 34244 21286 34296 21292
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35820 21078 35848 21354
rect 35900 21344 35952 21350
rect 35900 21286 35952 21292
rect 35808 21072 35860 21078
rect 35808 21014 35860 21020
rect 35912 20874 35940 21286
rect 35900 20868 35952 20874
rect 35900 20810 35952 20816
rect 36360 20868 36412 20874
rect 36360 20810 36412 20816
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 36174 4040 36230 4049
rect 36174 3975 36176 3984
rect 36228 3975 36230 3984
rect 36176 3946 36228 3952
rect 36268 3936 36320 3942
rect 36266 3904 36268 3913
rect 36320 3904 36322 3913
rect 34934 3836 35242 3856
rect 36266 3839 36322 3848
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33874 3632 33930 3641
rect 33874 3567 33876 3576
rect 33928 3567 33930 3576
rect 33876 3538 33928 3544
rect 33874 3496 33930 3505
rect 33874 3431 33876 3440
rect 33928 3431 33930 3440
rect 33876 3402 33928 3408
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35544 2650 35572 2790
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 33784 2576 33836 2582
rect 33784 2518 33836 2524
rect 35624 2508 35676 2514
rect 35624 2450 35676 2456
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 35636 2106 35664 2450
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 35624 2100 35676 2106
rect 35624 2042 35676 2048
rect 36096 800 36124 2314
rect 36188 1902 36216 2790
rect 36372 2514 36400 20810
rect 38396 16574 38424 23666
rect 39776 22778 39804 47126
rect 39960 45554 39988 49200
rect 41248 47410 41276 49200
rect 40512 47382 41276 47410
rect 40132 47048 40184 47054
rect 40132 46990 40184 46996
rect 40040 45892 40092 45898
rect 40040 45834 40092 45840
rect 39868 45526 39988 45554
rect 39868 45422 39896 45526
rect 39856 45416 39908 45422
rect 39856 45358 39908 45364
rect 40052 44878 40080 45834
rect 40040 44872 40092 44878
rect 40040 44814 40092 44820
rect 40052 24818 40080 44814
rect 40144 26450 40172 46990
rect 40316 44872 40368 44878
rect 40316 44814 40368 44820
rect 40328 37194 40356 44814
rect 40316 37188 40368 37194
rect 40316 37130 40368 37136
rect 40132 26444 40184 26450
rect 40132 26386 40184 26392
rect 40512 24857 40540 47382
rect 42260 46442 42288 49286
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49314 46470 50000
rect 46216 49286 46470 49314
rect 42248 46436 42300 46442
rect 42248 46378 42300 46384
rect 41052 46368 41104 46374
rect 41052 46310 41104 46316
rect 41064 46034 41092 46310
rect 42536 46034 42564 49200
rect 43180 47122 43208 49200
rect 43168 47116 43220 47122
rect 43168 47058 43220 47064
rect 42708 46980 42760 46986
rect 42708 46922 42760 46928
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 41052 46028 41104 46034
rect 41052 45970 41104 45976
rect 42524 46028 42576 46034
rect 42524 45970 42576 45976
rect 41236 45892 41288 45898
rect 41236 45834 41288 45840
rect 40684 45348 40736 45354
rect 40684 45290 40736 45296
rect 40696 44470 40724 45290
rect 41248 45082 41276 45834
rect 42628 45626 42656 46446
rect 42616 45620 42668 45626
rect 42616 45562 42668 45568
rect 42720 45558 42748 46922
rect 43824 45966 43852 49200
rect 44468 47410 44496 49200
rect 44192 47382 44496 47410
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 42708 45552 42760 45558
rect 42708 45494 42760 45500
rect 43996 45552 44048 45558
rect 43996 45494 44048 45500
rect 44008 45370 44036 45494
rect 44192 45490 44220 47382
rect 44456 45892 44508 45898
rect 44456 45834 44508 45840
rect 44180 45484 44232 45490
rect 44180 45426 44232 45432
rect 44008 45354 44312 45370
rect 42800 45348 42852 45354
rect 42800 45290 42852 45296
rect 44008 45348 44324 45354
rect 44008 45342 44272 45348
rect 41236 45076 41288 45082
rect 41236 45018 41288 45024
rect 40684 44464 40736 44470
rect 40684 44406 40736 44412
rect 40498 24848 40554 24857
rect 40040 24812 40092 24818
rect 40498 24783 40554 24792
rect 40040 24754 40092 24760
rect 40408 24608 40460 24614
rect 40408 24550 40460 24556
rect 40420 24274 40448 24550
rect 40408 24268 40460 24274
rect 40408 24210 40460 24216
rect 40224 24200 40276 24206
rect 40224 24142 40276 24148
rect 40236 23866 40264 24142
rect 40224 23860 40276 23866
rect 40224 23802 40276 23808
rect 40236 23186 40264 23802
rect 42812 23798 42840 45290
rect 44008 26382 44036 45342
rect 44272 45290 44324 45296
rect 44088 45280 44140 45286
rect 44088 45222 44140 45228
rect 43996 26376 44048 26382
rect 43996 26318 44048 26324
rect 44100 24954 44128 45222
rect 44272 44872 44324 44878
rect 44272 44814 44324 44820
rect 44284 38214 44312 44814
rect 44272 38208 44324 38214
rect 44272 38150 44324 38156
rect 44180 31272 44232 31278
rect 44180 31214 44232 31220
rect 44088 24948 44140 24954
rect 44088 24890 44140 24896
rect 43352 24200 43404 24206
rect 43352 24142 43404 24148
rect 43536 24200 43588 24206
rect 43536 24142 43588 24148
rect 43364 23866 43392 24142
rect 43352 23860 43404 23866
rect 43352 23802 43404 23808
rect 42800 23792 42852 23798
rect 42800 23734 42852 23740
rect 42616 23724 42668 23730
rect 42616 23666 42668 23672
rect 42628 23322 42656 23666
rect 42616 23316 42668 23322
rect 42616 23258 42668 23264
rect 42812 23254 42840 23734
rect 42800 23248 42852 23254
rect 42800 23190 42852 23196
rect 43364 23186 43392 23802
rect 40224 23180 40276 23186
rect 40224 23122 40276 23128
rect 41420 23180 41472 23186
rect 41420 23122 41472 23128
rect 43352 23180 43404 23186
rect 43352 23122 43404 23128
rect 40684 23112 40736 23118
rect 40684 23054 40736 23060
rect 40696 22778 40724 23054
rect 39764 22772 39816 22778
rect 39764 22714 39816 22720
rect 40684 22772 40736 22778
rect 40684 22714 40736 22720
rect 39776 22438 39804 22714
rect 40132 22636 40184 22642
rect 40132 22578 40184 22584
rect 39764 22432 39816 22438
rect 39764 22374 39816 22380
rect 40144 22030 40172 22578
rect 40316 22432 40368 22438
rect 40316 22374 40368 22380
rect 40328 22030 40356 22374
rect 40132 22024 40184 22030
rect 40132 21966 40184 21972
rect 40316 22024 40368 22030
rect 40316 21966 40368 21972
rect 40592 21956 40644 21962
rect 40592 21898 40644 21904
rect 40408 20392 40460 20398
rect 40408 20334 40460 20340
rect 40420 20058 40448 20334
rect 40408 20052 40460 20058
rect 40408 19994 40460 20000
rect 40500 18760 40552 18766
rect 40500 18702 40552 18708
rect 40512 18290 40540 18702
rect 40500 18284 40552 18290
rect 40500 18226 40552 18232
rect 38396 16546 38516 16574
rect 38488 5302 38516 16546
rect 40512 12434 40540 18226
rect 40420 12406 40540 12434
rect 40224 5704 40276 5710
rect 40224 5646 40276 5652
rect 40236 5370 40264 5646
rect 40316 5568 40368 5574
rect 40316 5510 40368 5516
rect 40224 5364 40276 5370
rect 40224 5306 40276 5312
rect 36544 5296 36596 5302
rect 36544 5238 36596 5244
rect 38476 5296 38528 5302
rect 38476 5238 38528 5244
rect 36556 4010 36584 5238
rect 38384 4276 38436 4282
rect 38384 4218 38436 4224
rect 37648 4208 37700 4214
rect 37648 4150 37700 4156
rect 36636 4140 36688 4146
rect 36636 4082 36688 4088
rect 36912 4140 36964 4146
rect 36912 4082 36964 4088
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 36544 3392 36596 3398
rect 36544 3334 36596 3340
rect 36556 2854 36584 3334
rect 36648 3194 36676 4082
rect 36924 4049 36952 4082
rect 36910 4040 36966 4049
rect 36910 3975 36966 3984
rect 37660 3194 37688 4150
rect 38396 4078 38424 4218
rect 38488 4214 38516 5238
rect 40328 5234 40356 5510
rect 40316 5228 40368 5234
rect 40316 5170 40368 5176
rect 40420 5114 40448 12406
rect 40328 5086 40448 5114
rect 39764 5024 39816 5030
rect 39764 4966 39816 4972
rect 39776 4690 39804 4966
rect 40224 4820 40276 4826
rect 40224 4762 40276 4768
rect 39764 4684 39816 4690
rect 39764 4626 39816 4632
rect 39488 4548 39540 4554
rect 39488 4490 39540 4496
rect 38476 4208 38528 4214
rect 38476 4150 38528 4156
rect 39500 4078 39528 4490
rect 38384 4072 38436 4078
rect 38384 4014 38436 4020
rect 39488 4072 39540 4078
rect 39488 4014 39540 4020
rect 39672 4072 39724 4078
rect 39672 4014 39724 4020
rect 39948 4072 40000 4078
rect 39948 4014 40000 4020
rect 39304 3664 39356 3670
rect 39304 3606 39356 3612
rect 37832 3528 37884 3534
rect 37832 3470 37884 3476
rect 36636 3188 36688 3194
rect 36636 3130 36688 3136
rect 37648 3188 37700 3194
rect 37648 3130 37700 3136
rect 37844 3058 37872 3470
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 38028 3126 38056 3334
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 39316 2990 39344 3606
rect 39500 2990 39528 4014
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 39488 2984 39540 2990
rect 39488 2926 39540 2932
rect 36544 2848 36596 2854
rect 36544 2790 36596 2796
rect 36360 2508 36412 2514
rect 36360 2450 36412 2456
rect 39684 2446 39712 4014
rect 39960 3534 39988 4014
rect 40132 3936 40184 3942
rect 40132 3878 40184 3884
rect 40144 3534 40172 3878
rect 40236 3602 40264 4762
rect 40224 3596 40276 3602
rect 40224 3538 40276 3544
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 39948 2508 40000 2514
rect 39948 2450 40000 2456
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 36176 1896 36228 1902
rect 36176 1838 36228 1844
rect 38028 800 38056 2314
rect 39316 800 39344 2314
rect 39960 800 39988 2450
rect 40328 1970 40356 5086
rect 40500 5024 40552 5030
rect 40500 4966 40552 4972
rect 40512 4690 40540 4966
rect 40500 4684 40552 4690
rect 40500 4626 40552 4632
rect 40604 4214 40632 21898
rect 40684 20324 40736 20330
rect 40684 20266 40736 20272
rect 40696 19922 40724 20266
rect 40684 19916 40736 19922
rect 40684 19858 40736 19864
rect 41144 19712 41196 19718
rect 41144 19654 41196 19660
rect 40684 18760 40736 18766
rect 40684 18702 40736 18708
rect 40696 18290 40724 18702
rect 41052 18624 41104 18630
rect 41052 18566 41104 18572
rect 40684 18284 40736 18290
rect 40684 18226 40736 18232
rect 40960 18284 41012 18290
rect 40960 18226 41012 18232
rect 40972 17542 41000 18226
rect 41064 18222 41092 18566
rect 41052 18216 41104 18222
rect 41052 18158 41104 18164
rect 41064 17814 41092 18158
rect 41052 17808 41104 17814
rect 41052 17750 41104 17756
rect 40960 17536 41012 17542
rect 40960 17478 41012 17484
rect 41156 16574 41184 19654
rect 41432 19446 41460 23122
rect 43076 23112 43128 23118
rect 43076 23054 43128 23060
rect 43088 22234 43116 23054
rect 43548 22982 43576 24142
rect 43812 24064 43864 24070
rect 43812 24006 43864 24012
rect 43824 23730 43852 24006
rect 43812 23724 43864 23730
rect 43812 23666 43864 23672
rect 43720 23656 43772 23662
rect 43720 23598 43772 23604
rect 43732 23118 43760 23598
rect 43720 23112 43772 23118
rect 43720 23054 43772 23060
rect 43536 22976 43588 22982
rect 43536 22918 43588 22924
rect 43076 22228 43128 22234
rect 43076 22170 43128 22176
rect 42892 22160 42944 22166
rect 42892 22102 42944 22108
rect 42904 21690 42932 22102
rect 43444 22024 43496 22030
rect 43444 21966 43496 21972
rect 43076 21956 43128 21962
rect 43076 21898 43128 21904
rect 42892 21684 42944 21690
rect 42892 21626 42944 21632
rect 43088 21622 43116 21898
rect 43352 21888 43404 21894
rect 43352 21830 43404 21836
rect 43076 21616 43128 21622
rect 42352 21554 42748 21570
rect 43076 21558 43128 21564
rect 42340 21548 42760 21554
rect 42392 21542 42708 21548
rect 42340 21490 42392 21496
rect 42708 21490 42760 21496
rect 41880 20392 41932 20398
rect 41880 20334 41932 20340
rect 41420 19440 41472 19446
rect 41420 19382 41472 19388
rect 41696 18760 41748 18766
rect 41696 18702 41748 18708
rect 41328 18080 41380 18086
rect 41328 18022 41380 18028
rect 41340 17882 41368 18022
rect 41328 17876 41380 17882
rect 41328 17818 41380 17824
rect 41708 17746 41736 18702
rect 41696 17740 41748 17746
rect 41696 17682 41748 17688
rect 41236 17536 41288 17542
rect 41236 17478 41288 17484
rect 41248 17134 41276 17478
rect 41788 17332 41840 17338
rect 41788 17274 41840 17280
rect 41236 17128 41288 17134
rect 41236 17070 41288 17076
rect 41156 16546 41276 16574
rect 41248 16114 41276 16546
rect 41236 16108 41288 16114
rect 41236 16050 41288 16056
rect 40776 5228 40828 5234
rect 40776 5170 40828 5176
rect 40960 5228 41012 5234
rect 40960 5170 41012 5176
rect 40788 4282 40816 5170
rect 40776 4276 40828 4282
rect 40776 4218 40828 4224
rect 40592 4208 40644 4214
rect 40592 4150 40644 4156
rect 40408 3936 40460 3942
rect 40408 3878 40460 3884
rect 40498 3904 40554 3913
rect 40420 3670 40448 3878
rect 40498 3839 40554 3848
rect 40512 3670 40540 3839
rect 40408 3664 40460 3670
rect 40408 3606 40460 3612
rect 40500 3664 40552 3670
rect 40500 3606 40552 3612
rect 40408 2984 40460 2990
rect 40408 2926 40460 2932
rect 40420 2446 40448 2926
rect 40604 2650 40632 4150
rect 40868 4140 40920 4146
rect 40868 4082 40920 4088
rect 40776 3528 40828 3534
rect 40776 3470 40828 3476
rect 40788 3194 40816 3470
rect 40880 3398 40908 4082
rect 40972 3738 41000 5170
rect 41248 4214 41276 16050
rect 41420 15904 41472 15910
rect 41420 15846 41472 15852
rect 41432 15570 41460 15846
rect 41420 15564 41472 15570
rect 41420 15506 41472 15512
rect 41236 4208 41288 4214
rect 41236 4150 41288 4156
rect 40960 3732 41012 3738
rect 40960 3674 41012 3680
rect 41420 3732 41472 3738
rect 41420 3674 41472 3680
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 40868 3392 40920 3398
rect 40868 3334 40920 3340
rect 41340 3194 41368 3402
rect 40776 3188 40828 3194
rect 40776 3130 40828 3136
rect 41328 3188 41380 3194
rect 41328 3130 41380 3136
rect 40592 2644 40644 2650
rect 40592 2586 40644 2592
rect 40776 2644 40828 2650
rect 40776 2586 40828 2592
rect 40408 2440 40460 2446
rect 40408 2382 40460 2388
rect 40592 2440 40644 2446
rect 40592 2382 40644 2388
rect 40316 1964 40368 1970
rect 40316 1906 40368 1912
rect 40604 800 40632 2382
rect 40684 2372 40736 2378
rect 40684 2314 40736 2320
rect 40696 2106 40724 2314
rect 40788 2310 40816 2586
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 40776 2304 40828 2310
rect 40776 2246 40828 2252
rect 40684 2100 40736 2106
rect 40684 2042 40736 2048
rect 41248 800 41276 2382
rect 41432 2378 41460 3674
rect 41604 3120 41656 3126
rect 41604 3062 41656 3068
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 41524 2650 41552 2994
rect 41512 2644 41564 2650
rect 41512 2586 41564 2592
rect 41616 2378 41644 3062
rect 41800 2394 41828 17274
rect 41892 2990 41920 20334
rect 42156 20052 42208 20058
rect 42156 19994 42208 20000
rect 42168 19446 42196 19994
rect 42248 19848 42300 19854
rect 42248 19790 42300 19796
rect 42260 19446 42288 19790
rect 42156 19440 42208 19446
rect 42156 19382 42208 19388
rect 42248 19440 42300 19446
rect 42248 19382 42300 19388
rect 42168 4690 42196 19382
rect 42260 17814 42288 19382
rect 42248 17808 42300 17814
rect 42248 17750 42300 17756
rect 42156 4684 42208 4690
rect 42156 4626 42208 4632
rect 42168 3602 42196 4626
rect 42156 3596 42208 3602
rect 42156 3538 42208 3544
rect 41880 2984 41932 2990
rect 41880 2926 41932 2932
rect 42352 2514 42380 21490
rect 43364 21418 43392 21830
rect 42800 21412 42852 21418
rect 42800 21354 42852 21360
rect 43352 21412 43404 21418
rect 43352 21354 43404 21360
rect 42812 20466 42840 21354
rect 43456 21010 43484 21966
rect 44192 21554 44220 31214
rect 44468 30122 44496 45834
rect 45112 45626 45140 49200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 45620 45152 45626
rect 45100 45562 45152 45568
rect 45100 45416 45152 45422
rect 45100 45358 45152 45364
rect 45112 45082 45140 45358
rect 45100 45076 45152 45082
rect 45100 45018 45152 45024
rect 45008 44872 45060 44878
rect 45008 44814 45060 44820
rect 44456 30116 44508 30122
rect 44456 30058 44508 30064
rect 44272 24812 44324 24818
rect 44272 24754 44324 24760
rect 44284 24138 44312 24754
rect 44272 24132 44324 24138
rect 44272 24074 44324 24080
rect 45020 23798 45048 44814
rect 45204 44402 45232 46990
rect 45468 46980 45520 46986
rect 45468 46922 45520 46928
rect 45376 46504 45428 46510
rect 45376 46446 45428 46452
rect 45388 45014 45416 46446
rect 45376 45008 45428 45014
rect 45376 44950 45428 44956
rect 45480 44538 45508 46922
rect 45652 46436 45704 46442
rect 45652 46378 45704 46384
rect 45560 45824 45612 45830
rect 45560 45766 45612 45772
rect 45468 44532 45520 44538
rect 45468 44474 45520 44480
rect 45192 44396 45244 44402
rect 45192 44338 45244 44344
rect 45572 36582 45600 45766
rect 45664 45554 45692 46378
rect 45756 45966 45784 49200
rect 45836 46096 45888 46102
rect 45836 46038 45888 46044
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45664 45526 45784 45554
rect 45756 44402 45784 45526
rect 45848 44742 45876 46038
rect 46216 45626 46244 49286
rect 46358 49200 46470 49286
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 46386 47016 46442 47025
rect 46386 46951 46442 46960
rect 46296 45960 46348 45966
rect 46296 45902 46348 45908
rect 46204 45620 46256 45626
rect 46204 45562 46256 45568
rect 45836 44736 45888 44742
rect 45836 44678 45888 44684
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45928 44328 45980 44334
rect 45928 44270 45980 44276
rect 45560 36576 45612 36582
rect 45560 36518 45612 36524
rect 45940 32502 45968 44270
rect 46308 43246 46336 45902
rect 46296 43240 46348 43246
rect 46296 43182 46348 43188
rect 46296 42696 46348 42702
rect 46296 42638 46348 42644
rect 46308 42226 46336 42638
rect 46296 42220 46348 42226
rect 46296 42162 46348 42168
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 46020 38956 46072 38962
rect 46020 38898 46072 38904
rect 45928 32496 45980 32502
rect 45928 32438 45980 32444
rect 46032 31090 46060 38898
rect 46112 33584 46164 33590
rect 46112 33526 46164 33532
rect 46124 31414 46152 33526
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46204 32360 46256 32366
rect 46204 32302 46256 32308
rect 46216 32065 46244 32302
rect 46202 32056 46258 32065
rect 46202 31991 46258 32000
rect 46308 31890 46336 32846
rect 46296 31884 46348 31890
rect 46296 31826 46348 31832
rect 46112 31408 46164 31414
rect 46112 31350 46164 31356
rect 45940 31062 46060 31090
rect 45834 28656 45890 28665
rect 45834 28591 45890 28600
rect 45652 28076 45704 28082
rect 45652 28018 45704 28024
rect 45664 27470 45692 28018
rect 45652 27464 45704 27470
rect 45652 27406 45704 27412
rect 45664 26994 45692 27406
rect 45744 27328 45796 27334
rect 45744 27270 45796 27276
rect 45652 26988 45704 26994
rect 45652 26930 45704 26936
rect 45664 26586 45692 26930
rect 45468 26580 45520 26586
rect 45468 26522 45520 26528
rect 45652 26580 45704 26586
rect 45652 26522 45704 26528
rect 45480 26382 45508 26522
rect 45664 26450 45692 26522
rect 45652 26444 45704 26450
rect 45652 26386 45704 26392
rect 45468 26376 45520 26382
rect 45468 26318 45520 26324
rect 45192 25832 45244 25838
rect 45192 25774 45244 25780
rect 45204 25430 45232 25774
rect 45192 25424 45244 25430
rect 45192 25366 45244 25372
rect 45480 25294 45508 26318
rect 45468 25288 45520 25294
rect 45468 25230 45520 25236
rect 45560 25152 45612 25158
rect 45560 25094 45612 25100
rect 45572 24834 45600 25094
rect 45100 24812 45152 24818
rect 45100 24754 45152 24760
rect 45480 24806 45600 24834
rect 45664 24818 45692 26386
rect 45756 25974 45784 27270
rect 45848 26042 45876 28591
rect 45836 26036 45888 26042
rect 45836 25978 45888 25984
rect 45940 25974 45968 31062
rect 46020 26376 46072 26382
rect 46020 26318 46072 26324
rect 45744 25968 45796 25974
rect 45744 25910 45796 25916
rect 45928 25968 45980 25974
rect 45928 25910 45980 25916
rect 45940 25378 45968 25910
rect 46032 25498 46060 26318
rect 46020 25492 46072 25498
rect 46020 25434 46072 25440
rect 45940 25350 46060 25378
rect 45928 25288 45980 25294
rect 45928 25230 45980 25236
rect 45652 24812 45704 24818
rect 45112 24138 45140 24754
rect 45480 24206 45508 24806
rect 45652 24754 45704 24760
rect 45652 24676 45704 24682
rect 45652 24618 45704 24624
rect 45468 24200 45520 24206
rect 45468 24142 45520 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 45100 24132 45152 24138
rect 45100 24074 45152 24080
rect 44364 23792 44416 23798
rect 44364 23734 44416 23740
rect 45008 23792 45060 23798
rect 45008 23734 45060 23740
rect 44376 23118 44404 23734
rect 45112 23338 45140 24074
rect 45376 23792 45428 23798
rect 45376 23734 45428 23740
rect 45020 23310 45140 23338
rect 44364 23112 44416 23118
rect 44364 23054 44416 23060
rect 44272 22500 44324 22506
rect 44272 22442 44324 22448
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 43536 21344 43588 21350
rect 43536 21286 43588 21292
rect 43444 21004 43496 21010
rect 43444 20946 43496 20952
rect 42800 20460 42852 20466
rect 42800 20402 42852 20408
rect 42616 20256 42668 20262
rect 42616 20198 42668 20204
rect 42628 19922 42656 20198
rect 42616 19916 42668 19922
rect 42616 19858 42668 19864
rect 42812 19378 42840 20402
rect 43076 20392 43128 20398
rect 43076 20334 43128 20340
rect 43088 19378 43116 20334
rect 43456 19990 43484 20946
rect 43548 20942 43576 21286
rect 44284 21078 44312 22442
rect 44272 21072 44324 21078
rect 44272 21014 44324 21020
rect 44088 21004 44140 21010
rect 44088 20946 44140 20952
rect 43536 20936 43588 20942
rect 43536 20878 43588 20884
rect 44100 20534 44128 20946
rect 44088 20528 44140 20534
rect 44088 20470 44140 20476
rect 43720 20460 43772 20466
rect 43720 20402 43772 20408
rect 43732 20058 43760 20402
rect 43812 20392 43864 20398
rect 43812 20334 43864 20340
rect 43720 20052 43772 20058
rect 43720 19994 43772 20000
rect 43444 19984 43496 19990
rect 43444 19926 43496 19932
rect 43260 19848 43312 19854
rect 43260 19790 43312 19796
rect 43444 19848 43496 19854
rect 43444 19790 43496 19796
rect 42800 19372 42852 19378
rect 42800 19314 42852 19320
rect 43076 19372 43128 19378
rect 43076 19314 43128 19320
rect 42708 18624 42760 18630
rect 42708 18566 42760 18572
rect 42720 18290 42748 18566
rect 42708 18284 42760 18290
rect 42708 18226 42760 18232
rect 42616 17536 42668 17542
rect 42616 17478 42668 17484
rect 42628 17202 42656 17478
rect 42616 17196 42668 17202
rect 42616 17138 42668 17144
rect 42984 17060 43036 17066
rect 42984 17002 43036 17008
rect 42996 16658 43024 17002
rect 42984 16652 43036 16658
rect 42984 16594 43036 16600
rect 42892 15564 42944 15570
rect 42892 15506 42944 15512
rect 42904 12434 42932 15506
rect 42812 12406 42932 12434
rect 42616 5568 42668 5574
rect 42616 5510 42668 5516
rect 42628 5302 42656 5510
rect 42616 5296 42668 5302
rect 42616 5238 42668 5244
rect 42812 3942 42840 12406
rect 42892 7336 42944 7342
rect 42892 7278 42944 7284
rect 42904 4690 42932 7278
rect 43088 6458 43116 19314
rect 43272 19310 43300 19790
rect 43456 19514 43484 19790
rect 43732 19786 43760 19994
rect 43720 19780 43772 19786
rect 43720 19722 43772 19728
rect 43824 19514 43852 20334
rect 43444 19508 43496 19514
rect 43444 19450 43496 19456
rect 43812 19508 43864 19514
rect 43812 19450 43864 19456
rect 44180 19440 44232 19446
rect 44180 19382 44232 19388
rect 43904 19372 43956 19378
rect 43904 19314 43956 19320
rect 44088 19372 44140 19378
rect 44088 19314 44140 19320
rect 43168 19304 43220 19310
rect 43168 19246 43220 19252
rect 43260 19304 43312 19310
rect 43260 19246 43312 19252
rect 43180 19174 43208 19246
rect 43168 19168 43220 19174
rect 43168 19110 43220 19116
rect 43272 18766 43300 19246
rect 43260 18760 43312 18766
rect 43260 18702 43312 18708
rect 43812 18760 43864 18766
rect 43812 18702 43864 18708
rect 43720 18692 43772 18698
rect 43720 18634 43772 18640
rect 43732 18290 43760 18634
rect 43720 18284 43772 18290
rect 43720 18226 43772 18232
rect 43444 18216 43496 18222
rect 43444 18158 43496 18164
rect 43456 15638 43484 18158
rect 43732 17746 43760 18226
rect 43720 17740 43772 17746
rect 43720 17682 43772 17688
rect 43824 17678 43852 18702
rect 43916 17882 43944 19314
rect 43996 19168 44048 19174
rect 43996 19110 44048 19116
rect 44008 18766 44036 19110
rect 43996 18760 44048 18766
rect 43996 18702 44048 18708
rect 43996 18216 44048 18222
rect 43996 18158 44048 18164
rect 43904 17876 43956 17882
rect 43904 17818 43956 17824
rect 43812 17672 43864 17678
rect 43812 17614 43864 17620
rect 44008 16658 44036 18158
rect 44100 18154 44128 19314
rect 44192 18766 44220 19382
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 44192 18426 44220 18702
rect 44180 18420 44232 18426
rect 44180 18362 44232 18368
rect 44192 18306 44220 18362
rect 44192 18278 44312 18306
rect 44180 18216 44232 18222
rect 44180 18158 44232 18164
rect 44088 18148 44140 18154
rect 44088 18090 44140 18096
rect 44192 17814 44220 18158
rect 44180 17808 44232 17814
rect 44180 17750 44232 17756
rect 44284 17678 44312 18278
rect 44272 17672 44324 17678
rect 44272 17614 44324 17620
rect 43996 16652 44048 16658
rect 43996 16594 44048 16600
rect 43444 15632 43496 15638
rect 43444 15574 43496 15580
rect 43076 6452 43128 6458
rect 43076 6394 43128 6400
rect 43536 5704 43588 5710
rect 43536 5646 43588 5652
rect 42892 4684 42944 4690
rect 42892 4626 42944 4632
rect 42904 4554 42932 4626
rect 42892 4548 42944 4554
rect 42892 4490 42944 4496
rect 43076 4548 43128 4554
rect 43076 4490 43128 4496
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 42984 3936 43036 3942
rect 42984 3878 43036 3884
rect 42996 3126 43024 3878
rect 43088 3534 43116 4490
rect 43548 3738 43576 5646
rect 43812 3936 43864 3942
rect 43812 3878 43864 3884
rect 43536 3732 43588 3738
rect 43536 3674 43588 3680
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 42984 3120 43036 3126
rect 42984 3062 43036 3068
rect 43088 2514 43116 3470
rect 43824 3194 43852 3878
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 43812 3188 43864 3194
rect 43812 3130 43864 3136
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 42340 2508 42392 2514
rect 42340 2450 42392 2456
rect 43076 2508 43128 2514
rect 43076 2450 43128 2456
rect 41420 2372 41472 2378
rect 41420 2314 41472 2320
rect 41604 2372 41656 2378
rect 41800 2366 42564 2394
rect 41604 2314 41656 2320
rect 42536 800 42564 2366
rect 43180 800 43208 2926
rect 44100 2922 44128 3334
rect 44088 2916 44140 2922
rect 44088 2858 44140 2864
rect 44284 2774 44312 17614
rect 44376 5302 44404 23054
rect 45020 22094 45048 23310
rect 45284 22636 45336 22642
rect 45284 22578 45336 22584
rect 45020 22066 45140 22094
rect 44640 21344 44692 21350
rect 44640 21286 44692 21292
rect 44652 20534 44680 21286
rect 44640 20528 44692 20534
rect 44640 20470 44692 20476
rect 45008 19712 45060 19718
rect 45008 19654 45060 19660
rect 45020 18766 45048 19654
rect 45008 18760 45060 18766
rect 45008 18702 45060 18708
rect 45020 17678 45048 18702
rect 45008 17672 45060 17678
rect 45008 17614 45060 17620
rect 44548 17060 44600 17066
rect 44548 17002 44600 17008
rect 44560 16590 44588 17002
rect 44548 16584 44600 16590
rect 44548 16526 44600 16532
rect 44364 5296 44416 5302
rect 44364 5238 44416 5244
rect 44376 4690 44404 5238
rect 44364 4684 44416 4690
rect 44364 4626 44416 4632
rect 44560 3534 44588 16526
rect 45112 13938 45140 22066
rect 45192 22024 45244 22030
rect 45192 21966 45244 21972
rect 45204 21554 45232 21966
rect 45296 21894 45324 22578
rect 45284 21888 45336 21894
rect 45284 21830 45336 21836
rect 45192 21548 45244 21554
rect 45192 21490 45244 21496
rect 45296 21418 45324 21830
rect 45284 21412 45336 21418
rect 45284 21354 45336 21360
rect 45388 20074 45416 23734
rect 45480 23730 45508 24142
rect 45572 23866 45600 24142
rect 45560 23860 45612 23866
rect 45560 23802 45612 23808
rect 45468 23724 45520 23730
rect 45468 23666 45520 23672
rect 45480 23118 45508 23666
rect 45468 23112 45520 23118
rect 45468 23054 45520 23060
rect 45572 22098 45600 23802
rect 45664 22778 45692 24618
rect 45836 23044 45888 23050
rect 45836 22986 45888 22992
rect 45652 22772 45704 22778
rect 45652 22714 45704 22720
rect 45664 22642 45692 22714
rect 45652 22636 45704 22642
rect 45652 22578 45704 22584
rect 45652 22432 45704 22438
rect 45652 22374 45704 22380
rect 45744 22432 45796 22438
rect 45744 22374 45796 22380
rect 45560 22092 45612 22098
rect 45560 22034 45612 22040
rect 45664 21962 45692 22374
rect 45652 21956 45704 21962
rect 45652 21898 45704 21904
rect 45468 21888 45520 21894
rect 45756 21842 45784 22374
rect 45468 21830 45520 21836
rect 45480 21350 45508 21830
rect 45572 21814 45784 21842
rect 45572 21622 45600 21814
rect 45560 21616 45612 21622
rect 45848 21570 45876 22986
rect 45560 21558 45612 21564
rect 45664 21542 45876 21570
rect 45468 21344 45520 21350
rect 45468 21286 45520 21292
rect 45388 20046 45508 20074
rect 45376 19304 45428 19310
rect 45376 19246 45428 19252
rect 45388 18970 45416 19246
rect 45376 18964 45428 18970
rect 45376 18906 45428 18912
rect 45284 18760 45336 18766
rect 45284 18702 45336 18708
rect 45296 17610 45324 18702
rect 45284 17604 45336 17610
rect 45284 17546 45336 17552
rect 45100 13932 45152 13938
rect 45100 13874 45152 13880
rect 45296 12434 45324 17546
rect 45480 17066 45508 20046
rect 45560 19848 45612 19854
rect 45560 19790 45612 19796
rect 45572 18465 45600 19790
rect 45558 18456 45614 18465
rect 45558 18391 45614 18400
rect 45664 18358 45692 21542
rect 45940 21434 45968 25230
rect 46032 24138 46060 25350
rect 46020 24132 46072 24138
rect 46020 24074 46072 24080
rect 46020 22568 46072 22574
rect 46020 22510 46072 22516
rect 46032 21690 46060 22510
rect 46020 21684 46072 21690
rect 46020 21626 46072 21632
rect 45756 21406 45968 21434
rect 45756 20602 45784 21406
rect 45836 21344 45888 21350
rect 45836 21286 45888 21292
rect 45848 20942 45876 21286
rect 45836 20936 45888 20942
rect 45836 20878 45888 20884
rect 45928 20800 45980 20806
rect 45928 20742 45980 20748
rect 45744 20596 45796 20602
rect 45744 20538 45796 20544
rect 45756 19922 45784 20538
rect 45836 20392 45888 20398
rect 45836 20334 45888 20340
rect 45848 19990 45876 20334
rect 45836 19984 45888 19990
rect 45836 19926 45888 19932
rect 45744 19916 45796 19922
rect 45744 19858 45796 19864
rect 45848 19310 45876 19926
rect 45940 19922 45968 20742
rect 45928 19916 45980 19922
rect 45928 19858 45980 19864
rect 45836 19304 45888 19310
rect 45836 19246 45888 19252
rect 45848 18358 45876 19246
rect 45652 18352 45704 18358
rect 45652 18294 45704 18300
rect 45836 18352 45888 18358
rect 45836 18294 45888 18300
rect 45468 17060 45520 17066
rect 45468 17002 45520 17008
rect 45468 16652 45520 16658
rect 45468 16594 45520 16600
rect 45296 12406 45416 12434
rect 45100 8492 45152 8498
rect 45100 8434 45152 8440
rect 45112 8090 45140 8434
rect 45284 8288 45336 8294
rect 45284 8230 45336 8236
rect 45100 8084 45152 8090
rect 45100 8026 45152 8032
rect 44824 7880 44876 7886
rect 44824 7822 44876 7828
rect 44836 7478 44864 7822
rect 45296 7818 45324 8230
rect 45388 7954 45416 12406
rect 45376 7948 45428 7954
rect 45376 7890 45428 7896
rect 45192 7812 45244 7818
rect 45192 7754 45244 7760
rect 45284 7812 45336 7818
rect 45284 7754 45336 7760
rect 45204 7546 45232 7754
rect 45192 7540 45244 7546
rect 45192 7482 45244 7488
rect 44824 7472 44876 7478
rect 44824 7414 44876 7420
rect 44836 4690 44864 7414
rect 45388 7342 45416 7890
rect 45376 7336 45428 7342
rect 45376 7278 45428 7284
rect 44824 4684 44876 4690
rect 44824 4626 44876 4632
rect 44548 3528 44600 3534
rect 44548 3470 44600 3476
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 45204 3058 45232 3470
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45480 2774 45508 16594
rect 45560 16448 45612 16454
rect 45560 16390 45612 16396
rect 45572 15745 45600 16390
rect 45558 15736 45614 15745
rect 45558 15671 45614 15680
rect 45664 10674 45692 18294
rect 45652 10668 45704 10674
rect 45652 10610 45704 10616
rect 46124 9450 46152 31350
rect 46400 26926 46428 46951
rect 47044 46646 47072 49200
rect 47688 47054 47716 49200
rect 48134 47696 48190 47705
rect 48134 47631 48190 47640
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47032 46640 47084 46646
rect 47032 46582 47084 46588
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47216 46368 47268 46374
rect 47964 46345 47992 46514
rect 47216 46310 47268 46316
rect 47950 46336 48006 46345
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46492 45082 46520 45834
rect 46480 45076 46532 45082
rect 46480 45018 46532 45024
rect 47032 44940 47084 44946
rect 47032 44882 47084 44888
rect 46756 44736 46808 44742
rect 46756 44678 46808 44684
rect 46572 44396 46624 44402
rect 46572 44338 46624 44344
rect 46480 32836 46532 32842
rect 46480 32778 46532 32784
rect 46492 32434 46520 32778
rect 46480 32428 46532 32434
rect 46480 32370 46532 32376
rect 46480 32224 46532 32230
rect 46480 32166 46532 32172
rect 46492 31890 46520 32166
rect 46480 31884 46532 31890
rect 46480 31826 46532 31832
rect 46584 27130 46612 44338
rect 46768 41138 46796 44678
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 46952 43858 46980 44134
rect 46940 43852 46992 43858
rect 46940 43794 46992 43800
rect 47044 43314 47072 44882
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 46940 41540 46992 41546
rect 46940 41482 46992 41488
rect 46952 41274 46980 41482
rect 46940 41268 46992 41274
rect 46940 41210 46992 41216
rect 46756 41132 46808 41138
rect 46756 41074 46808 41080
rect 46572 27124 46624 27130
rect 46572 27066 46624 27072
rect 46388 26920 46440 26926
rect 46388 26862 46440 26868
rect 46296 25696 46348 25702
rect 46296 25638 46348 25644
rect 46308 25362 46336 25638
rect 46296 25356 46348 25362
rect 46296 25298 46348 25304
rect 46388 24812 46440 24818
rect 46388 24754 46440 24760
rect 46204 24744 46256 24750
rect 46204 24686 46256 24692
rect 46216 23905 46244 24686
rect 46202 23896 46258 23905
rect 46202 23831 46258 23840
rect 46296 23656 46348 23662
rect 46296 23598 46348 23604
rect 46204 22568 46256 22574
rect 46202 22536 46204 22545
rect 46256 22536 46258 22545
rect 46202 22471 46258 22480
rect 46202 21856 46258 21865
rect 46202 21791 46258 21800
rect 46216 21554 46244 21791
rect 46204 21548 46256 21554
rect 46204 21490 46256 21496
rect 46308 20330 46336 23598
rect 46400 23225 46428 24754
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46480 24132 46532 24138
rect 46480 24074 46532 24080
rect 46386 23216 46442 23225
rect 46386 23151 46442 23160
rect 46296 20324 46348 20330
rect 46296 20266 46348 20272
rect 46492 19786 46520 24074
rect 46480 19780 46532 19786
rect 46480 19722 46532 19728
rect 46296 17672 46348 17678
rect 46296 17614 46348 17620
rect 46308 16794 46336 17614
rect 46388 17128 46440 17134
rect 46388 17070 46440 17076
rect 46296 16788 46348 16794
rect 46296 16730 46348 16736
rect 46400 16114 46428 17070
rect 46388 16108 46440 16114
rect 46388 16050 46440 16056
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 46308 12850 46336 13262
rect 46296 12844 46348 12850
rect 46296 12786 46348 12792
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46480 10464 46532 10470
rect 46480 10406 46532 10412
rect 46308 10130 46336 10406
rect 46492 10130 46520 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46480 10124 46532 10130
rect 46480 10066 46532 10072
rect 46112 9444 46164 9450
rect 46112 9386 46164 9392
rect 45560 8288 45612 8294
rect 45558 8256 45560 8265
rect 45612 8256 45614 8265
rect 45558 8191 45614 8200
rect 46584 4826 46612 27066
rect 46664 26784 46716 26790
rect 46664 26726 46716 26732
rect 46676 23254 46704 26726
rect 46664 23248 46716 23254
rect 46664 23190 46716 23196
rect 46768 20466 46796 41074
rect 46940 39364 46992 39370
rect 46940 39306 46992 39312
rect 46952 39098 46980 39306
rect 46940 39092 46992 39098
rect 46940 39034 46992 39040
rect 46940 38344 46992 38350
rect 46940 38286 46992 38292
rect 46952 37126 46980 38286
rect 46940 37120 46992 37126
rect 46940 37062 46992 37068
rect 47124 34944 47176 34950
rect 47124 34886 47176 34892
rect 47136 32978 47164 34886
rect 47124 32972 47176 32978
rect 47124 32914 47176 32920
rect 46846 31376 46902 31385
rect 46846 31311 46902 31320
rect 46860 30394 46888 31311
rect 46848 30388 46900 30394
rect 46848 30330 46900 30336
rect 46846 30016 46902 30025
rect 46846 29951 46902 29960
rect 46860 29782 46888 29951
rect 46848 29776 46900 29782
rect 46848 29718 46900 29724
rect 46940 28552 46992 28558
rect 46940 28494 46992 28500
rect 46952 27606 46980 28494
rect 46940 27600 46992 27606
rect 46940 27542 46992 27548
rect 46846 26616 46902 26625
rect 46846 26551 46902 26560
rect 46860 25838 46888 26551
rect 46848 25832 46900 25838
rect 46848 25774 46900 25780
rect 46940 22092 46992 22098
rect 46940 22034 46992 22040
rect 46756 20460 46808 20466
rect 46756 20402 46808 20408
rect 46952 20398 46980 22034
rect 46940 20392 46992 20398
rect 46940 20334 46992 20340
rect 46848 19236 46900 19242
rect 46848 19178 46900 19184
rect 46860 18290 46888 19178
rect 47228 18630 47256 46310
rect 47950 46271 48006 46280
rect 48148 46034 48176 47631
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 48136 46028 48188 46034
rect 48136 45970 48188 45976
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 47584 45348 47636 45354
rect 47584 45290 47636 45296
rect 47596 42226 47624 45290
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 47676 44804 47728 44810
rect 47676 44746 47728 44752
rect 47688 44538 47716 44746
rect 47676 44532 47728 44538
rect 47676 44474 47728 44480
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 47584 42220 47636 42226
rect 48134 42191 48190 42200
rect 47584 42162 47636 42168
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 40730 47716 41618
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 48044 41132 48096 41138
rect 48044 41074 48096 41080
rect 47952 40928 48004 40934
rect 48056 40905 48084 41074
rect 47952 40870 48004 40876
rect 48042 40896 48098 40905
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47676 38956 47728 38962
rect 47676 38898 47728 38904
rect 47688 38865 47716 38898
rect 47860 38888 47912 38894
rect 47674 38856 47730 38865
rect 47860 38830 47912 38836
rect 47674 38791 47730 38800
rect 47584 37868 47636 37874
rect 47584 37810 47636 37816
rect 47308 33312 47360 33318
rect 47308 33254 47360 33260
rect 47320 32842 47348 33254
rect 47400 32972 47452 32978
rect 47400 32914 47452 32920
rect 47308 32836 47360 32842
rect 47308 32778 47360 32784
rect 47412 31414 47440 32914
rect 47492 32428 47544 32434
rect 47492 32370 47544 32376
rect 47400 31408 47452 31414
rect 47400 31350 47452 31356
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47320 29345 47348 29582
rect 47306 29336 47362 29345
rect 47306 29271 47362 29280
rect 47400 28008 47452 28014
rect 47400 27950 47452 27956
rect 47308 26444 47360 26450
rect 47308 26386 47360 26392
rect 47216 18624 47268 18630
rect 47216 18566 47268 18572
rect 46848 18284 46900 18290
rect 46848 18226 46900 18232
rect 47216 18284 47268 18290
rect 47320 18272 47348 26386
rect 47412 24750 47440 27950
rect 47504 24818 47532 32370
rect 47596 28082 47624 37810
rect 47676 37664 47728 37670
rect 47676 37606 47728 37612
rect 47688 37194 47716 37606
rect 47676 37188 47728 37194
rect 47676 37130 47728 37136
rect 47872 35894 47900 38830
rect 47688 35866 47900 35894
rect 47964 35894 47992 40870
rect 48042 40831 48098 40840
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48226 39536 48282 39545
rect 48136 39500 48188 39506
rect 48226 39471 48282 39480
rect 48136 39442 48188 39448
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48148 37330 48176 38111
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 47964 35866 48084 35894
rect 47584 28076 47636 28082
rect 47584 28018 47636 28024
rect 47688 27962 47716 35866
rect 47860 34400 47912 34406
rect 47860 34342 47912 34348
rect 47872 33318 47900 34342
rect 47952 33992 48004 33998
rect 47952 33934 48004 33940
rect 47964 33425 47992 33934
rect 47950 33416 48006 33425
rect 47950 33351 48006 33360
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 47768 29640 47820 29646
rect 47768 29582 47820 29588
rect 47596 27934 47716 27962
rect 47596 26518 47624 27934
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27538 47716 27814
rect 47676 27532 47728 27538
rect 47676 27474 47728 27480
rect 47584 26512 47636 26518
rect 47584 26454 47636 26460
rect 47676 26308 47728 26314
rect 47676 26250 47728 26256
rect 47688 24818 47716 26250
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47676 24812 47728 24818
rect 47676 24754 47728 24760
rect 47400 24744 47452 24750
rect 47400 24686 47452 24692
rect 47268 18244 47348 18272
rect 47216 18226 47268 18232
rect 46940 18080 46992 18086
rect 46940 18022 46992 18028
rect 46952 17746 46980 18022
rect 46940 17740 46992 17746
rect 46940 17682 46992 17688
rect 46848 17128 46900 17134
rect 46846 17096 46848 17105
rect 46900 17096 46902 17105
rect 46846 17031 46902 17040
rect 46940 13728 46992 13734
rect 46940 13670 46992 13676
rect 46952 13394 46980 13670
rect 46940 13388 46992 13394
rect 46940 13330 46992 13336
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10810 46980 11018
rect 46940 10804 46992 10810
rect 46940 10746 46992 10752
rect 46664 10668 46716 10674
rect 46664 10610 46716 10616
rect 46572 4820 46624 4826
rect 46572 4762 46624 4768
rect 46676 4622 46704 10610
rect 46664 4616 46716 4622
rect 46664 4558 46716 4564
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3602 46336 3878
rect 46492 3602 46520 4422
rect 46860 4185 46888 4558
rect 46846 4176 46902 4185
rect 46756 4140 46808 4146
rect 46846 4111 46902 4120
rect 46756 4082 46808 4088
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 44192 2746 44312 2774
rect 45112 2746 45508 2774
rect 44192 2582 44220 2746
rect 44180 2576 44232 2582
rect 44180 2518 44232 2524
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 45112 800 45140 2746
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 45468 2304 45520 2310
rect 45468 2246 45520 2252
rect 45480 2038 45508 2246
rect 45468 2032 45520 2038
rect 45468 1974 45520 1980
rect 46400 800 46428 2314
rect 30484 734 30788 762
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46768 105 46796 4082
rect 47228 4078 47256 18226
rect 47412 12434 47440 24686
rect 47676 23520 47728 23526
rect 47676 23462 47728 23468
rect 47688 23186 47716 23462
rect 47676 23180 47728 23186
rect 47676 23122 47728 23128
rect 47584 22772 47636 22778
rect 47584 22714 47636 22720
rect 47596 21554 47624 22714
rect 47780 22574 47808 29582
rect 47950 25936 48006 25945
rect 47950 25871 48006 25880
rect 47964 25362 47992 25871
rect 47952 25356 48004 25362
rect 47952 25298 48004 25304
rect 48056 23594 48084 35866
rect 48136 35080 48188 35086
rect 48136 35022 48188 35028
rect 48148 34785 48176 35022
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48148 34105 48176 34546
rect 48134 34096 48190 34105
rect 48134 34031 48190 34040
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48148 31890 48176 32671
rect 48136 31884 48188 31890
rect 48136 31826 48188 31832
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48136 26308 48188 26314
rect 48136 26250 48188 26256
rect 48148 25265 48176 26250
rect 48134 25256 48190 25265
rect 48134 25191 48190 25200
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48044 23588 48096 23594
rect 48044 23530 48096 23536
rect 48148 23186 48176 24511
rect 48240 24274 48268 39471
rect 48228 24268 48280 24274
rect 48228 24210 48280 24216
rect 48136 23180 48188 23186
rect 48136 23122 48188 23128
rect 47860 22636 47912 22642
rect 47860 22578 47912 22584
rect 48044 22636 48096 22642
rect 48044 22578 48096 22584
rect 47768 22568 47820 22574
rect 47768 22510 47820 22516
rect 47780 21894 47808 22510
rect 47768 21888 47820 21894
rect 47768 21830 47820 21836
rect 47584 21548 47636 21554
rect 47584 21490 47636 21496
rect 47872 21486 47900 22578
rect 48056 21554 48084 22578
rect 48044 21548 48096 21554
rect 48044 21490 48096 21496
rect 47860 21480 47912 21486
rect 47860 21422 47912 21428
rect 47676 20868 47728 20874
rect 47676 20810 47728 20816
rect 47688 20602 47716 20810
rect 47676 20596 47728 20602
rect 47676 20538 47728 20544
rect 47584 19236 47636 19242
rect 47584 19178 47636 19184
rect 47596 18970 47624 19178
rect 47584 18964 47636 18970
rect 47584 18906 47636 18912
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47688 18426 47716 18634
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47872 12434 47900 21422
rect 47952 19372 48004 19378
rect 47952 19314 48004 19320
rect 47964 18630 47992 19314
rect 48056 19310 48084 21490
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48044 19304 48096 19310
rect 48044 19246 48096 19252
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48044 18964 48096 18970
rect 48044 18906 48096 18912
rect 47952 18624 48004 18630
rect 47952 18566 48004 18572
rect 47412 12406 47624 12434
rect 47596 10674 47624 12406
rect 47688 12406 47900 12434
rect 47584 10668 47636 10674
rect 47584 10610 47636 10616
rect 47308 7880 47360 7886
rect 47308 7822 47360 7828
rect 47320 7585 47348 7822
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47216 4072 47268 4078
rect 47216 4014 47268 4020
rect 46940 3936 46992 3942
rect 46940 3878 46992 3884
rect 46952 3670 46980 3878
rect 46940 3664 46992 3670
rect 46940 3606 46992 3612
rect 47596 2854 47624 10610
rect 47688 7954 47716 12406
rect 47858 9616 47914 9625
rect 47858 9551 47860 9560
rect 47912 9551 47914 9560
rect 47860 9522 47912 9528
rect 47766 8936 47822 8945
rect 47766 8871 47768 8880
rect 47820 8871 47822 8880
rect 47768 8842 47820 8848
rect 47676 7948 47728 7954
rect 47676 7890 47728 7896
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 47964 6225 47992 6258
rect 47950 6216 48006 6225
rect 47950 6151 48006 6160
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 47768 4208 47820 4214
rect 47768 4150 47820 4156
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47584 2848 47636 2854
rect 47584 2790 47636 2796
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 47780 1465 47808 4150
rect 47872 3505 47900 5170
rect 47858 3496 47914 3505
rect 47858 3431 47914 3440
rect 48056 3194 48084 18906
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 48148 16425 48176 17546
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 48148 12345 48176 13194
rect 48134 12336 48190 12345
rect 48134 12271 48190 12280
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48134 6831 48190 6840
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 48320 3052 48372 3058
rect 48320 2994 48372 3000
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 47766 1456 47822 1465
rect 47766 1391 47822 1400
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48056 785 48084 2382
rect 48332 800 48360 2994
rect 48976 800 49004 3402
rect 48042 776 48098 785
rect 48042 711 48098 720
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1858 47640 1914 47696
rect 3514 46960 3570 47016
rect 1398 42880 1454 42936
rect 1398 40160 1454 40216
rect 1582 35400 1638 35456
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 32680 1638 32736
rect 1858 41520 1914 41576
rect 1398 23160 1454 23216
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 1398 17720 1454 17776
rect 1398 12280 1454 12336
rect 2962 46280 3018 46336
rect 2778 36760 2834 36816
rect 2962 32000 3018 32056
rect 3422 44920 3478 44976
rect 3330 39480 3386 39536
rect 2226 19080 2282 19136
rect 3330 28600 3386 28656
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 8206 46980 8262 47016
rect 8206 46960 8208 46980
rect 8208 46960 8260 46980
rect 8260 46960 8262 46980
rect 3606 43560 3662 43616
rect 3790 31320 3846 31376
rect 3974 19760 4030 19816
rect 2962 18400 3018 18456
rect 2778 16360 2834 16416
rect 2778 15000 2834 15056
rect 3514 17076 3516 17096
rect 3516 17076 3568 17096
rect 3568 17076 3570 17096
rect 3514 17040 3570 17076
rect 3422 10240 3478 10296
rect 3422 7520 3478 7576
rect 3974 13640 4030 13696
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4986 19896 5042 19952
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3698 6840 3754 6896
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3514 3440 3570 3496
rect 3422 1400 3478 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 13910 28484 13966 28520
rect 13910 28464 13912 28484
rect 13912 28464 13964 28484
rect 13964 28464 13966 28484
rect 15382 28500 15384 28520
rect 15384 28500 15436 28520
rect 15436 28500 15438 28520
rect 15382 28464 15438 28500
rect 17498 28464 17554 28520
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 22006 32136 22062 32192
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 21086 28600 21142 28656
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 18418 3612 18420 3632
rect 18420 3612 18472 3632
rect 18472 3612 18474 3632
rect 18418 3576 18474 3612
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 21454 27240 21510 27296
rect 21270 24812 21326 24848
rect 21270 24792 21272 24812
rect 21272 24792 21324 24812
rect 21324 24792 21326 24812
rect 22190 26988 22246 27024
rect 22190 26968 22192 26988
rect 22192 26968 22244 26988
rect 22244 26968 22246 26988
rect 22834 27276 22836 27296
rect 22836 27276 22888 27296
rect 22888 27276 22890 27296
rect 22834 27240 22890 27276
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 25226 32544 25282 32600
rect 24674 31864 24730 31920
rect 25778 32836 25834 32872
rect 25778 32816 25780 32836
rect 25780 32816 25832 32836
rect 25832 32816 25834 32836
rect 25870 27820 25872 27840
rect 25872 27820 25924 27840
rect 25924 27820 25926 27840
rect 25870 27784 25926 27820
rect 26606 28600 26662 28656
rect 27802 32816 27858 32872
rect 27066 32136 27122 32192
rect 26330 3576 26386 3632
rect 28078 31900 28080 31920
rect 28080 31900 28132 31920
rect 28132 31900 28134 31920
rect 28078 31864 28134 31900
rect 27986 27820 27988 27840
rect 27988 27820 28040 27840
rect 28040 27820 28042 27840
rect 27986 27784 28042 27820
rect 28814 32544 28870 32600
rect 28998 32444 29000 32464
rect 29000 32444 29052 32464
rect 29052 32444 29054 32464
rect 28998 32408 29054 32444
rect 28722 28600 28778 28656
rect 29642 32408 29698 32464
rect 27986 19896 28042 19952
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 3054 720 3110 776
rect 33690 3596 33746 3632
rect 33690 3576 33692 3596
rect 33692 3576 33744 3596
rect 33744 3576 33746 3596
rect 32954 3476 32956 3496
rect 32956 3476 33008 3496
rect 33008 3476 33010 3496
rect 32954 3440 33010 3476
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 36174 4004 36230 4040
rect 36174 3984 36176 4004
rect 36176 3984 36228 4004
rect 36228 3984 36230 4004
rect 36266 3884 36268 3904
rect 36268 3884 36320 3904
rect 36320 3884 36322 3904
rect 36266 3848 36322 3884
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 33874 3596 33930 3632
rect 33874 3576 33876 3596
rect 33876 3576 33928 3596
rect 33928 3576 33930 3596
rect 33874 3460 33930 3496
rect 33874 3440 33876 3460
rect 33876 3440 33928 3460
rect 33928 3440 33930 3460
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 40498 24792 40554 24848
rect 36910 3984 36966 4040
rect 40498 3848 40554 3904
rect 46386 46960 46442 47016
rect 46202 32000 46258 32056
rect 45834 28600 45890 28656
rect 45558 18400 45614 18456
rect 45558 15680 45614 15736
rect 48134 47640 48190 47696
rect 46202 23840 46258 23896
rect 46202 22516 46204 22536
rect 46204 22516 46256 22536
rect 46256 22516 46258 22536
rect 46202 22480 46258 22516
rect 46202 21800 46258 21856
rect 46386 23160 46442 23216
rect 45558 8236 45560 8256
rect 45560 8236 45612 8256
rect 45612 8236 45614 8256
rect 45558 8200 45614 8236
rect 46846 31320 46902 31376
rect 46846 29960 46902 30016
rect 46846 26560 46902 26616
rect 47950 46280 48006 46336
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 47674 38800 47730 38856
rect 47306 29280 47362 29336
rect 48042 40840 48098 40896
rect 48134 40160 48190 40216
rect 48226 39480 48282 39536
rect 48134 38120 48190 38176
rect 47950 33360 48006 33416
rect 46846 17076 46848 17096
rect 46848 17076 46900 17096
rect 46900 17076 46902 17096
rect 46846 17040 46902 17076
rect 46846 4120 46902 4176
rect 47950 25880 48006 25936
rect 48134 34720 48190 34776
rect 48134 34040 48190 34096
rect 48134 32680 48190 32736
rect 48134 27920 48190 27976
rect 48134 25200 48190 25256
rect 48134 24520 48190 24576
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 47306 7520 47362 7576
rect 47858 9580 47914 9616
rect 47858 9560 47860 9580
rect 47860 9560 47912 9580
rect 47912 9560 47914 9580
rect 47766 8900 47822 8936
rect 47766 8880 47768 8900
rect 47768 8880 47820 8900
rect 47820 8880 47822 8900
rect 47950 6160 48006 6216
rect 47858 3440 47914 3496
rect 48134 16360 48190 16416
rect 48134 12280 48190 12336
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 48134 6840 48190 6896
rect 47766 1400 47822 1456
rect 46754 40 46810 96
rect 48042 720 48098 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1853 47698 1919 47701
rect 0 47696 1919 47698
rect 0 47640 1858 47696
rect 1914 47640 1919 47696
rect 0 47638 1919 47640
rect 0 47548 800 47638
rect 1853 47635 1919 47638
rect 48129 47698 48195 47701
rect 49200 47698 50000 47788
rect 48129 47696 50000 47698
rect 48129 47640 48134 47696
rect 48190 47640 50000 47696
rect 48129 47638 50000 47640
rect 48129 47635 48195 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3509 47018 3575 47021
rect 0 47016 3575 47018
rect 0 46960 3514 47016
rect 3570 46960 3575 47016
rect 0 46958 3575 46960
rect 0 46868 800 46958
rect 3509 46955 3575 46958
rect 8201 47018 8267 47021
rect 22318 47018 22324 47020
rect 8201 47016 22324 47018
rect 8201 46960 8206 47016
rect 8262 46960 22324 47016
rect 8201 46958 22324 46960
rect 8201 46955 8267 46958
rect 22318 46956 22324 46958
rect 22388 46956 22394 47020
rect 46381 47018 46447 47021
rect 49200 47018 50000 47108
rect 46381 47016 50000 47018
rect 46381 46960 46386 47016
rect 46442 46960 50000 47016
rect 46381 46958 50000 46960
rect 46381 46955 46447 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2957 46338 3023 46341
rect 0 46336 3023 46338
rect 0 46280 2962 46336
rect 3018 46280 3023 46336
rect 0 46278 3023 46280
rect 0 46188 800 46278
rect 2957 46275 3023 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3417 44978 3483 44981
rect 0 44976 3483 44978
rect 0 44920 3422 44976
rect 3478 44920 3483 44976
rect 0 44918 3483 44920
rect 0 44828 800 44918
rect 3417 44915 3483 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3601 43618 3667 43621
rect 0 43616 3667 43618
rect 0 43560 3606 43616
rect 3662 43560 3667 43616
rect 0 43558 3667 43560
rect 0 43468 800 43558
rect 3601 43555 3667 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 48037 40898 48103 40901
rect 49200 40898 50000 40988
rect 48037 40896 50000 40898
rect 48037 40840 48042 40896
rect 48098 40840 50000 40896
rect 48037 40838 50000 40840
rect 48037 40835 48103 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1393 40218 1459 40221
rect 0 40216 1459 40218
rect 0 40160 1398 40216
rect 1454 40160 1459 40216
rect 0 40158 1459 40160
rect 0 40068 800 40158
rect 1393 40155 1459 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3325 39538 3391 39541
rect 0 39536 3391 39538
rect 0 39480 3330 39536
rect 3386 39480 3391 39536
rect 0 39478 3391 39480
rect 0 39388 800 39478
rect 3325 39475 3391 39478
rect 48221 39538 48287 39541
rect 49200 39538 50000 39628
rect 48221 39536 50000 39538
rect 48221 39480 48226 39536
rect 48282 39480 50000 39536
rect 48221 39478 50000 39480
rect 48221 39475 48287 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47669 38858 47735 38861
rect 49200 38858 50000 38948
rect 47669 38856 50000 38858
rect 47669 38800 47674 38856
rect 47730 38800 50000 38856
rect 47669 38798 50000 38800
rect 47669 38795 47735 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48129 34098 48195 34101
rect 49200 34098 50000 34188
rect 48129 34096 50000 34098
rect 48129 34040 48134 34096
rect 48190 34040 50000 34096
rect 48129 34038 50000 34040
rect 48129 34035 48195 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 47945 33418 48011 33421
rect 49200 33418 50000 33508
rect 47945 33416 50000 33418
rect 47945 33360 47950 33416
rect 48006 33360 50000 33416
rect 47945 33358 50000 33360
rect 47945 33355 48011 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 25773 32874 25839 32877
rect 27797 32874 27863 32877
rect 25773 32872 27863 32874
rect 0 32738 800 32828
rect 25773 32816 25778 32872
rect 25834 32816 27802 32872
rect 27858 32816 27863 32872
rect 25773 32814 27863 32816
rect 25773 32811 25839 32814
rect 27797 32811 27863 32814
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 25221 32602 25287 32605
rect 28809 32602 28875 32605
rect 25221 32600 28875 32602
rect 25221 32544 25226 32600
rect 25282 32544 28814 32600
rect 28870 32544 28875 32600
rect 49200 32588 50000 32678
rect 25221 32542 28875 32544
rect 25221 32539 25287 32542
rect 28809 32539 28875 32542
rect 28993 32466 29059 32469
rect 29637 32466 29703 32469
rect 28993 32464 29703 32466
rect 28993 32408 28998 32464
rect 29054 32408 29642 32464
rect 29698 32408 29703 32464
rect 28993 32406 29703 32408
rect 28993 32403 29059 32406
rect 29637 32403 29703 32406
rect 22001 32194 22067 32197
rect 27061 32194 27127 32197
rect 22001 32192 27127 32194
rect 0 32058 800 32148
rect 22001 32136 22006 32192
rect 22062 32136 27066 32192
rect 27122 32136 27127 32192
rect 22001 32134 27127 32136
rect 22001 32131 22067 32134
rect 27061 32131 27127 32134
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 2957 32058 3023 32061
rect 0 32056 3023 32058
rect 0 32000 2962 32056
rect 3018 32000 3023 32056
rect 0 31998 3023 32000
rect 0 31908 800 31998
rect 2957 31995 3023 31998
rect 46197 32058 46263 32061
rect 49200 32058 50000 32148
rect 46197 32056 50000 32058
rect 46197 32000 46202 32056
rect 46258 32000 50000 32056
rect 46197 31998 50000 32000
rect 46197 31995 46263 31998
rect 24669 31922 24735 31925
rect 28073 31922 28139 31925
rect 24669 31920 28139 31922
rect 24669 31864 24674 31920
rect 24730 31864 28078 31920
rect 28134 31864 28139 31920
rect 49200 31908 50000 31998
rect 24669 31862 28139 31864
rect 24669 31859 24735 31862
rect 28073 31859 28139 31862
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3785 31378 3851 31381
rect 0 31376 3851 31378
rect 0 31320 3790 31376
rect 3846 31320 3851 31376
rect 0 31318 3851 31320
rect 0 31228 800 31318
rect 3785 31315 3851 31318
rect 46841 31378 46907 31381
rect 49200 31378 50000 31468
rect 46841 31376 50000 31378
rect 46841 31320 46846 31376
rect 46902 31320 50000 31376
rect 46841 31318 50000 31320
rect 46841 31315 46907 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 46841 30018 46907 30021
rect 49200 30018 50000 30108
rect 46841 30016 50000 30018
rect 46841 29960 46846 30016
rect 46902 29960 50000 30016
rect 46841 29958 50000 29960
rect 46841 29955 46907 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47301 29338 47367 29341
rect 49200 29338 50000 29428
rect 47301 29336 50000 29338
rect 47301 29280 47306 29336
rect 47362 29280 50000 29336
rect 47301 29278 50000 29280
rect 47301 29275 47367 29278
rect 49200 29188 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3325 28658 3391 28661
rect 0 28656 3391 28658
rect 0 28600 3330 28656
rect 3386 28600 3391 28656
rect 0 28598 3391 28600
rect 0 28508 800 28598
rect 3325 28595 3391 28598
rect 21081 28658 21147 28661
rect 26601 28658 26667 28661
rect 28717 28658 28783 28661
rect 21081 28656 28783 28658
rect 21081 28600 21086 28656
rect 21142 28600 26606 28656
rect 26662 28600 28722 28656
rect 28778 28600 28783 28656
rect 21081 28598 28783 28600
rect 21081 28595 21147 28598
rect 26601 28595 26667 28598
rect 28717 28595 28783 28598
rect 45829 28658 45895 28661
rect 49200 28658 50000 28748
rect 45829 28656 50000 28658
rect 45829 28600 45834 28656
rect 45890 28600 50000 28656
rect 45829 28598 50000 28600
rect 45829 28595 45895 28598
rect 13905 28522 13971 28525
rect 15377 28522 15443 28525
rect 17493 28522 17559 28525
rect 13905 28520 17559 28522
rect 13905 28464 13910 28520
rect 13966 28464 15382 28520
rect 15438 28464 17498 28520
rect 17554 28464 17559 28520
rect 49200 28508 50000 28598
rect 13905 28462 17559 28464
rect 13905 28459 13971 28462
rect 15377 28459 15443 28462
rect 17493 28459 17559 28462
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 25865 27842 25931 27845
rect 27981 27842 28047 27845
rect 25865 27840 28047 27842
rect 25865 27784 25870 27840
rect 25926 27784 27986 27840
rect 28042 27784 28047 27840
rect 49200 27828 50000 27918
rect 25865 27782 28047 27784
rect 25865 27779 25931 27782
rect 27981 27779 28047 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 21449 27298 21515 27301
rect 22829 27298 22895 27301
rect 21449 27296 22895 27298
rect 21449 27240 21454 27296
rect 21510 27240 22834 27296
rect 22890 27240 22895 27296
rect 21449 27238 22895 27240
rect 21449 27235 21515 27238
rect 22829 27235 22895 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 22185 27026 22251 27029
rect 22318 27026 22324 27028
rect 22185 27024 22324 27026
rect 22185 26968 22190 27024
rect 22246 26968 22324 27024
rect 22185 26966 22324 26968
rect 22185 26963 22251 26966
rect 22318 26964 22324 26966
rect 22388 26964 22394 27028
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 46841 26618 46907 26621
rect 49200 26618 50000 26708
rect 46841 26616 50000 26618
rect 46841 26560 46846 26616
rect 46902 26560 50000 26616
rect 46841 26558 50000 26560
rect 46841 26555 46907 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 47945 25938 48011 25941
rect 49200 25938 50000 26028
rect 47945 25936 50000 25938
rect 47945 25880 47950 25936
rect 48006 25880 50000 25936
rect 47945 25878 50000 25880
rect 47945 25875 48011 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 48129 25258 48195 25261
rect 49200 25258 50000 25348
rect 48129 25256 50000 25258
rect 48129 25200 48134 25256
rect 48190 25200 50000 25256
rect 48129 25198 50000 25200
rect 48129 25195 48195 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 21265 24850 21331 24853
rect 40493 24850 40559 24853
rect 21265 24848 40559 24850
rect 21265 24792 21270 24848
rect 21326 24792 40498 24848
rect 40554 24792 40559 24848
rect 21265 24790 40559 24792
rect 21265 24787 21331 24790
rect 40493 24787 40559 24790
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46197 23898 46263 23901
rect 49200 23898 50000 23988
rect 46197 23896 50000 23898
rect 46197 23840 46202 23896
rect 46258 23840 50000 23896
rect 46197 23838 50000 23840
rect 46197 23835 46263 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23068 800 23158
rect 1393 23155 1459 23158
rect 46381 23218 46447 23221
rect 49200 23218 50000 23308
rect 46381 23216 50000 23218
rect 46381 23160 46386 23216
rect 46442 23160 50000 23216
rect 46381 23158 50000 23160
rect 46381 23155 46447 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46197 22538 46263 22541
rect 49200 22538 50000 22628
rect 46197 22536 50000 22538
rect 46197 22480 46202 22536
rect 46258 22480 50000 22536
rect 46197 22478 50000 22480
rect 46197 22475 46263 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 46197 21858 46263 21861
rect 49200 21858 50000 21948
rect 46197 21856 50000 21858
rect 46197 21800 46202 21856
rect 46258 21800 50000 21856
rect 46197 21798 50000 21800
rect 46197 21795 46263 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 4981 19954 5047 19957
rect 27981 19954 28047 19957
rect 4981 19952 28047 19954
rect 0 19818 800 19908
rect 4981 19896 4986 19952
rect 5042 19896 27986 19952
rect 28042 19896 28047 19952
rect 4981 19894 28047 19896
rect 4981 19891 5047 19894
rect 27981 19891 28047 19894
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19668 800 19758
rect 3969 19755 4035 19758
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 2957 18458 3023 18461
rect 0 18456 3023 18458
rect 0 18400 2962 18456
rect 3018 18400 3023 18456
rect 0 18398 3023 18400
rect 0 18308 800 18398
rect 2957 18395 3023 18398
rect 45553 18458 45619 18461
rect 49200 18458 50000 18548
rect 45553 18456 50000 18458
rect 45553 18400 45558 18456
rect 45614 18400 50000 18456
rect 45553 18398 50000 18400
rect 45553 18395 45619 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3509 17098 3575 17101
rect 0 17096 3575 17098
rect 0 17040 3514 17096
rect 3570 17040 3575 17096
rect 0 17038 3575 17040
rect 0 16948 800 17038
rect 3509 17035 3575 17038
rect 46841 17098 46907 17101
rect 49200 17098 50000 17188
rect 46841 17096 50000 17098
rect 46841 17040 46846 17096
rect 46902 17040 50000 17096
rect 46841 17038 50000 17040
rect 46841 17035 46907 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16268 800 16358
rect 2773 16355 2839 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3969 13698 4035 13701
rect 0 13696 4035 13698
rect 0 13640 3974 13696
rect 4030 13640 4035 13696
rect 0 13638 4035 13640
rect 0 13548 800 13638
rect 3969 13635 4035 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 3417 10298 3483 10301
rect 0 10296 3483 10298
rect 0 10240 3422 10296
rect 3478 10240 3483 10296
rect 0 10238 3483 10240
rect 0 10148 800 10238
rect 3417 10235 3483 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 47853 9618 47919 9621
rect 49200 9618 50000 9708
rect 47853 9616 50000 9618
rect 47853 9560 47858 9616
rect 47914 9560 50000 9616
rect 47853 9558 50000 9560
rect 47853 9555 47919 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 45553 8258 45619 8261
rect 49200 8258 50000 8348
rect 45553 8256 50000 8258
rect 45553 8200 45558 8256
rect 45614 8200 50000 8256
rect 45553 8198 50000 8200
rect 45553 8195 45619 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3417 7578 3483 7581
rect 0 7576 3483 7578
rect 0 7520 3422 7576
rect 3478 7520 3483 7576
rect 0 7518 3483 7520
rect 0 7428 800 7518
rect 3417 7515 3483 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3693 6898 3759 6901
rect 0 6896 3759 6898
rect 0 6840 3698 6896
rect 3754 6840 3759 6896
rect 0 6838 3759 6840
rect 0 6748 800 6838
rect 3693 6835 3759 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 47945 6218 48011 6221
rect 49200 6218 50000 6308
rect 47945 6216 50000 6218
rect 47945 6160 47950 6216
rect 48006 6160 50000 6216
rect 47945 6158 50000 6160
rect 47945 6155 48011 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 36169 4042 36235 4045
rect 36905 4042 36971 4045
rect 36169 4040 36971 4042
rect 36169 3984 36174 4040
rect 36230 3984 36910 4040
rect 36966 3984 36971 4040
rect 49200 4028 50000 4118
rect 36169 3982 36971 3984
rect 36169 3979 36235 3982
rect 36905 3979 36971 3982
rect 36261 3906 36327 3909
rect 40493 3906 40559 3909
rect 36261 3904 40559 3906
rect 36261 3848 36266 3904
rect 36322 3848 40498 3904
rect 40554 3848 40559 3904
rect 36261 3846 40559 3848
rect 36261 3843 36327 3846
rect 40493 3843 40559 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 18413 3634 18479 3637
rect 26325 3634 26391 3637
rect 18413 3632 26391 3634
rect 0 3498 800 3588
rect 18413 3576 18418 3632
rect 18474 3576 26330 3632
rect 26386 3576 26391 3632
rect 18413 3574 26391 3576
rect 18413 3571 18479 3574
rect 26325 3571 26391 3574
rect 33685 3634 33751 3637
rect 33869 3634 33935 3637
rect 33685 3632 33935 3634
rect 33685 3576 33690 3632
rect 33746 3576 33874 3632
rect 33930 3576 33935 3632
rect 33685 3574 33935 3576
rect 33685 3571 33751 3574
rect 33869 3571 33935 3574
rect 3509 3498 3575 3501
rect 0 3496 3575 3498
rect 0 3440 3514 3496
rect 3570 3440 3575 3496
rect 0 3438 3575 3440
rect 0 3348 800 3438
rect 3509 3435 3575 3438
rect 32949 3498 33015 3501
rect 33869 3498 33935 3501
rect 32949 3496 33935 3498
rect 32949 3440 32954 3496
rect 33010 3440 33874 3496
rect 33930 3440 33935 3496
rect 32949 3438 33935 3440
rect 32949 3435 33015 3438
rect 33869 3435 33935 3438
rect 47853 3498 47919 3501
rect 49200 3498 50000 3588
rect 47853 3496 50000 3498
rect 47853 3440 47858 3496
rect 47914 3440 50000 3496
rect 47853 3438 50000 3440
rect 47853 3435 47919 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2668 800 2908
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1308 800 1398
rect 3417 1395 3483 1398
rect 47761 1458 47827 1461
rect 49200 1458 50000 1548
rect 47761 1456 50000 1458
rect 47761 1400 47766 1456
rect 47822 1400 50000 1456
rect 47761 1398 50000 1400
rect 47761 1395 47827 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 3049 778 3115 781
rect 0 776 3115 778
rect 0 720 3054 776
rect 3110 720 3115 776
rect 0 718 3115 720
rect 0 628 800 718
rect 3049 715 3115 718
rect 48037 778 48103 781
rect 49200 778 50000 868
rect 48037 776 50000 778
rect 48037 720 48042 776
rect 48098 720 50000 776
rect 48037 718 50000 720
rect 48037 715 48103 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 22324 46956 22388 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 22324 26964 22388 27028
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 22323 47020 22389 47021
rect 22323 46956 22324 47020
rect 22388 46956 22389 47020
rect 22323 46955 22389 46956
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 22326 27029 22386 46955
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 22323 27028 22389 27029
rect 22323 26964 22324 27028
rect 22388 26964 22389 27028
rect 22323 26963 22389 26964
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 40020 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 43608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform -1 0 30728 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 27968 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 43792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 38640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1644511149
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_89
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_200
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1644511149
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_314
timestamp 1644511149
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1644511149
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_430
timestamp 1644511149
transform 1 0 40664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1644511149
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1644511149
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_452
timestamp 1644511149
transform 1 0 42688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_460
timestamp 1644511149
transform 1 0 43424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_60
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_176
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_191
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_258
timestamp 1644511149
transform 1 0 24840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_296
timestamp 1644511149
transform 1 0 28336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_308
timestamp 1644511149
transform 1 0 29440 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_320
timestamp 1644511149
transform 1 0 30544 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_366
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_420
timestamp 1644511149
transform 1 0 39744 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_424
timestamp 1644511149
transform 1 0 40112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1644511149
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_440
timestamp 1644511149
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_474
timestamp 1644511149
transform 1 0 44712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_18
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1644511149
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1644511149
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp 1644511149
transform 1 0 11960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_134
timestamp 1644511149
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1644511149
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1644511149
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1644511149
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_224
timestamp 1644511149
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_231
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_237
timestamp 1644511149
transform 1 0 22908 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_261
timestamp 1644511149
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1644511149
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1644511149
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_397
timestamp 1644511149
transform 1 0 37628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_407
timestamp 1644511149
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1644511149
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_427
timestamp 1644511149
transform 1 0 40388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_452
timestamp 1644511149
transform 1 0 42688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_462
timestamp 1644511149
transform 1 0 43608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_31
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_89
timestamp 1644511149
transform 1 0 9292 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_97
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_101
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1644511149
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_136
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1644511149
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_185
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1644511149
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_407
timestamp 1644511149
transform 1 0 38548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_415
timestamp 1644511149
transform 1 0 39284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_425
timestamp 1644511149
transform 1 0 40204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_434
timestamp 1644511149
transform 1 0 41032 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_446
timestamp 1644511149
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_458
timestamp 1644511149
transform 1 0 43240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_465
timestamp 1644511149
transform 1 0 43884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_477
timestamp 1644511149
transform 1 0 44988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_492
timestamp 1644511149
transform 1 0 46368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_92
timestamp 1644511149
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_104
timestamp 1644511149
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_116
timestamp 1644511149
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_128
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1644511149
transform 1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1644511149
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1644511149
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1644511149
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_261
timestamp 1644511149
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_285
timestamp 1644511149
transform 1 0 27324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp 1644511149
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1644511149
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_425
timestamp 1644511149
transform 1 0 40204 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_447
timestamp 1644511149
transform 1 0 42228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_466
timestamp 1644511149
transform 1 0 43976 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_474
timestamp 1644511149
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_189
timestamp 1644511149
transform 1 0 18492 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_194
timestamp 1644511149
transform 1 0 18952 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_206
timestamp 1644511149
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1644511149
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_410
timestamp 1644511149
transform 1 0 38824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_418
timestamp 1644511149
transform 1 0 39560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_422
timestamp 1644511149
transform 1 0 39928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_436
timestamp 1644511149
transform 1 0 41216 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_462
timestamp 1644511149
transform 1 0 43608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_466
timestamp 1644511149
transform 1 0 43976 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_478
timestamp 1644511149
transform 1 0 45080 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_490
timestamp 1644511149
transform 1 0 46184 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1644511149
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_428
timestamp 1644511149
transform 1 0 40480 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_440
timestamp 1644511149
transform 1 0 41584 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_448
timestamp 1644511149
transform 1 0 42320 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_454
timestamp 1644511149
transform 1 0 42872 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1644511149
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1644511149
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_486
timestamp 1644511149
transform 1 0 45816 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_498
timestamp 1644511149
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_461
timestamp 1644511149
transform 1 0 43516 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_464
timestamp 1644511149
transform 1 0 43792 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_472
timestamp 1644511149
transform 1 0 44528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_491
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_499
timestamp 1644511149
transform 1 0 47012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_479
timestamp 1644511149
transform 1 0 45172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_491
timestamp 1644511149
transform 1 0 46276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_505
timestamp 1644511149
transform 1 0 47564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1644511149
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_489
timestamp 1644511149
transform 1 0 46092 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_493
timestamp 1644511149
transform 1 0 46460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_172
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_183
timestamp 1644511149
transform 1 0 17940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_236
timestamp 1644511149
transform 1 0 22816 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_202
timestamp 1644511149
transform 1 0 19688 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_246
timestamp 1644511149
transform 1 0 23736 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_258
timestamp 1644511149
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1644511149
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1644511149
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1644511149
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_218
timestamp 1644511149
transform 1 0 21160 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_226
timestamp 1644511149
transform 1 0 21896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_190
timestamp 1644511149
transform 1 0 18584 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_202
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1644511149
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1644511149
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_246
timestamp 1644511149
transform 1 0 23736 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_258
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1644511149
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1644511149
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_500
timestamp 1644511149
transform 1 0 47104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1644511149
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_171
timestamp 1644511149
transform 1 0 16836 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1644511149
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1644511149
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_225
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1644511149
transform 1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1644511149
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_145
timestamp 1644511149
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_152
timestamp 1644511149
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1644511149
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_204
timestamp 1644511149
transform 1 0 19872 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_216
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_229
timestamp 1644511149
transform 1 0 22172 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_240
timestamp 1644511149
transform 1 0 23184 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_252
timestamp 1644511149
transform 1 0 24288 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_264
timestamp 1644511149
transform 1 0 25392 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_147
timestamp 1644511149
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_168
timestamp 1644511149
transform 1 0 16560 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_176
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_257
timestamp 1644511149
transform 1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1644511149
transform 1 0 13340 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1644511149
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_146
timestamp 1644511149
transform 1 0 14536 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_150
timestamp 1644511149
transform 1 0 14904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1644511149
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_210
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1644511149
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_232
timestamp 1644511149
transform 1 0 22448 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_236
timestamp 1644511149
transform 1 0 22816 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1644511149
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1644511149
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_435
timestamp 1644511149
transform 1 0 41124 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_439
timestamp 1644511149
transform 1 0 41492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1644511149
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_162
timestamp 1644511149
transform 1 0 16008 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_174
timestamp 1644511149
transform 1 0 17112 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_184
timestamp 1644511149
transform 1 0 18032 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_200
timestamp 1644511149
transform 1 0 19504 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_212
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_220
timestamp 1644511149
transform 1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1644511149
transform 1 0 21988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_239
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_262
timestamp 1644511149
transform 1 0 25208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_274
timestamp 1644511149
transform 1 0 26312 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_285
timestamp 1644511149
transform 1 0 27324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_297
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1644511149
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_472
timestamp 1644511149
transform 1 0 44528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_498
timestamp 1644511149
transform 1 0 46920 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_507
timestamp 1644511149
transform 1 0 47748 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_515
timestamp 1644511149
transform 1 0 48484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_143
timestamp 1644511149
transform 1 0 14260 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1644511149
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_155
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1644511149
transform 1 0 16928 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1644511149
transform 1 0 18032 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1644511149
transform 1 0 19136 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_204
timestamp 1644511149
transform 1 0 19872 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_211
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_233
timestamp 1644511149
transform 1 0 22540 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1644511149
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_265
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_303
timestamp 1644511149
transform 1 0 28980 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_315
timestamp 1644511149
transform 1 0 30084 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_327
timestamp 1644511149
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_456
timestamp 1644511149
transform 1 0 43056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_468
timestamp 1644511149
transform 1 0 44160 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_476
timestamp 1644511149
transform 1 0 44896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_14
timestamp 1644511149
transform 1 0 2392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1644511149
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_152
timestamp 1644511149
transform 1 0 15088 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_164
timestamp 1644511149
transform 1 0 16192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1644511149
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_223
timestamp 1644511149
transform 1 0 21620 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_235
timestamp 1644511149
transform 1 0 22724 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1644511149
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_256
timestamp 1644511149
transform 1 0 24656 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_268
timestamp 1644511149
transform 1 0 25760 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_280
timestamp 1644511149
transform 1 0 26864 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_286
timestamp 1644511149
transform 1 0 27416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_317
timestamp 1644511149
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_341
timestamp 1644511149
transform 1 0 32476 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_353
timestamp 1644511149
transform 1 0 33580 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1644511149
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_429
timestamp 1644511149
transform 1 0 40572 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_437
timestamp 1644511149
transform 1 0 41308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_451
timestamp 1644511149
transform 1 0 42596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_482
timestamp 1644511149
transform 1 0 45448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_490
timestamp 1644511149
transform 1 0 46184 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_36
timestamp 1644511149
transform 1 0 4416 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_48
timestamp 1644511149
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1644511149
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1644511149
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1644511149
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_174
timestamp 1644511149
transform 1 0 17112 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1644511149
transform 1 0 17848 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_186
timestamp 1644511149
transform 1 0 18216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1644511149
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_215
timestamp 1644511149
transform 1 0 20884 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1644511149
transform 1 0 22448 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_244
timestamp 1644511149
transform 1 0 23552 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_262
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1644511149
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_309
timestamp 1644511149
transform 1 0 29532 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_315
timestamp 1644511149
transform 1 0 30084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_340
timestamp 1644511149
transform 1 0 32384 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_352
timestamp 1644511149
transform 1 0 33488 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_364
timestamp 1644511149
transform 1 0 34592 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_376
timestamp 1644511149
transform 1 0 35696 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1644511149
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_425
timestamp 1644511149
transform 1 0 40204 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_430
timestamp 1644511149
transform 1 0 40664 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_436
timestamp 1644511149
transform 1 0 41216 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_462
timestamp 1644511149
transform 1 0 43608 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_487
timestamp 1644511149
transform 1 0 45908 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_495
timestamp 1644511149
transform 1 0 46644 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_161
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_175
timestamp 1644511149
transform 1 0 17204 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1644511149
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_214
timestamp 1644511149
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_239
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1644511149
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_283
timestamp 1644511149
transform 1 0 27140 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_296
timestamp 1644511149
transform 1 0 28336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_303
timestamp 1644511149
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_331
timestamp 1644511149
transform 1 0 31556 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_343
timestamp 1644511149
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_355
timestamp 1644511149
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_427
timestamp 1644511149
transform 1 0 40388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_431
timestamp 1644511149
transform 1 0 40756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_443
timestamp 1644511149
transform 1 0 41860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_452
timestamp 1644511149
transform 1 0 42688 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1644511149
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_480
timestamp 1644511149
transform 1 0 45264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1644511149
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_129
timestamp 1644511149
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_133
timestamp 1644511149
transform 1 0 13340 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1644511149
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_155
timestamp 1644511149
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_196
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1644511149
transform 1 0 22448 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_244
timestamp 1644511149
transform 1 0 23552 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_252
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_260
timestamp 1644511149
transform 1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_268
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_289
timestamp 1644511149
transform 1 0 27692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_297
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_304
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_308
timestamp 1644511149
transform 1 0 29440 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_330
timestamp 1644511149
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_352
timestamp 1644511149
transform 1 0 33488 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_364
timestamp 1644511149
transform 1 0 34592 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_376
timestamp 1644511149
transform 1 0 35696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1644511149
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_453
timestamp 1644511149
transform 1 0 42780 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_459
timestamp 1644511149
transform 1 0 43332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_466
timestamp 1644511149
transform 1 0 43976 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_478
timestamp 1644511149
transform 1 0 45080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1644511149
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1644511149
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1644511149
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_159
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_171
timestamp 1644511149
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_175
timestamp 1644511149
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_183
timestamp 1644511149
transform 1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_205
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1644511149
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1644511149
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_256
timestamp 1644511149
transform 1 0 24656 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_283
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_291
timestamp 1644511149
transform 1 0 27876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_317
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_340
timestamp 1644511149
transform 1 0 32384 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_352
timestamp 1644511149
transform 1 0 33488 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_425
timestamp 1644511149
transform 1 0 40204 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_429
timestamp 1644511149
transform 1 0 40572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_441
timestamp 1644511149
transform 1 0 41676 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_449
timestamp 1644511149
transform 1 0 42412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_462
timestamp 1644511149
transform 1 0 43608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_481
timestamp 1644511149
transform 1 0 45356 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_506
timestamp 1644511149
transform 1 0 47656 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_514
timestamp 1644511149
transform 1 0 48392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_121
timestamp 1644511149
transform 1 0 12236 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_131
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_155
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1644511149
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_203
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1644511149
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_232
timestamp 1644511149
transform 1 0 22448 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_239
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_251
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_255
timestamp 1644511149
transform 1 0 24564 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_260
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_272
timestamp 1644511149
transform 1 0 26128 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_284
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_325
timestamp 1644511149
transform 1 0 31004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_350
timestamp 1644511149
transform 1 0 33304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_354
timestamp 1644511149
transform 1 0 33672 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_366
timestamp 1644511149
transform 1 0 34776 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_378
timestamp 1644511149
transform 1 0 35880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1644511149
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1644511149
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_454
timestamp 1644511149
transform 1 0 42872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_471
timestamp 1644511149
transform 1 0 44436 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_106
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_118
timestamp 1644511149
transform 1 0 11960 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp 1644511149
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1644511149
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_152
timestamp 1644511149
transform 1 0 15088 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_164
timestamp 1644511149
transform 1 0 16192 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_170
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_176
timestamp 1644511149
transform 1 0 17296 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1644511149
transform 1 0 17664 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_212
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_224
timestamp 1644511149
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_279
timestamp 1644511149
transform 1 0 26772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_290
timestamp 1644511149
transform 1 0 27784 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1644511149
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_317
timestamp 1644511149
transform 1 0 30268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_323
timestamp 1644511149
transform 1 0 30820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_344
timestamp 1644511149
transform 1 0 32752 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_356
timestamp 1644511149
transform 1 0 33856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 1644511149
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_379
timestamp 1644511149
transform 1 0 35972 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_391
timestamp 1644511149
transform 1 0 37076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_415
timestamp 1644511149
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_453
timestamp 1644511149
transform 1 0 42780 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_480
timestamp 1644511149
transform 1 0 45264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1644511149
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_103
timestamp 1644511149
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_145
timestamp 1644511149
transform 1 0 14444 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_184
timestamp 1644511149
transform 1 0 18032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_188
timestamp 1644511149
transform 1 0 18400 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_192
timestamp 1644511149
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_204
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_212
timestamp 1644511149
transform 1 0 20608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1644511149
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_234
timestamp 1644511149
transform 1 0 22632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_259
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1644511149
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_306
timestamp 1644511149
transform 1 0 29256 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_318
timestamp 1644511149
transform 1 0 30360 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1644511149
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_357
timestamp 1644511149
transform 1 0 33948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_370
timestamp 1644511149
transform 1 0 35144 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_382
timestamp 1644511149
transform 1 0 36248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1644511149
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_452
timestamp 1644511149
transform 1 0 42688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_462
timestamp 1644511149
transform 1 0 43608 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_469
timestamp 1644511149
transform 1 0 44252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_476
timestamp 1644511149
transform 1 0 44896 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_486
timestamp 1644511149
transform 1 0 45816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_88
timestamp 1644511149
transform 1 0 9200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_95
timestamp 1644511149
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1644511149
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_132
timestamp 1644511149
transform 1 0 13248 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_164
timestamp 1644511149
transform 1 0 16192 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1644511149
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_217
timestamp 1644511149
transform 1 0 21068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_229
timestamp 1644511149
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_237
timestamp 1644511149
transform 1 0 22908 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1644511149
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_285
timestamp 1644511149
transform 1 0 27324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_291
timestamp 1644511149
transform 1 0 27876 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1644511149
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_336
timestamp 1644511149
transform 1 0 32016 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_348
timestamp 1644511149
transform 1 0 33120 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_368
timestamp 1644511149
transform 1 0 34960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_380
timestamp 1644511149
transform 1 0 36064 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_392
timestamp 1644511149
transform 1 0 37168 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_404
timestamp 1644511149
transform 1 0 38272 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_429
timestamp 1644511149
transform 1 0 40572 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_441
timestamp 1644511149
transform 1 0 41676 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_453
timestamp 1644511149
transform 1 0 42780 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_460
timestamp 1644511149
transform 1 0 43424 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1644511149
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_481
timestamp 1644511149
transform 1 0 45356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_506
timestamp 1644511149
transform 1 0 47656 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_514
timestamp 1644511149
transform 1 0 48392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_101
timestamp 1644511149
transform 1 0 10396 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_126
timestamp 1644511149
transform 1 0 12696 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_157
timestamp 1644511149
transform 1 0 15548 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1644511149
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_180
timestamp 1644511149
transform 1 0 17664 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_188
timestamp 1644511149
transform 1 0 18400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_198
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_210
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_246
timestamp 1644511149
transform 1 0 23736 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_271
timestamp 1644511149
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_284
timestamp 1644511149
transform 1 0 27232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_291
timestamp 1644511149
transform 1 0 27876 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_299
timestamp 1644511149
transform 1 0 28612 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_307
timestamp 1644511149
transform 1 0 29348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_321
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1644511149
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_357
timestamp 1644511149
transform 1 0 33948 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_369
timestamp 1644511149
transform 1 0 35052 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_381
timestamp 1644511149
transform 1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1644511149
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_423
timestamp 1644511149
transform 1 0 40020 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_431
timestamp 1644511149
transform 1 0 40756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_443
timestamp 1644511149
transform 1 0 41860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_477
timestamp 1644511149
transform 1 0 44988 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_486
timestamp 1644511149
transform 1 0 45816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1644511149
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_111
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_147
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_176
timestamp 1644511149
transform 1 0 17296 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_183
timestamp 1644511149
transform 1 0 17940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1644511149
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_239
timestamp 1644511149
transform 1 0 23092 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_259
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_280
timestamp 1644511149
transform 1 0 26864 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_291
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_299
timestamp 1644511149
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_315
timestamp 1644511149
transform 1 0 30084 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_323
timestamp 1644511149
transform 1 0 30820 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_347
timestamp 1644511149
transform 1 0 33028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_354
timestamp 1644511149
transform 1 0 33672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1644511149
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_427
timestamp 1644511149
transform 1 0 40388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_452
timestamp 1644511149
transform 1 0 42688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_464
timestamp 1644511149
transform 1 0 43792 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_471
timestamp 1644511149
transform 1 0 44436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_487
timestamp 1644511149
transform 1 0 45908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_31
timestamp 1644511149
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1644511149
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_87
timestamp 1644511149
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_99
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_119
timestamp 1644511149
transform 1 0 12052 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_131
timestamp 1644511149
transform 1 0 13156 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1644511149
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_180
timestamp 1644511149
transform 1 0 17664 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_184
timestamp 1644511149
transform 1 0 18032 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_201
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_207
timestamp 1644511149
transform 1 0 20148 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1644511149
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1644511149
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_228
timestamp 1644511149
transform 1 0 22080 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_240
timestamp 1644511149
transform 1 0 23184 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_252
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_264
timestamp 1644511149
transform 1 0 25392 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_298
timestamp 1644511149
transform 1 0 28520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_306
timestamp 1644511149
transform 1 0 29256 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_312
timestamp 1644511149
transform 1 0 29808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_321
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_346
timestamp 1644511149
transform 1 0 32936 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_354
timestamp 1644511149
transform 1 0 33672 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_360
timestamp 1644511149
transform 1 0 34224 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_372
timestamp 1644511149
transform 1 0 35328 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_384
timestamp 1644511149
transform 1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_421
timestamp 1644511149
transform 1 0 39836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_440
timestamp 1644511149
transform 1 0 41584 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_458
timestamp 1644511149
transform 1 0 43240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_469
timestamp 1644511149
transform 1 0 44252 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_475
timestamp 1644511149
transform 1 0 44804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_482
timestamp 1644511149
transform 1 0 45448 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_495
timestamp 1644511149
transform 1 0 46644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_101
timestamp 1644511149
transform 1 0 10396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1644511149
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_120
timestamp 1644511149
transform 1 0 12144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_129
timestamp 1644511149
transform 1 0 12972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_144
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_148
timestamp 1644511149
transform 1 0 14720 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_156
timestamp 1644511149
transform 1 0 15456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_164
timestamp 1644511149
transform 1 0 16192 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_200
timestamp 1644511149
transform 1 0 19504 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1644511149
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1644511149
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_261
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1644511149
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1644511149
transform 1 0 27048 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_294
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1644511149
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_318
timestamp 1644511149
transform 1 0 30360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1644511149
transform 1 0 31188 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1644511149
transform 1 0 33396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_368
timestamp 1644511149
transform 1 0 34960 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_380
timestamp 1644511149
transform 1 0 36064 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_392
timestamp 1644511149
transform 1 0 37168 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_404
timestamp 1644511149
transform 1 0 38272 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1644511149
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_446
timestamp 1644511149
transform 1 0 42136 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_458
timestamp 1644511149
transform 1 0 43240 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_462
timestamp 1644511149
transform 1 0 43608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_472
timestamp 1644511149
transform 1 0 44528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_487
timestamp 1644511149
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_102
timestamp 1644511149
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1644511149
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1644511149
transform 1 0 11960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_126
timestamp 1644511149
transform 1 0 12696 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_159
timestamp 1644511149
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_197
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_231
timestamp 1644511149
transform 1 0 22356 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_255
timestamp 1644511149
transform 1 0 24564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1644511149
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_300
timestamp 1644511149
transform 1 0 28704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_310
timestamp 1644511149
transform 1 0 29624 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_316
timestamp 1644511149
transform 1 0 30176 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_323
timestamp 1644511149
transform 1 0 30820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1644511149
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_355
timestamp 1644511149
transform 1 0 33764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_376
timestamp 1644511149
transform 1 0 35696 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1644511149
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_425
timestamp 1644511149
transform 1 0 40204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_469
timestamp 1644511149
transform 1 0 44252 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_474
timestamp 1644511149
transform 1 0 44712 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_481
timestamp 1644511149
transform 1 0 45356 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1644511149
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_115
timestamp 1644511149
transform 1 0 11684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_122
timestamp 1644511149
transform 1 0 12328 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1644511149
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1644511149
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_154
timestamp 1644511149
transform 1 0 15272 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_161
timestamp 1644511149
transform 1 0 15916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_173
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_227
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_263
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_279
timestamp 1644511149
transform 1 0 26772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_291
timestamp 1644511149
transform 1 0 27876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_299
timestamp 1644511149
transform 1 0 28612 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_317
timestamp 1644511149
transform 1 0 30268 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_330
timestamp 1644511149
transform 1 0 31464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_340
timestamp 1644511149
transform 1 0 32384 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_347
timestamp 1644511149
transform 1 0 33028 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_369
timestamp 1644511149
transform 1 0 35052 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_381
timestamp 1644511149
transform 1 0 36156 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_393
timestamp 1644511149
transform 1 0 37260 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_405
timestamp 1644511149
transform 1 0 38364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_417
timestamp 1644511149
transform 1 0 39468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_472
timestamp 1644511149
transform 1 0 44528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_485
timestamp 1644511149
transform 1 0 45724 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_510
timestamp 1644511149
transform 1 0 48024 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_97
timestamp 1644511149
transform 1 0 10028 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_101
timestamp 1644511149
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1644511149
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_117
timestamp 1644511149
transform 1 0 11868 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_129
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_135
timestamp 1644511149
transform 1 0 13524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_148
timestamp 1644511149
transform 1 0 14720 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_156
timestamp 1644511149
transform 1 0 15456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_177
timestamp 1644511149
transform 1 0 17388 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_187
timestamp 1644511149
transform 1 0 18308 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_194
timestamp 1644511149
transform 1 0 18952 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_206
timestamp 1644511149
transform 1 0 20056 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_215
timestamp 1644511149
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_233
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_239
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_252
timestamp 1644511149
transform 1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_263
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_267
timestamp 1644511149
transform 1 0 25668 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_290
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_294
timestamp 1644511149
transform 1 0 28152 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_302
timestamp 1644511149
transform 1 0 28888 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_312
timestamp 1644511149
transform 1 0 29808 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_320
timestamp 1644511149
transform 1 0 30544 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1644511149
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_357
timestamp 1644511149
transform 1 0 33948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_381
timestamp 1644511149
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1644511149
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1644511149
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_105
timestamp 1644511149
transform 1 0 10764 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_111
timestamp 1644511149
transform 1 0 11316 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_115
timestamp 1644511149
transform 1 0 11684 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_119
timestamp 1644511149
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_127
timestamp 1644511149
transform 1 0 12788 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1644511149
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_154
timestamp 1644511149
transform 1 0 15272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_178
timestamp 1644511149
transform 1 0 17480 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_185
timestamp 1644511149
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1644511149
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_219
timestamp 1644511149
transform 1 0 21252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_241
timestamp 1644511149
transform 1 0 23276 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_273
timestamp 1644511149
transform 1 0 26220 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_278
timestamp 1644511149
transform 1 0 26680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1644511149
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_313
timestamp 1644511149
transform 1 0 29900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_325
timestamp 1644511149
transform 1 0 31004 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_335
timestamp 1644511149
transform 1 0 31924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_346
timestamp 1644511149
transform 1 0 32936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_350
timestamp 1644511149
transform 1 0 33304 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_472
timestamp 1644511149
transform 1 0 44528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_481
timestamp 1644511149
transform 1 0 45356 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_486
timestamp 1644511149
transform 1 0 45816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_490
timestamp 1644511149
transform 1 0 46184 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1644511149
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_96
timestamp 1644511149
transform 1 0 9936 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_102
timestamp 1644511149
transform 1 0 10488 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1644511149
transform 1 0 10948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_133
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_141
timestamp 1644511149
transform 1 0 14076 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_148
timestamp 1644511149
transform 1 0 14720 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_158
timestamp 1644511149
transform 1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1644511149
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_175
timestamp 1644511149
transform 1 0 17204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_179
timestamp 1644511149
transform 1 0 17572 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_204
timestamp 1644511149
transform 1 0 19872 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_212
timestamp 1644511149
transform 1 0 20608 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_234
timestamp 1644511149
transform 1 0 22632 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_255
timestamp 1644511149
transform 1 0 24564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_267
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_271
timestamp 1644511149
transform 1 0 26036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_289
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_299
timestamp 1644511149
transform 1 0 28612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_312
timestamp 1644511149
transform 1 0 29808 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_316
timestamp 1644511149
transform 1 0 30176 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_320
timestamp 1644511149
transform 1 0 30544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_479
timestamp 1644511149
transform 1 0 45172 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_500
timestamp 1644511149
transform 1 0 47104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_508
timestamp 1644511149
transform 1 0 47840 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_89
timestamp 1644511149
transform 1 0 9292 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_111
timestamp 1644511149
transform 1 0 11316 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_122
timestamp 1644511149
transform 1 0 12328 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_130
timestamp 1644511149
transform 1 0 13064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_162
timestamp 1644511149
transform 1 0 16008 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_174
timestamp 1644511149
transform 1 0 17112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_182
timestamp 1644511149
transform 1 0 17848 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1644511149
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1644511149
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_261
timestamp 1644511149
transform 1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_272
timestamp 1644511149
transform 1 0 26128 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_280
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_286
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_294
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1644511149
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_314
timestamp 1644511149
transform 1 0 29992 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_323
timestamp 1644511149
transform 1 0 30820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_330
timestamp 1644511149
transform 1 0 31464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_334
timestamp 1644511149
transform 1 0 31832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_343
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1644511149
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_385
timestamp 1644511149
transform 1 0 36524 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_397
timestamp 1644511149
transform 1 0 37628 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_409
timestamp 1644511149
transform 1 0 38732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1644511149
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_483
timestamp 1644511149
transform 1 0 45540 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_487
timestamp 1644511149
transform 1 0 45908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_101
timestamp 1644511149
transform 1 0 10396 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_136
timestamp 1644511149
transform 1 0 13616 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_148
timestamp 1644511149
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_158
timestamp 1644511149
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1644511149
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_189
timestamp 1644511149
transform 1 0 18492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_201
timestamp 1644511149
transform 1 0 19596 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_209
timestamp 1644511149
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_231
timestamp 1644511149
transform 1 0 22356 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_239
timestamp 1644511149
transform 1 0 23092 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1644511149
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_255
timestamp 1644511149
transform 1 0 24564 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_260
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_264
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_269
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_289
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_295
timestamp 1644511149
transform 1 0 28244 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_300
timestamp 1644511149
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_307
timestamp 1644511149
transform 1 0 29348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_314
timestamp 1644511149
transform 1 0 29992 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_324
timestamp 1644511149
transform 1 0 30912 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_343
timestamp 1644511149
transform 1 0 32660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_351
timestamp 1644511149
transform 1 0 33396 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_358
timestamp 1644511149
transform 1 0 34040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_366
timestamp 1644511149
transform 1 0 34776 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_370
timestamp 1644511149
transform 1 0 35144 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_374
timestamp 1644511149
transform 1 0 35512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1644511149
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1644511149
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_96
timestamp 1644511149
transform 1 0 9936 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_104
timestamp 1644511149
transform 1 0 10672 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_112
timestamp 1644511149
transform 1 0 11408 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_124
timestamp 1644511149
transform 1 0 12512 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_148
timestamp 1644511149
transform 1 0 14720 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_159
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_167
timestamp 1644511149
transform 1 0 16468 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_179
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1644511149
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_218
timestamp 1644511149
transform 1 0 21160 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_229
timestamp 1644511149
transform 1 0 22172 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1644511149
transform 1 0 23092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_281
timestamp 1644511149
transform 1 0 26956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_298
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1644511149
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_315
timestamp 1644511149
transform 1 0 30084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_324
timestamp 1644511149
transform 1 0 30912 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_332
timestamp 1644511149
transform 1 0 31648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_339
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_353
timestamp 1644511149
transform 1 0 33580 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1644511149
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_386
timestamp 1644511149
transform 1 0 36616 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_398
timestamp 1644511149
transform 1 0 37720 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_410
timestamp 1644511149
transform 1 0 38824 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_418
timestamp 1644511149
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_507
timestamp 1644511149
transform 1 0 47748 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_515
timestamp 1644511149
transform 1 0 48484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1644511149
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_130
timestamp 1644511149
transform 1 0 13064 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_138
timestamp 1644511149
transform 1 0 13800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_142
timestamp 1644511149
transform 1 0 14168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_148
timestamp 1644511149
transform 1 0 14720 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_154
timestamp 1644511149
transform 1 0 15272 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1644511149
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_175
timestamp 1644511149
transform 1 0 17204 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_183
timestamp 1644511149
transform 1 0 17940 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_206
timestamp 1644511149
transform 1 0 20056 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1644511149
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_242
timestamp 1644511149
transform 1 0 23368 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_250
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_262
timestamp 1644511149
transform 1 0 25208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_285
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_309
timestamp 1644511149
transform 1 0 29532 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_322
timestamp 1644511149
transform 1 0 30728 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_345
timestamp 1644511149
transform 1 0 32844 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_358
timestamp 1644511149
transform 1 0 34040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1644511149
transform 1 0 34868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1644511149
transform 1 0 35972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_117
timestamp 1644511149
transform 1 0 11868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_125
timestamp 1644511149
transform 1 0 12604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1644511149
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_160
timestamp 1644511149
transform 1 0 15824 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_184
timestamp 1644511149
transform 1 0 18032 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_240
timestamp 1644511149
transform 1 0 23184 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_269
timestamp 1644511149
transform 1 0 25852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_278
timestamp 1644511149
transform 1 0 26680 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_282
timestamp 1644511149
transform 1 0 27048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_291
timestamp 1644511149
transform 1 0 27876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_297
timestamp 1644511149
transform 1 0 28428 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_319
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_328
timestamp 1644511149
transform 1 0 31280 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_336
timestamp 1644511149
transform 1 0 32016 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_343
timestamp 1644511149
transform 1 0 32660 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_349
timestamp 1644511149
transform 1 0 33212 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_372
timestamp 1644511149
transform 1 0 35328 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_384
timestamp 1644511149
transform 1 0 36432 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_396
timestamp 1644511149
transform 1 0 37536 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_408
timestamp 1644511149
transform 1 0 38640 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_133
timestamp 1644511149
transform 1 0 13340 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_144
timestamp 1644511149
transform 1 0 14352 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_151
timestamp 1644511149
transform 1 0 14996 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_157
timestamp 1644511149
transform 1 0 15548 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1644511149
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_213
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_260
timestamp 1644511149
transform 1 0 25024 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1644511149
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_311
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_359
timestamp 1644511149
transform 1 0 34132 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_383
timestamp 1644511149
transform 1 0 36340 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_118
timestamp 1644511149
transform 1 0 11960 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_131
timestamp 1644511149
transform 1 0 13156 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_148
timestamp 1644511149
transform 1 0 14720 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_155
timestamp 1644511149
transform 1 0 15364 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1644511149
transform 1 0 17664 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_239
timestamp 1644511149
transform 1 0 23092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_259
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_270
timestamp 1644511149
transform 1 0 25944 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1644511149
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1644511149
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_331
timestamp 1644511149
transform 1 0 31556 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_343
timestamp 1644511149
transform 1 0 32660 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1644511149
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_30
timestamp 1644511149
transform 1 0 3864 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_42
timestamp 1644511149
transform 1 0 4968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1644511149
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_96
timestamp 1644511149
transform 1 0 9936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_116
timestamp 1644511149
transform 1 0 11776 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_128
timestamp 1644511149
transform 1 0 12880 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_156
timestamp 1644511149
transform 1 0 15456 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1644511149
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_173
timestamp 1644511149
transform 1 0 17020 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_185
timestamp 1644511149
transform 1 0 18124 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_246
timestamp 1644511149
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_250
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1644511149
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_287
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_292
timestamp 1644511149
transform 1 0 27968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_304
timestamp 1644511149
transform 1 0 29072 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_312
timestamp 1644511149
transform 1 0 29808 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_320
timestamp 1644511149
transform 1 0 30544 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_345
timestamp 1644511149
transform 1 0 32844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_368
timestamp 1644511149
transform 1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_380
timestamp 1644511149
transform 1 0 36064 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_396
timestamp 1644511149
transform 1 0 37536 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_408
timestamp 1644511149
transform 1 0 38640 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_420
timestamp 1644511149
transform 1 0 39744 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_432
timestamp 1644511149
transform 1 0 40848 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_444
timestamp 1644511149
transform 1 0 41952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_500
timestamp 1644511149
transform 1 0 47104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_89
timestamp 1644511149
transform 1 0 9292 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_111
timestamp 1644511149
transform 1 0 11316 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_117
timestamp 1644511149
transform 1 0 11868 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_128
timestamp 1644511149
transform 1 0 12880 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_156
timestamp 1644511149
transform 1 0 15456 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_168
timestamp 1644511149
transform 1 0 16560 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_180
timestamp 1644511149
transform 1 0 17664 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_205
timestamp 1644511149
transform 1 0 19964 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_211
timestamp 1644511149
transform 1 0 20516 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_218
timestamp 1644511149
transform 1 0 21160 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_224
timestamp 1644511149
transform 1 0 21712 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_231
timestamp 1644511149
transform 1 0 22356 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_243
timestamp 1644511149
transform 1 0 23460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_262
timestamp 1644511149
transform 1 0 25208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_266
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_274
timestamp 1644511149
transform 1 0 26312 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_286
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_293
timestamp 1644511149
transform 1 0 28060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1644511149
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_336
timestamp 1644511149
transform 1 0 32016 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_348
timestamp 1644511149
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_368
timestamp 1644511149
transform 1 0 34960 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_376
timestamp 1644511149
transform 1 0 35696 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_398
timestamp 1644511149
transform 1 0 37720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_410
timestamp 1644511149
transform 1 0 38824 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1644511149
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_11
timestamp 1644511149
transform 1 0 2116 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_36
timestamp 1644511149
transform 1 0 4416 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_48
timestamp 1644511149
transform 1 0 5520 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_134
timestamp 1644511149
transform 1 0 13432 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_145
timestamp 1644511149
transform 1 0 14444 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_157
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1644511149
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1644511149
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_243
timestamp 1644511149
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_255
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_270
timestamp 1644511149
transform 1 0 25944 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1644511149
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_297
timestamp 1644511149
transform 1 0 28428 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_311
timestamp 1644511149
transform 1 0 29716 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_318
timestamp 1644511149
transform 1 0 30360 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_326
timestamp 1644511149
transform 1 0 31096 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_331
timestamp 1644511149
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_344
timestamp 1644511149
transform 1 0 32752 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_348
timestamp 1644511149
transform 1 0 33120 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_354
timestamp 1644511149
transform 1 0 33672 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_366
timestamp 1644511149
transform 1 0 34776 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_378
timestamp 1644511149
transform 1 0 35880 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 1644511149
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_402
timestamp 1644511149
transform 1 0 38088 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_414
timestamp 1644511149
transform 1 0 39192 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_426
timestamp 1644511149
transform 1 0 40296 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_438
timestamp 1644511149
transform 1 0 41400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1644511149
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_489
timestamp 1644511149
transform 1 0 46092 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1644511149
transform 1 0 4048 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1644511149
transform 1 0 5152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1644511149
transform 1 0 6256 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1644511149
transform 1 0 7360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_119
timestamp 1644511149
transform 1 0 12052 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_131
timestamp 1644511149
transform 1 0 13156 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_163
timestamp 1644511149
transform 1 0 16100 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_175
timestamp 1644511149
transform 1 0 17204 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_187
timestamp 1644511149
transform 1 0 18308 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_217
timestamp 1644511149
transform 1 0 21068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_225
timestamp 1644511149
transform 1 0 21804 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_238
timestamp 1644511149
transform 1 0 23000 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1644511149
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_263
timestamp 1644511149
transform 1 0 25300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_267
timestamp 1644511149
transform 1 0 25668 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_275
timestamp 1644511149
transform 1 0 26404 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_286
timestamp 1644511149
transform 1 0 27416 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_295
timestamp 1644511149
transform 1 0 28244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_299
timestamp 1644511149
transform 1 0 28612 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_313
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_319
timestamp 1644511149
transform 1 0 30452 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1644511149
transform 1 0 31188 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_339
timestamp 1644511149
transform 1 0 32292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_347
timestamp 1644511149
transform 1 0 33028 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1644511149
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_374
timestamp 1644511149
transform 1 0 35512 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_386
timestamp 1644511149
transform 1 0 36616 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_398
timestamp 1644511149
transform 1 0 37720 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_410
timestamp 1644511149
transform 1 0 38824 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_418
timestamp 1644511149
transform 1 0 39560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_495
timestamp 1644511149
transform 1 0 46644 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_23
timestamp 1644511149
transform 1 0 3220 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_35
timestamp 1644511149
transform 1 0 4324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1644511149
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_141
timestamp 1644511149
transform 1 0 14076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_163
timestamp 1644511149
transform 1 0 16100 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_267
timestamp 1644511149
transform 1 0 25668 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1644511149
transform 1 0 27416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_299
timestamp 1644511149
transform 1 0 28612 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_308
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_315
timestamp 1644511149
transform 1 0 30084 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_343
timestamp 1644511149
transform 1 0 32660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_352
timestamp 1644511149
transform 1 0 33488 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_358
timestamp 1644511149
transform 1 0 34040 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1644511149
transform 1 0 35972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_511
timestamp 1644511149
transform 1 0 48116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_515
timestamp 1644511149
transform 1 0 48484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_213
timestamp 1644511149
transform 1 0 20700 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_217
timestamp 1644511149
transform 1 0 21068 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_225
timestamp 1644511149
transform 1 0 21804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_235
timestamp 1644511149
transform 1 0 22724 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_242
timestamp 1644511149
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1644511149
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_283
timestamp 1644511149
transform 1 0 27140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_295
timestamp 1644511149
transform 1 0 28244 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_319
timestamp 1644511149
transform 1 0 30452 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_325
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_346
timestamp 1644511149
transform 1 0 32936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_353
timestamp 1644511149
transform 1 0 33580 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_361
timestamp 1644511149
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_507
timestamp 1644511149
transform 1 0 47748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_245
timestamp 1644511149
transform 1 0 23644 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_260
timestamp 1644511149
transform 1 0 25024 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_285
timestamp 1644511149
transform 1 0 27324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_297
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_303
timestamp 1644511149
transform 1 0 28980 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_311
timestamp 1644511149
transform 1 0 29716 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 1644511149
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1644511149
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_6
timestamp 1644511149
transform 1 0 1656 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_10
timestamp 1644511149
transform 1 0 2024 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_14
timestamp 1644511149
transform 1 0 2392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1644511149
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_238
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_258
timestamp 1644511149
transform 1 0 24840 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_266
timestamp 1644511149
transform 1 0 25576 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_276
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_318
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_334
timestamp 1644511149
transform 1 0 31832 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_346
timestamp 1644511149
transform 1 0 32936 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1644511149
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_11
timestamp 1644511149
transform 1 0 2116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_23
timestamp 1644511149
transform 1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_35
timestamp 1644511149
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 1644511149
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1644511149
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_252
timestamp 1644511149
transform 1 0 24288 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_287
timestamp 1644511149
transform 1 0 27508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_299
timestamp 1644511149
transform 1 0 28612 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_307
timestamp 1644511149
transform 1 0 29348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1644511149
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_241
timestamp 1644511149
transform 1 0 23276 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1644511149
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_270
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_274
timestamp 1644511149
transform 1 0 26312 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_282
timestamp 1644511149
transform 1 0 27048 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_294
timestamp 1644511149
transform 1 0 28152 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1644511149
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_269
timestamp 1644511149
transform 1 0 25852 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_290
timestamp 1644511149
transform 1 0 27784 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_294
timestamp 1644511149
transform 1 0 28152 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1644511149
transform 1 0 29256 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1644511149
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_271
timestamp 1644511149
transform 1 0 26036 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_283
timestamp 1644511149
transform 1 0 27140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_295
timestamp 1644511149
transform 1 0 28244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_271
timestamp 1644511149
transform 1 0 26036 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_292
timestamp 1644511149
transform 1 0 27968 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_507
timestamp 1644511149
transform 1 0 47748 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_515
timestamp 1644511149
transform 1 0 48484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_269
timestamp 1644511149
transform 1 0 25852 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_274
timestamp 1644511149
transform 1 0 26312 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1644511149
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_14
timestamp 1644511149
transform 1 0 2392 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_26
timestamp 1644511149
transform 1 0 3496 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_38
timestamp 1644511149
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1644511149
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1644511149
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_312
timestamp 1644511149
transform 1 0 29808 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_324
timestamp 1644511149
transform 1 0 30912 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_336
timestamp 1644511149
transform 1 0 32016 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_348
timestamp 1644511149
transform 1 0 33120 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_360
timestamp 1644511149
transform 1 0 34224 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_412
timestamp 1644511149
transform 1 0 39008 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_425
timestamp 1644511149
transform 1 0 40204 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_429
timestamp 1644511149
transform 1 0 40572 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_441
timestamp 1644511149
transform 1 0 41676 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_453
timestamp 1644511149
transform 1 0 42780 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_465
timestamp 1644511149
transform 1 0 43884 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1644511149
transform 1 0 3864 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1644511149
transform 1 0 4968 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1644511149
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_101
timestamp 1644511149
transform 1 0 10396 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_133
timestamp 1644511149
transform 1 0 13340 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_139
timestamp 1644511149
transform 1 0 13892 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_151
timestamp 1644511149
transform 1 0 14996 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_163
timestamp 1644511149
transform 1 0 16100 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_216
timestamp 1644511149
transform 1 0 20976 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_454
timestamp 1644511149
transform 1 0 42872 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_469
timestamp 1644511149
transform 1 0 44252 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_494
timestamp 1644511149
transform 1 0 46552 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_502
timestamp 1644511149
transform 1 0 47288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1644511149
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1644511149
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_32
timestamp 1644511149
transform 1 0 4048 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_39
timestamp 1644511149
transform 1 0 4692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_51
timestamp 1644511149
transform 1 0 5796 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_63
timestamp 1644511149
transform 1 0 6900 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_75
timestamp 1644511149
transform 1 0 8004 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_122
timestamp 1644511149
transform 1 0 12328 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_134
timestamp 1644511149
transform 1 0 13432 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_202
timestamp 1644511149
transform 1 0 19688 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_234
timestamp 1644511149
transform 1 0 22632 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_246
timestamp 1644511149
transform 1 0 23736 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_344
timestamp 1644511149
transform 1 0 32752 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_353
timestamp 1644511149
transform 1 0 33580 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_361
timestamp 1644511149
transform 1 0 34316 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_405
timestamp 1644511149
transform 1 0 38364 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_417
timestamp 1644511149
transform 1 0 39468 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_455
timestamp 1644511149
transform 1 0 42964 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_463
timestamp 1644511149
transform 1 0 43700 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_13
timestamp 1644511149
transform 1 0 2300 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_20
timestamp 1644511149
transform 1 0 2944 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_45
timestamp 1644511149
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1644511149
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_131
timestamp 1644511149
transform 1 0 13156 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_156
timestamp 1644511149
transform 1 0 15456 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_228
timestamp 1644511149
transform 1 0 22080 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_240
timestamp 1644511149
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_252
timestamp 1644511149
transform 1 0 24288 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_362
timestamp 1644511149
transform 1 0 34408 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_374
timestamp 1644511149
transform 1 0 35512 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_386
timestamp 1644511149
transform 1 0 36616 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_422
timestamp 1644511149
transform 1 0 39928 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1644511149
transform 1 0 6900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_117
timestamp 1644511149
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_149
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_161
timestamp 1644511149
transform 1 0 15916 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_185
timestamp 1644511149
transform 1 0 18124 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_192
timestamp 1644511149
transform 1 0 18768 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_259
timestamp 1644511149
transform 1 0 24932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_266
timestamp 1644511149
transform 1 0 25576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1644511149
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_323
timestamp 1644511149
transform 1 0 30820 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_329
timestamp 1644511149
transform 1 0 31372 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1644511149
transform 1 0 31924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_405
timestamp 1644511149
transform 1 0 38364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1644511149
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_444
timestamp 1644511149
transform 1 0 41952 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_471
timestamp 1644511149
transform 1 0 44436 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0591_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31832 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0597_
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0598_
timestamp 1644511149
transform 1 0 35880 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0599_
timestamp 1644511149
transform 1 0 28520 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0600_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0601_
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0602_
timestamp 1644511149
transform 1 0 25760 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0603_
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20884 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0605_
timestamp 1644511149
transform 1 0 20608 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0606_
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0607_
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0608_
timestamp 1644511149
transform 1 0 27324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18676 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0613_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0614_
timestamp 1644511149
transform 1 0 13064 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0616_
timestamp 1644511149
transform 1 0 17572 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0618_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0619_
timestamp 1644511149
transform 1 0 15088 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0620_
timestamp 1644511149
transform 1 0 14628 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21620 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0623_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0626_
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0627_
timestamp 1644511149
transform 1 0 20056 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1644511149
transform 1 0 22172 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19872 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0630_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0632_
timestamp 1644511149
transform 1 0 17940 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0634_
timestamp 1644511149
transform 1 0 18400 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0635_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0636_
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0637_
timestamp 1644511149
transform 1 0 17020 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0639_
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0641_
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0644_
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1644511149
transform 1 0 18676 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0646_
timestamp 1644511149
transform 1 0 15088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0647_
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0648_
timestamp 1644511149
transform 1 0 14260 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0649_
timestamp 1644511149
transform 1 0 13432 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0650_
timestamp 1644511149
transform 1 0 15272 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0653_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1644511149
transform 1 0 12696 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1644511149
transform 1 0 16928 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0658_
timestamp 1644511149
transform 1 0 15364 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1644511149
transform 1 0 16744 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14812 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1644511149
transform 1 0 15824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0663_
timestamp 1644511149
transform 1 0 12512 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0664_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13800 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1644511149
transform 1 0 12328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11408 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0667_
timestamp 1644511149
transform 1 0 11684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1644511149
transform 1 0 12604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0669_
timestamp 1644511149
transform 1 0 11960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0670_
timestamp 1644511149
transform 1 0 11408 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1644511149
transform 1 0 12880 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1644511149
transform 1 0 12052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0673_
timestamp 1644511149
transform 1 0 10764 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1644511149
transform 1 0 11776 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0675_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0676_
timestamp 1644511149
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0677_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0678_
timestamp 1644511149
transform 1 0 11040 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1644511149
transform 1 0 12052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0680_
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0681_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10488 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1644511149
transform 1 0 12420 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0683_
timestamp 1644511149
transform 1 0 11592 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1644511149
transform 1 0 9752 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0691_
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0692_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0694_
timestamp 1644511149
transform 1 0 14904 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0695_
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1644511149
transform 1 0 14996 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0697_
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0698_
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1644511149
transform 1 0 15088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0700_
timestamp 1644511149
transform 1 0 13524 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1644511149
transform 1 0 14628 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0703_
timestamp 1644511149
transform 1 0 23828 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0704_
timestamp 1644511149
transform 1 0 17204 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0705_
timestamp 1644511149
transform 1 0 15272 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0706_
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0707_
timestamp 1644511149
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1644511149
transform 1 0 19320 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0709_
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0710_
timestamp 1644511149
transform 1 0 17572 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0712_
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0714_
timestamp 1644511149
transform 1 0 24840 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0715_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0716_
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0718_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0721_
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1644511149
transform 1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0726_
timestamp 1644511149
transform 1 0 24380 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0729_
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0730_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 29072 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0733_
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1644511149
transform 1 0 29716 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0736_
timestamp 1644511149
transform 1 0 28336 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0737_
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1644511149
transform 1 0 22816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0740_
timestamp 1644511149
transform 1 0 29716 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0741_
timestamp 1644511149
transform 1 0 29256 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0742_
timestamp 1644511149
transform 1 0 26404 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0743_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24196 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0745_
timestamp 1644511149
transform 1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0746_
timestamp 1644511149
transform 1 0 24932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0747_
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0748_
timestamp 1644511149
transform 1 0 26128 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0749_
timestamp 1644511149
transform 1 0 28520 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0750_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 1644511149
transform 1 0 29808 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0752_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1644511149
transform 1 0 23000 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0754_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0755_
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0756_
timestamp 1644511149
transform 1 0 28152 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0757_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _0758_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0759_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0760_
timestamp 1644511149
transform 1 0 33672 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0761_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0762_
timestamp 1644511149
transform 1 0 29624 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0763_
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0764_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21528 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0765_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0766_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0767_
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1644511149
transform 1 0 23276 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0769_
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0770_
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0771_
timestamp 1644511149
transform 1 0 22080 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0772_
timestamp 1644511149
transform 1 0 28704 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0773_
timestamp 1644511149
transform 1 0 28060 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0774_
timestamp 1644511149
transform 1 0 31188 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0775_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1644511149
transform 1 0 21344 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0777_
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0778_
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0779_
timestamp 1644511149
transform 1 0 27048 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0780_
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0782_
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0783_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29256 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0784_
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0785_
timestamp 1644511149
transform 1 0 22816 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0786_
timestamp 1644511149
transform 1 0 21896 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0787_
timestamp 1644511149
transform 1 0 25760 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0789_
timestamp 1644511149
transform 1 0 27784 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0790_
timestamp 1644511149
transform 1 0 26404 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0792_
timestamp 1644511149
transform 1 0 23460 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0793_
timestamp 1644511149
transform 1 0 29440 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0794_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1644511149
transform 1 0 26036 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0796_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0798_
timestamp 1644511149
transform 1 0 27600 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0799_
timestamp 1644511149
transform 1 0 26772 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0800_
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0801_
timestamp 1644511149
transform 1 0 27784 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0802_
timestamp 1644511149
transform 1 0 30084 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0803_
timestamp 1644511149
transform 1 0 28428 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0804_
timestamp 1644511149
transform 1 0 24288 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0805_
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0806_
timestamp 1644511149
transform 1 0 33028 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0807_
timestamp 1644511149
transform 1 0 30636 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0809_
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 1644511149
transform 1 0 29992 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29716 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0812_
timestamp 1644511149
transform 1 0 29624 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0813_
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1644511149
transform 1 0 33304 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0815_
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0816_
timestamp 1644511149
transform 1 0 33396 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0817_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32384 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0820_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0821_
timestamp 1644511149
transform 1 0 34408 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0823_
timestamp 1644511149
transform 1 0 31096 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1644511149
transform 1 0 31188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0825_
timestamp 1644511149
transform 1 0 30084 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0826_
timestamp 1644511149
transform 1 0 36156 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 1644511149
transform 1 0 36432 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0829_
timestamp 1644511149
transform 1 0 31832 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0830_
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0831_
timestamp 1644511149
transform 1 0 31924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0832_
timestamp 1644511149
transform 1 0 30820 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0833_
timestamp 1644511149
transform 1 0 33028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0834_
timestamp 1644511149
transform 1 0 32200 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0835_
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0836_
timestamp 1644511149
transform 1 0 33304 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1644511149
transform 1 0 33396 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0838_
timestamp 1644511149
transform 1 0 33304 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0839_
timestamp 1644511149
transform 1 0 31648 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 1644511149
transform 1 0 30544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1644511149
transform 1 0 30452 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0842_
timestamp 1644511149
transform 1 0 29900 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0843_
timestamp 1644511149
transform 1 0 27048 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0844_
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0845_
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0847_
timestamp 1644511149
transform 1 0 25576 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0848_
timestamp 1644511149
transform 1 0 24380 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0849_
timestamp 1644511149
transform 1 0 25300 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1644511149
transform 1 0 25668 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0851_
timestamp 1644511149
transform 1 0 24656 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1644511149
transform 1 0 30176 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0853_
timestamp 1644511149
transform 1 0 30728 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0856_
timestamp 1644511149
transform 1 0 32292 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0857_
timestamp 1644511149
transform 1 0 33396 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0858_
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0859_
timestamp 1644511149
transform 1 0 31188 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0861_
timestamp 1644511149
transform 1 0 30084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0862_
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0863_
timestamp 1644511149
transform 1 0 29624 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0864_
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0865_
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0866_
timestamp 1644511149
transform 1 0 31004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0867_
timestamp 1644511149
transform 1 0 30176 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0868_
timestamp 1644511149
transform 1 0 31004 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform 1 0 28152 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0872_
timestamp 1644511149
transform 1 0 28244 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0873_
timestamp 1644511149
transform 1 0 33396 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0874_
timestamp 1644511149
transform 1 0 26404 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0875_
timestamp 1644511149
transform 1 0 25392 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0876_
timestamp 1644511149
transform 1 0 25944 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 1644511149
transform 1 0 27600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0878_
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0879_
timestamp 1644511149
transform 1 0 28704 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0880_
timestamp 1644511149
transform 1 0 28612 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0883_
timestamp 1644511149
transform 1 0 25760 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0884_
timestamp 1644511149
transform 1 0 45448 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  _0885_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43516 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 38640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 42596 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45264 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 13616 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 20056 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0903_
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0909_
timestamp 1644511149
transform 1 0 45356 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44896 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 43976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45816 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 2760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 28796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0922_
timestamp 1644511149
transform 1 0 45356 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 23368 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0928_
timestamp 1644511149
transform 1 0 45080 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 41216 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 40296 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0934_
timestamp 1644511149
transform 1 0 43976 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 45080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 40296 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 38732 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 33304 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1644511149
transform 1 0 25944 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0941_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0947_
timestamp 1644511149
transform 1 0 25668 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 10488 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 2760 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0953_
timestamp 1644511149
transform 1 0 26128 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 42964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0959_
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 38088 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0965_
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 40296 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 30544 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0971_
timestamp 1644511149
transform 1 0 17940 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0972_
timestamp 1644511149
transform 1 0 16744 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 17664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0978_
timestamp 1644511149
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 14536 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 9568 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0984_
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 14168 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0990_
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0996_
timestamp 1644511149
transform 1 0 16652 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform 1 0 20516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 45632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1003_
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1004_
timestamp 1644511149
transform 1 0 21068 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43424 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1010_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1011_
timestamp 1644511149
transform 1 0 45264 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform 1 0 45632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1013_
timestamp 1644511149
transform 1 0 45080 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1014_
timestamp 1644511149
transform 1 0 45356 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1016_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1644511149
transform 1 0 44712 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1018_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1019_
timestamp 1644511149
transform 1 0 40204 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1644511149
transform 1 0 40112 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1021_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40112 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1022_
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1644511149
transform 1 0 40296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1024_
timestamp 1644511149
transform 1 0 40020 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1644511149
transform 1 0 41308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1026_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_2  _1027_
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _1028_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _1029_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1644511149
transform 1 0 26864 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 1644511149
transform 1 0 40388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1033_
timestamp 1644511149
transform 1 0 40480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1034_
timestamp 1644511149
transform 1 0 40756 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1035_
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1644511149
transform 1 0 42412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1039_
timestamp 1644511149
transform 1 0 41308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1040_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 1644511149
transform 1 0 42596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1042_
timestamp 1644511149
transform 1 0 42872 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1644511149
transform 1 0 43976 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _1044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41676 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1045_
timestamp 1644511149
transform 1 0 43700 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1046_
timestamp 1644511149
transform 1 0 43240 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1047_
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1048_
timestamp 1644511149
transform 1 0 43976 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1049_
timestamp 1644511149
transform 1 0 43056 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_2  _1050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42688 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _1051_
timestamp 1644511149
transform 1 0 43056 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1052_
timestamp 1644511149
transform 1 0 44160 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 1644511149
transform 1 0 42780 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1644511149
transform 1 0 43332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1055_
timestamp 1644511149
transform 1 0 43056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1056_
timestamp 1644511149
transform 1 0 43608 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1057_
timestamp 1644511149
transform 1 0 43056 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1058_
timestamp 1644511149
transform 1 0 39928 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1059_
timestamp 1644511149
transform 1 0 40940 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1060_
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1061_
timestamp 1644511149
transform 1 0 28152 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1062_
timestamp 1644511149
transform 1 0 28704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1063_
timestamp 1644511149
transform 1 0 31096 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1065_
timestamp 1644511149
transform 1 0 25576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1067_
timestamp 1644511149
transform 1 0 2668 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1069_
timestamp 1644511149
transform 1 0 43976 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1644511149
transform 1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1071_
timestamp 1644511149
transform 1 0 33396 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1073_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1075_
timestamp 1644511149
transform 1 0 43056 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1644511149
transform 1 0 42596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1077_
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1079_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1644511149
transform 1 0 27508 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1644511149
transform 1 0 27600 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1644511149
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1644511149
transform 1 0 33396 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1644511149
transform 1 0 32660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1644511149
transform 1 0 32752 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1644511149
transform 1 0 34776 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1089_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1644511149
transform 1 0 32384 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 35052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1095_
timestamp 1644511149
transform 1 0 34408 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 35880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 35236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 35236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1101_
timestamp 1644511149
transform 1 0 24472 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1644511149
transform 1 0 30728 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 31556 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1644511149
transform 1 0 24748 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1644511149
transform 1 0 28704 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 25668 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1107_
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 23092 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 20240 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 20884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1113_
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 20608 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 23276 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1644511149
transform 1 0 22080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1119_
timestamp 1644511149
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1120_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1121_
timestamp 1644511149
transform 1 0 21620 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1122_
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1123_
timestamp 1644511149
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1124_
timestamp 1644511149
transform 1 0 18400 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1125_
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1126_
timestamp 1644511149
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1127_
timestamp 1644511149
transform 1 0 14352 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1128_
timestamp 1644511149
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1644511149
transform 1 0 13064 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1130_
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1131_
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1132_
timestamp 1644511149
transform 1 0 10580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1133_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1134_
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1644511149
transform 1 0 10120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1136_
timestamp 1644511149
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1137_
timestamp 1644511149
transform 1 0 10672 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1139_
timestamp 1644511149
transform 1 0 10764 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1140_
timestamp 1644511149
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1644511149
transform 1 0 14720 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1142_
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1143_
timestamp 1644511149
transform 1 0 15456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1144_
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1145_
timestamp 1644511149
transform 1 0 15824 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1146_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1147_
timestamp 1644511149
transform 1 0 15824 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1149_
timestamp 1644511149
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1644511149
transform 1 0 16928 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1152_
timestamp 1644511149
transform 1 0 20976 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1153_
timestamp 1644511149
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1154_
timestamp 1644511149
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1155_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1644511149
transform 1 0 25024 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1644511149
transform 1 0 33856 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1644511149
transform 1 0 31188 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1644511149
transform 1 0 34500 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1644511149
transform 1 0 34776 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1644511149
transform 1 0 35880 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1644511149
transform 1 0 33120 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1644511149
transform 1 0 34132 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1644511149
transform 1 0 29624 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1644511149
transform 1 0 31096 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1644511149
transform 1 0 27232 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1644511149
transform 1 0 24656 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1644511149
transform 1 0 22448 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1644511149
transform 1 0 19136 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1644511149
transform 1 0 19504 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1644511149
transform 1 0 19320 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1644511149
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1644511149
transform 1 0 22724 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25024 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1190_
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1193_
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1644511149
transform 1 0 18032 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1644511149
transform 1 0 14720 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1196_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1200_
timestamp 1644511149
transform 1 0 10212 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1644511149
transform 1 0 11408 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1644511149
transform 1 0 9844 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1204_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1205_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1644511149
transform 1 0 13616 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1208_
timestamp 1644511149
transform 1 0 15732 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1644511149
transform 1 0 16192 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1644511149
transform 1 0 15640 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1212_
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1214_
timestamp 1644511149
transform 1 0 16560 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1215_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1216_
timestamp 1644511149
transform 1 0 17204 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1217_
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1220_
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1221__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1222__82
timestamp 1644511149
transform 1 0 32476 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1223__83
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1224__84
timestamp 1644511149
transform 1 0 47472 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1225__85
timestamp 1644511149
transform 1 0 47472 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1226__86
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1227__87
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1228__88
timestamp 1644511149
transform 1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1229__89
timestamp 1644511149
transform 1 0 10488 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1230__90
timestamp 1644511149
transform 1 0 25300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1231__91
timestamp 1644511149
transform 1 0 47472 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1232__92
timestamp 1644511149
transform 1 0 2668 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1233__93
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1234__94
timestamp 1644511149
transform 1 0 4416 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1235__95
timestamp 1644511149
transform 1 0 1840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1236__96
timestamp 1644511149
transform 1 0 43608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1237__97
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1238__98
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1239__99
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1240__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1241__101
timestamp 1644511149
transform 1 0 38088 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1242__102
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1243__103
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1244__104
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1245__105
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1246__106
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1247__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1248__108
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1249__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1250__110
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1251__111
timestamp 1644511149
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1252__112
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1253__113
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1254__114
timestamp 1644511149
transform 1 0 45632 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1255__115
timestamp 1644511149
transform 1 0 37904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1256__116
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1257__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1258__118
timestamp 1644511149
transform 1 0 12880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1259__119
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1260__120
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1261__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1262__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1263__123
timestamp 1644511149
transform 1 0 46368 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1264__124
timestamp 1644511149
transform 1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1265__125
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1266__126
timestamp 1644511149
transform 1 0 19412 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1267__127
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1268__128
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1269__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1270__130
timestamp 1644511149
transform 1 0 46184 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1271__131
timestamp 1644511149
transform 1 0 1840 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1272__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1273__133
timestamp 1644511149
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1274__134
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1275__135
timestamp 1644511149
transform 1 0 43240 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1277_
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1278_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1279_
timestamp 1644511149
transform 1 0 41216 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1280_
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1281_
timestamp 1644511149
transform 1 0 40020 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1282_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1644511149
transform 1 0 40204 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1644511149
transform 1 0 38640 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1644511149
transform 1 0 32476 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 20700 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 10396 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 1932 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 3312 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 42780 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 41032 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 45172 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 21988 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 16376 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1315_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1316_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1317_
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1318_
timestamp 1644511149
transform 1 0 14260 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1319_
timestamp 1644511149
transform 1 0 8648 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1320_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1321_
timestamp 1644511149
transform 1 0 13616 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1322_
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1323_
timestamp 1644511149
transform 1 0 9384 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1324_
timestamp 1644511149
transform 1 0 14168 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1325_
timestamp 1644511149
transform 1 0 14168 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1326_
timestamp 1644511149
transform 1 0 9108 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1327_
timestamp 1644511149
transform 1 0 9384 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1328_
timestamp 1644511149
transform 1 0 13800 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1329_
timestamp 1644511149
transform 1 0 17940 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1330_
timestamp 1644511149
transform 1 0 18124 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1331_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1332_
timestamp 1644511149
transform 1 0 13892 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1333_
timestamp 1644511149
transform 1 0 19412 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1334_
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1335_
timestamp 1644511149
transform 1 0 20240 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1336_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1337_
timestamp 1644511149
transform 1 0 30544 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1338_
timestamp 1644511149
transform 1 0 24104 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1339_
timestamp 1644511149
transform 1 0 23000 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1340_
timestamp 1644511149
transform 1 0 9292 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1341_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1342_
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1343_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1344_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1345_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1346_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 37812 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 42504 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 13524 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 46276 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 46276 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 27692 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 25484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 30544 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 24564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 31280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 31188 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1644511149
transform 1 0 18216 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 47288 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 44436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 37444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1644511149
transform 1 0 47840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1644511149
transform 1 0 47840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1644511149
transform 1 0 46736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1644511149
transform 1 0 46184 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1644511149
transform 1 0 46184 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 31004 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1644511149
transform 1 0 43884 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46184 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 45080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40204 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 40756 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 40296 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 40940 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 40204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 39652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 18032 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 19320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31556 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 25392 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45080 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ext_inputs\[4\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 25392 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35144 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42780 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37352 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 29532 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 29624 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 43976 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45724 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 45724 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 40756 0 1 22848
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
