magic
tech sky130A
magscale 1 2
timestamp 1654258838
<< viali >>
rect 16911 47141 16945 47175
rect 29929 47141 29963 47175
rect 47961 47141 47995 47175
rect 2053 47073 2087 47107
rect 30757 47073 30791 47107
rect 43177 47073 43211 47107
rect 47041 47073 47075 47107
rect 1777 47005 1811 47039
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6377 47005 6411 47039
rect 7297 47005 7331 47039
rect 9413 47005 9447 47039
rect 11713 47005 11747 47039
rect 12357 47005 12391 47039
rect 12633 47005 12667 47039
rect 15485 47005 15519 47039
rect 16681 47005 16715 47039
rect 20729 47005 20763 47039
rect 22017 47005 22051 47039
rect 28733 47005 28767 47039
rect 29745 47005 29779 47039
rect 31033 47005 31067 47039
rect 38393 47005 38427 47039
rect 40509 47005 40543 47039
rect 41889 47005 41923 47039
rect 42625 47005 42659 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 2789 46937 2823 46971
rect 4077 46937 4111 46971
rect 4997 46937 5031 46971
rect 6653 46937 6687 46971
rect 9597 46937 9631 46971
rect 11897 46937 11931 46971
rect 14565 46937 14599 46971
rect 15669 46937 15703 46971
rect 19717 46937 19751 46971
rect 20085 46937 20119 46971
rect 28549 46937 28583 46971
rect 40325 46937 40359 46971
rect 42809 46937 42843 46971
rect 45385 46937 45419 46971
rect 2881 46869 2915 46903
rect 7481 46869 7515 46903
rect 14657 46869 14691 46903
rect 21833 46869 21867 46903
rect 1869 46597 1903 46631
rect 5825 46597 5859 46631
rect 32321 46597 32355 46631
rect 38117 46529 38151 46563
rect 47961 46529 47995 46563
rect 3985 46461 4019 46495
rect 4169 46461 4203 46495
rect 13185 46461 13219 46495
rect 13645 46461 13679 46495
rect 13829 46461 13863 46495
rect 14289 46461 14323 46495
rect 18981 46461 19015 46495
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 26341 46461 26375 46495
rect 26985 46461 27019 46495
rect 27169 46461 27203 46495
rect 27721 46461 27755 46495
rect 31585 46461 31619 46495
rect 32137 46461 32171 46495
rect 32597 46461 32631 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 2053 46393 2087 46427
rect 2881 46325 2915 46359
rect 10701 46325 10735 46359
rect 25513 46325 25547 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 4445 46121 4479 46155
rect 5181 46121 5215 46155
rect 14197 46121 14231 46155
rect 18613 46121 18647 46155
rect 27629 46121 27663 46155
rect 38301 46121 38335 46155
rect 1409 45985 1443 46019
rect 2789 45985 2823 46019
rect 10425 45985 10459 46019
rect 11069 45985 11103 46019
rect 26249 45985 26283 46019
rect 41337 45985 41371 46019
rect 41889 45985 41923 46019
rect 46305 45985 46339 46019
rect 47041 45985 47075 46019
rect 5089 45917 5123 45951
rect 14105 45917 14139 45951
rect 18521 45917 18555 45951
rect 19533 45917 19567 45951
rect 20177 45917 20211 45951
rect 22017 45917 22051 45951
rect 25237 45917 25271 45951
rect 27537 45917 27571 45951
rect 38209 45917 38243 45951
rect 44005 45917 44039 45951
rect 45661 45917 45695 45951
rect 1593 45849 1627 45883
rect 10609 45849 10643 45883
rect 19625 45849 19659 45883
rect 20361 45849 20395 45883
rect 25421 45849 25455 45883
rect 41521 45849 41555 45883
rect 44189 45849 44223 45883
rect 46489 45849 46523 45883
rect 45753 45781 45787 45815
rect 2237 45577 2271 45611
rect 10609 45577 10643 45611
rect 26157 45577 26191 45611
rect 41429 45577 41463 45611
rect 42533 45577 42567 45611
rect 43637 45509 43671 45543
rect 44373 45509 44407 45543
rect 46581 45509 46615 45543
rect 47685 45509 47719 45543
rect 2145 45441 2179 45475
rect 10517 45441 10551 45475
rect 26065 45441 26099 45475
rect 41337 45441 41371 45475
rect 42441 45441 42475 45475
rect 43545 45441 43579 45475
rect 47593 45441 47627 45475
rect 44189 45373 44223 45407
rect 45385 45373 45419 45407
rect 46673 45237 46707 45271
rect 43085 45033 43119 45067
rect 44465 44897 44499 44931
rect 48145 44897 48179 44931
rect 38669 44829 38703 44863
rect 42993 44829 43027 44863
rect 45477 44829 45511 44863
rect 46305 44829 46339 44863
rect 45661 44761 45695 44795
rect 46489 44761 46523 44795
rect 38761 44693 38795 44727
rect 45661 44489 45695 44523
rect 47685 44489 47719 44523
rect 38761 44421 38795 44455
rect 44465 44353 44499 44387
rect 45109 44353 45143 44387
rect 45569 44353 45603 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 38577 44285 38611 44319
rect 40049 44285 40083 44319
rect 46305 44217 46339 44251
rect 46949 44149 46983 44183
rect 45845 43945 45879 43979
rect 46305 43809 46339 43843
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 26801 43741 26835 43775
rect 26893 43605 26927 43639
rect 1409 43265 1443 43299
rect 45937 43265 45971 43299
rect 46581 43265 46615 43299
rect 1593 43197 1627 43231
rect 47777 43061 47811 43095
rect 46305 42721 46339 42755
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 2145 41225 2179 41259
rect 46857 41225 46891 41259
rect 2053 41089 2087 41123
rect 46765 41089 46799 41123
rect 47961 41089 47995 41123
rect 48145 40953 48179 40987
rect 47685 40681 47719 40715
rect 1869 40409 1903 40443
rect 1961 40341 1995 40375
rect 47777 39797 47811 39831
rect 25421 39457 25455 39491
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 22477 39389 22511 39423
rect 25237 39389 25271 39423
rect 22569 39321 22603 39355
rect 46489 39321 46523 39355
rect 24869 39253 24903 39287
rect 25329 39253 25363 39287
rect 25053 39049 25087 39083
rect 20085 38981 20119 39015
rect 20729 38981 20763 39015
rect 19441 38913 19475 38947
rect 20913 38913 20947 38947
rect 24685 38913 24719 38947
rect 47685 38913 47719 38947
rect 22109 38845 22143 38879
rect 22385 38845 22419 38879
rect 23857 38845 23891 38879
rect 24593 38845 24627 38879
rect 47869 38845 47903 38879
rect 21097 38709 21131 38743
rect 22937 38505 22971 38539
rect 24409 38369 24443 38403
rect 18245 38301 18279 38335
rect 19441 38301 19475 38335
rect 20821 38301 20855 38335
rect 23121 38301 23155 38335
rect 23581 38301 23615 38335
rect 23765 38301 23799 38335
rect 27905 38301 27939 38335
rect 47685 38301 47719 38335
rect 18521 38233 18555 38267
rect 20085 38233 20119 38267
rect 21373 38233 21407 38267
rect 24685 38233 24719 38267
rect 23673 38165 23707 38199
rect 26157 38165 26191 38199
rect 27997 38165 28031 38199
rect 18705 37961 18739 37995
rect 20821 37961 20855 37995
rect 24593 37961 24627 37995
rect 25513 37961 25547 37995
rect 18521 37825 18555 37859
rect 19441 37825 19475 37859
rect 20729 37825 20763 37859
rect 24317 37825 24351 37859
rect 24409 37825 24443 37859
rect 24685 37825 24719 37859
rect 25421 37825 25455 37859
rect 26985 37825 27019 37859
rect 29193 37825 29227 37859
rect 47593 37825 47627 37859
rect 19717 37757 19751 37791
rect 24501 37757 24535 37791
rect 27261 37757 27295 37791
rect 28733 37621 28767 37655
rect 29285 37621 29319 37655
rect 47685 37621 47719 37655
rect 19625 37417 19659 37451
rect 25513 37417 25547 37451
rect 25421 37281 25455 37315
rect 27261 37281 27295 37315
rect 48145 37281 48179 37315
rect 2053 37213 2087 37247
rect 19441 37213 19475 37247
rect 21833 37213 21867 37247
rect 24501 37213 24535 37247
rect 25513 37213 25547 37247
rect 26801 37213 26835 37247
rect 30757 37213 30791 37247
rect 46305 37213 46339 37247
rect 25237 37145 25271 37179
rect 27537 37145 27571 37179
rect 46489 37145 46523 37179
rect 21925 37077 21959 37111
rect 24685 37077 24719 37111
rect 25697 37077 25731 37111
rect 26617 37077 26651 37111
rect 29009 37077 29043 37111
rect 30849 37077 30883 37111
rect 24961 36873 24995 36907
rect 26065 36873 26099 36907
rect 27077 36873 27111 36907
rect 27445 36873 27479 36907
rect 25421 36805 25455 36839
rect 1777 36737 1811 36771
rect 22017 36737 22051 36771
rect 22201 36737 22235 36771
rect 22293 36737 22327 36771
rect 24685 36737 24719 36771
rect 24777 36737 24811 36771
rect 25881 36737 25915 36771
rect 27261 36737 27295 36771
rect 27537 36737 27571 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 24961 36669 24995 36703
rect 25697 36669 25731 36703
rect 29561 36669 29595 36703
rect 29837 36669 29871 36703
rect 21833 36533 21867 36567
rect 25881 36533 25915 36567
rect 31309 36533 31343 36567
rect 2237 36329 2271 36363
rect 26433 36329 26467 36363
rect 27629 36329 27663 36363
rect 29561 36329 29595 36363
rect 23673 36261 23707 36295
rect 24961 36261 24995 36295
rect 27537 36261 27571 36295
rect 20913 36193 20947 36227
rect 23397 36193 23431 36227
rect 30021 36193 30055 36227
rect 30573 36193 30607 36227
rect 2145 36125 2179 36159
rect 19901 36125 19935 36159
rect 23305 36125 23339 36159
rect 24409 36125 24443 36159
rect 24685 36125 24719 36159
rect 24777 36125 24811 36159
rect 25421 36125 25455 36159
rect 26249 36125 26283 36159
rect 28089 36125 28123 36159
rect 29745 36125 29779 36159
rect 29837 36125 29871 36159
rect 30113 36125 30147 36159
rect 30757 36125 30791 36159
rect 32045 36125 32079 36159
rect 21189 36057 21223 36091
rect 24593 36057 24627 36091
rect 25605 36057 25639 36091
rect 27169 36057 27203 36091
rect 30941 36057 30975 36091
rect 19993 35989 20027 36023
rect 22661 35989 22695 36023
rect 25789 35989 25823 36023
rect 28181 35989 28215 36023
rect 32137 35989 32171 36023
rect 22569 35785 22603 35819
rect 27721 35785 27755 35819
rect 28381 35785 28415 35819
rect 28549 35785 28583 35819
rect 29745 35785 29779 35819
rect 29929 35785 29963 35819
rect 31217 35785 31251 35819
rect 19441 35717 19475 35751
rect 27077 35717 27111 35751
rect 28181 35717 28215 35751
rect 31033 35717 31067 35751
rect 1593 35649 1627 35683
rect 21833 35649 21867 35683
rect 22017 35649 22051 35683
rect 22201 35649 22235 35683
rect 22385 35649 22419 35683
rect 23213 35649 23247 35683
rect 23397 35649 23431 35683
rect 24593 35649 24627 35683
rect 25237 35649 25271 35683
rect 25513 35649 25547 35683
rect 27445 35649 27479 35683
rect 29870 35649 29904 35683
rect 30389 35649 30423 35683
rect 30849 35649 30883 35683
rect 48145 35649 48179 35683
rect 19165 35581 19199 35615
rect 20913 35581 20947 35615
rect 22109 35581 22143 35615
rect 23489 35581 23523 35615
rect 25329 35581 25363 35615
rect 27537 35581 27571 35615
rect 32137 35581 32171 35615
rect 32413 35581 32447 35615
rect 23029 35513 23063 35547
rect 30297 35513 30331 35547
rect 1409 35445 1443 35479
rect 24685 35445 24719 35479
rect 25513 35445 25547 35479
rect 25697 35445 25731 35479
rect 28365 35445 28399 35479
rect 33885 35445 33919 35479
rect 47961 35445 47995 35479
rect 21649 35241 21683 35275
rect 21833 35241 21867 35275
rect 22661 35241 22695 35275
rect 24777 35241 24811 35275
rect 26985 35241 27019 35275
rect 28089 35241 28123 35275
rect 28549 35241 28583 35275
rect 32505 35241 32539 35275
rect 26433 35173 26467 35207
rect 22569 35105 22603 35139
rect 30757 35105 30791 35139
rect 32045 35105 32079 35139
rect 32137 35105 32171 35139
rect 21281 35037 21315 35071
rect 21649 35037 21683 35071
rect 22661 35037 22695 35071
rect 24409 35037 24443 35071
rect 26249 35037 26283 35071
rect 27169 35037 27203 35071
rect 27261 35037 27295 35071
rect 27629 35037 27663 35071
rect 28273 35037 28307 35071
rect 28365 35037 28399 35071
rect 28641 35037 28675 35071
rect 29929 35037 29963 35071
rect 30113 35037 30147 35071
rect 30941 35037 30975 35071
rect 31033 35037 31067 35071
rect 31217 35037 31251 35071
rect 31309 35037 31343 35071
rect 31769 35037 31803 35071
rect 31953 35037 31987 35071
rect 32321 35037 32355 35071
rect 48145 35037 48179 35071
rect 22385 34969 22419 35003
rect 24593 34969 24627 35003
rect 27354 34969 27388 35003
rect 27471 34969 27505 35003
rect 22845 34901 22879 34935
rect 30021 34901 30055 34935
rect 47961 34901 47995 34935
rect 28917 34697 28951 34731
rect 29929 34697 29963 34731
rect 23121 34629 23155 34663
rect 30389 34629 30423 34663
rect 22201 34561 22235 34595
rect 22477 34561 22511 34595
rect 22937 34561 22971 34595
rect 24593 34561 24627 34595
rect 27537 34561 27571 34595
rect 28733 34561 28767 34595
rect 29561 34561 29595 34595
rect 30665 34561 30699 34595
rect 47777 34561 47811 34595
rect 18613 34493 18647 34527
rect 20361 34493 20395 34527
rect 22385 34493 22419 34527
rect 24685 34493 24719 34527
rect 27629 34493 27663 34527
rect 27813 34493 27847 34527
rect 29653 34493 29687 34527
rect 30573 34493 30607 34527
rect 18876 34357 18910 34391
rect 22017 34357 22051 34391
rect 23305 34357 23339 34391
rect 27721 34357 27755 34391
rect 29745 34357 29779 34391
rect 30389 34357 30423 34391
rect 30849 34357 30883 34391
rect 47593 34357 47627 34391
rect 19625 34153 19659 34187
rect 21557 34153 21591 34187
rect 22385 34153 22419 34187
rect 28733 34153 28767 34187
rect 31309 34153 31343 34187
rect 21189 34017 21223 34051
rect 24409 34017 24443 34051
rect 29929 34017 29963 34051
rect 31493 34017 31527 34051
rect 47133 34017 47167 34051
rect 47685 34017 47719 34051
rect 19533 33949 19567 33983
rect 20821 33949 20855 33983
rect 21005 33949 21039 33983
rect 21097 33949 21131 33983
rect 21373 33949 21407 33983
rect 22017 33949 22051 33983
rect 22385 33949 22419 33983
rect 23029 33949 23063 33983
rect 29745 33949 29779 33983
rect 30021 33949 30055 33983
rect 30481 33949 30515 33983
rect 31217 33949 31251 33983
rect 24685 33881 24719 33915
rect 27261 33881 27295 33915
rect 28641 33881 28675 33915
rect 47225 33881 47259 33915
rect 22569 33813 22603 33847
rect 23213 33813 23247 33847
rect 26157 33813 26191 33847
rect 27353 33813 27387 33847
rect 29561 33813 29595 33847
rect 30665 33813 30699 33847
rect 31493 33813 31527 33847
rect 23305 33609 23339 33643
rect 48053 33609 48087 33643
rect 23213 33541 23247 33575
rect 29285 33541 29319 33575
rect 1593 33473 1627 33507
rect 2237 33473 2271 33507
rect 19809 33473 19843 33507
rect 22017 33473 22051 33507
rect 24119 33473 24153 33507
rect 25237 33473 25271 33507
rect 25329 33473 25363 33507
rect 25605 33473 25639 33507
rect 46857 33473 46891 33507
rect 47593 33473 47627 33507
rect 2421 33405 2455 33439
rect 4077 33405 4111 33439
rect 22293 33405 22327 33439
rect 23949 33405 23983 33439
rect 29009 33405 29043 33439
rect 24409 33337 24443 33371
rect 1409 33269 1443 33303
rect 19901 33269 19935 33303
rect 21833 33269 21867 33303
rect 22201 33269 22235 33303
rect 25053 33269 25087 33303
rect 25513 33269 25547 33303
rect 30757 33269 30791 33303
rect 46949 33269 46983 33303
rect 47869 33269 47903 33303
rect 2789 33065 2823 33099
rect 3801 33065 3835 33099
rect 21925 33065 21959 33099
rect 23029 33065 23063 33099
rect 24777 33065 24811 33099
rect 28273 33065 28307 33099
rect 30757 33065 30791 33099
rect 29561 32997 29595 33031
rect 31401 32997 31435 33031
rect 1409 32929 1443 32963
rect 3157 32929 3191 32963
rect 19533 32929 19567 32963
rect 22385 32929 22419 32963
rect 24409 32929 24443 32963
rect 27537 32929 27571 32963
rect 30021 32929 30055 32963
rect 47593 32929 47627 32963
rect 1685 32861 1719 32895
rect 2697 32861 2731 32895
rect 3985 32861 4019 32895
rect 19257 32861 19291 32895
rect 22109 32861 22143 32895
rect 22201 32861 22235 32895
rect 22477 32861 22511 32895
rect 22937 32861 22971 32895
rect 23121 32861 23155 32895
rect 24593 32861 24627 32895
rect 24869 32861 24903 32895
rect 28181 32861 28215 32895
rect 29745 32861 29779 32895
rect 29837 32861 29871 32895
rect 30113 32861 30147 32895
rect 31309 32861 31343 32895
rect 31493 32861 31527 32895
rect 32321 32861 32355 32895
rect 32597 32861 32631 32895
rect 46857 32861 46891 32895
rect 47317 32861 47351 32895
rect 26709 32793 26743 32827
rect 27353 32793 27387 32827
rect 30665 32793 30699 32827
rect 32137 32793 32171 32827
rect 21005 32725 21039 32759
rect 26985 32725 27019 32759
rect 27445 32725 27479 32759
rect 32505 32725 32539 32759
rect 21281 32521 21315 32555
rect 23581 32521 23615 32555
rect 25053 32521 25087 32555
rect 30113 32521 30147 32555
rect 31585 32521 31619 32555
rect 31309 32453 31343 32487
rect 32413 32453 32447 32487
rect 18153 32385 18187 32419
rect 21005 32385 21039 32419
rect 22109 32385 22143 32419
rect 23121 32385 23155 32419
rect 23397 32385 23431 32419
rect 24041 32385 24075 32419
rect 24225 32385 24259 32419
rect 24961 32385 24995 32419
rect 27169 32385 27203 32419
rect 27905 32385 27939 32419
rect 29193 32385 29227 32419
rect 30021 32385 30055 32419
rect 31033 32385 31067 32419
rect 31217 32385 31251 32419
rect 31401 32385 31435 32419
rect 32137 32385 32171 32419
rect 47593 32385 47627 32419
rect 1777 32317 1811 32351
rect 1961 32317 1995 32351
rect 2789 32317 2823 32351
rect 18429 32317 18463 32351
rect 21281 32317 21315 32351
rect 21833 32317 21867 32351
rect 23213 32317 23247 32351
rect 29285 32317 29319 32351
rect 19901 32249 19935 32283
rect 21097 32181 21131 32215
rect 23121 32181 23155 32215
rect 24409 32181 24443 32215
rect 26985 32181 27019 32215
rect 27997 32181 28031 32215
rect 29561 32181 29595 32215
rect 33885 32181 33919 32215
rect 47685 32181 47719 32215
rect 1685 31977 1719 32011
rect 2237 31977 2271 32011
rect 19441 31977 19475 32011
rect 21925 31977 21959 32011
rect 22661 31977 22695 32011
rect 24777 31977 24811 32011
rect 25237 31977 25271 32011
rect 32505 31977 32539 32011
rect 33333 31977 33367 32011
rect 22201 31909 22235 31943
rect 3985 31841 4019 31875
rect 4629 31841 4663 31875
rect 21925 31841 21959 31875
rect 22845 31841 22879 31875
rect 24869 31841 24903 31875
rect 26065 31841 26099 31875
rect 26341 31841 26375 31875
rect 27813 31841 27847 31875
rect 32137 31841 32171 31875
rect 46305 31841 46339 31875
rect 46489 31841 46523 31875
rect 48145 31841 48179 31875
rect 2145 31773 2179 31807
rect 3801 31773 3835 31807
rect 17785 31773 17819 31807
rect 18245 31773 18279 31807
rect 19349 31773 19383 31807
rect 21833 31773 21867 31807
rect 22937 31773 22971 31807
rect 24777 31773 24811 31807
rect 25053 31773 25087 31807
rect 28273 31773 28307 31807
rect 29929 31773 29963 31807
rect 30113 31773 30147 31807
rect 32229 31773 32263 31807
rect 33241 31773 33275 31807
rect 22661 31705 22695 31739
rect 28365 31705 28399 31739
rect 18337 31637 18371 31671
rect 23121 31637 23155 31671
rect 30021 31637 30055 31671
rect 24685 31433 24719 31467
rect 28641 31433 28675 31467
rect 18521 31365 18555 31399
rect 26065 31365 26099 31399
rect 26265 31365 26299 31399
rect 29653 31365 29687 31399
rect 18337 31297 18371 31331
rect 22017 31297 22051 31331
rect 22845 31297 22879 31331
rect 23029 31297 23063 31331
rect 23765 31297 23799 31331
rect 23949 31297 23983 31331
rect 24041 31297 24075 31331
rect 24593 31297 24627 31331
rect 27353 31297 27387 31331
rect 30849 31297 30883 31331
rect 20177 31229 20211 31263
rect 22109 31229 22143 31263
rect 22385 31229 22419 31263
rect 31217 31229 31251 31263
rect 22845 31161 22879 31195
rect 29837 31161 29871 31195
rect 31309 31161 31343 31195
rect 23581 31093 23615 31127
rect 26249 31093 26283 31127
rect 26433 31093 26467 31127
rect 31014 31093 31048 31127
rect 31125 31093 31159 31127
rect 22477 30889 22511 30923
rect 23581 30889 23615 30923
rect 25789 30889 25823 30923
rect 27537 30889 27571 30923
rect 28181 30889 28215 30923
rect 33333 30821 33367 30855
rect 20453 30753 20487 30787
rect 23489 30753 23523 30787
rect 24961 30753 24995 30787
rect 27077 30753 27111 30787
rect 29561 30753 29595 30787
rect 31309 30753 31343 30787
rect 32229 30753 32263 30787
rect 34713 30753 34747 30787
rect 47685 30753 47719 30787
rect 20361 30685 20395 30719
rect 21833 30685 21867 30719
rect 21926 30685 21960 30719
rect 22201 30685 22235 30719
rect 22298 30685 22332 30719
rect 23213 30685 23247 30719
rect 25145 30685 25179 30719
rect 25789 30685 25823 30719
rect 25973 30685 26007 30719
rect 27169 30685 27203 30719
rect 27997 30685 28031 30719
rect 28825 30685 28859 30719
rect 31769 30685 31803 30719
rect 31861 30685 31895 30719
rect 32045 30685 32079 30719
rect 33149 30685 33183 30719
rect 33793 30685 33827 30719
rect 22109 30617 22143 30651
rect 29837 30617 29871 30651
rect 32965 30617 32999 30651
rect 34989 30617 35023 30651
rect 46857 30617 46891 30651
rect 46949 30617 46983 30651
rect 20729 30549 20763 30583
rect 23765 30549 23799 30583
rect 25329 30549 25363 30583
rect 28917 30549 28951 30583
rect 33885 30549 33919 30583
rect 36461 30549 36495 30583
rect 27261 30345 27295 30379
rect 29561 30345 29595 30379
rect 24133 30277 24167 30311
rect 29285 30277 29319 30311
rect 34161 30277 34195 30311
rect 34805 30277 34839 30311
rect 15117 30209 15151 30243
rect 19717 30209 19751 30243
rect 20545 30209 20579 30243
rect 20729 30209 20763 30243
rect 20821 30209 20855 30243
rect 21097 30209 21131 30243
rect 25053 30209 25087 30243
rect 25237 30209 25271 30243
rect 25329 30209 25363 30243
rect 27077 30209 27111 30243
rect 28181 30209 28215 30243
rect 28924 30209 28958 30243
rect 29055 30209 29089 30243
rect 29193 30209 29227 30243
rect 29423 30209 29457 30243
rect 30849 30209 30883 30243
rect 31033 30209 31067 30243
rect 32137 30209 32171 30243
rect 33425 30209 33459 30243
rect 33609 30209 33643 30243
rect 33701 30209 33735 30243
rect 33977 30209 34011 30243
rect 34713 30209 34747 30243
rect 17417 30141 17451 30175
rect 17601 30141 17635 30175
rect 19257 30141 19291 30175
rect 20913 30141 20947 30175
rect 32413 30141 32447 30175
rect 33793 30141 33827 30175
rect 15209 30005 15243 30039
rect 19809 30005 19843 30039
rect 21281 30005 21315 30039
rect 24225 30005 24259 30039
rect 24869 30005 24903 30039
rect 28365 30005 28399 30039
rect 30849 30005 30883 30039
rect 27077 29801 27111 29835
rect 28641 29801 28675 29835
rect 31585 29801 31619 29835
rect 32689 29801 32723 29835
rect 27261 29733 27295 29767
rect 31769 29733 31803 29767
rect 14933 29665 14967 29699
rect 16497 29665 16531 29699
rect 19533 29665 19567 29699
rect 32321 29665 32355 29699
rect 32597 29665 32631 29699
rect 33701 29665 33735 29699
rect 47593 29665 47627 29699
rect 14105 29597 14139 29631
rect 14749 29597 14783 29631
rect 19257 29597 19291 29631
rect 23029 29597 23063 29631
rect 23213 29597 23247 29631
rect 23305 29597 23339 29631
rect 23397 29597 23431 29631
rect 23581 29597 23615 29631
rect 24501 29597 24535 29631
rect 24649 29597 24683 29631
rect 25007 29597 25041 29631
rect 25605 29597 25639 29631
rect 27815 29597 27849 29631
rect 28457 29597 28491 29631
rect 30573 29597 30607 29631
rect 31401 29597 31435 29631
rect 31585 29597 31619 29631
rect 32229 29597 32263 29631
rect 32505 29597 32539 29631
rect 33333 29597 33367 29631
rect 33517 29597 33551 29631
rect 33609 29597 33643 29631
rect 33885 29597 33919 29631
rect 47317 29597 47351 29631
rect 24777 29529 24811 29563
rect 24869 29529 24903 29563
rect 26893 29529 26927 29563
rect 30757 29529 30791 29563
rect 14197 29461 14231 29495
rect 21005 29461 21039 29495
rect 23765 29461 23799 29495
rect 25145 29461 25179 29495
rect 25697 29461 25731 29495
rect 27093 29461 27127 29495
rect 27905 29461 27939 29495
rect 34069 29461 34103 29495
rect 10977 29257 11011 29291
rect 21925 29257 21959 29291
rect 25053 29257 25087 29291
rect 27721 29257 27755 29291
rect 28365 29257 28399 29291
rect 30297 29257 30331 29291
rect 31585 29257 31619 29291
rect 32965 29257 32999 29291
rect 35725 29257 35759 29291
rect 11805 29189 11839 29223
rect 14473 29189 14507 29223
rect 20177 29189 20211 29223
rect 23581 29189 23615 29223
rect 31217 29189 31251 29223
rect 34253 29189 34287 29223
rect 10609 29121 10643 29155
rect 19165 29121 19199 29155
rect 20085 29121 20119 29155
rect 20269 29121 20303 29155
rect 20913 29121 20947 29155
rect 21097 29121 21131 29155
rect 21833 29121 21867 29155
rect 22017 29121 22051 29155
rect 25881 29121 25915 29155
rect 27813 29121 27847 29155
rect 28273 29121 28307 29155
rect 29469 29121 29503 29155
rect 30113 29121 30147 29155
rect 31401 29121 31435 29155
rect 32413 29121 32447 29155
rect 33977 29121 34011 29155
rect 27537 29087 27571 29121
rect 10701 29053 10735 29087
rect 11529 29053 11563 29087
rect 14289 29053 14323 29087
rect 14749 29053 14783 29087
rect 16681 29053 16715 29087
rect 16865 29053 16899 29087
rect 17141 29053 17175 29087
rect 19257 29053 19291 29087
rect 21189 29053 21223 29087
rect 23305 29053 23339 29087
rect 32689 29053 32723 29087
rect 13277 28985 13311 29019
rect 27353 28985 27387 29019
rect 20729 28917 20763 28951
rect 25973 28917 26007 28951
rect 29561 28917 29595 28951
rect 32781 28917 32815 28951
rect 10701 28713 10735 28747
rect 12449 28713 12483 28747
rect 15853 28713 15887 28747
rect 16405 28713 16439 28747
rect 17417 28713 17451 28747
rect 21557 28713 21591 28747
rect 22845 28713 22879 28747
rect 26433 28713 26467 28747
rect 27077 28713 27111 28747
rect 30113 28713 30147 28747
rect 32137 28713 32171 28747
rect 32781 28713 32815 28747
rect 34805 28713 34839 28747
rect 10057 28645 10091 28679
rect 21005 28645 21039 28679
rect 27813 28645 27847 28679
rect 19257 28577 19291 28611
rect 19533 28577 19567 28611
rect 24961 28577 24995 28611
rect 30665 28577 30699 28611
rect 32229 28577 32263 28611
rect 32965 28577 32999 28611
rect 9965 28509 9999 28543
rect 10609 28509 10643 28543
rect 10793 28509 10827 28543
rect 11253 28509 11287 28543
rect 11437 28509 11471 28543
rect 12357 28509 12391 28543
rect 14105 28509 14139 28543
rect 16313 28509 16347 28543
rect 17325 28509 17359 28543
rect 18521 28509 18555 28543
rect 21465 28509 21499 28543
rect 21833 28509 21867 28543
rect 22661 28509 22695 28543
rect 23305 28509 23339 28543
rect 24685 28509 24719 28543
rect 27629 28509 27663 28543
rect 28457 28509 28491 28543
rect 29837 28509 29871 28543
rect 29989 28509 30023 28543
rect 30205 28509 30239 28543
rect 30849 28509 30883 28543
rect 31953 28509 31987 28543
rect 32689 28509 32723 28543
rect 34713 28509 34747 28543
rect 47685 28509 47719 28543
rect 14381 28441 14415 28475
rect 22477 28441 22511 28475
rect 26985 28441 27019 28475
rect 32965 28441 32999 28475
rect 11345 28373 11379 28407
rect 18613 28373 18647 28407
rect 22017 28373 22051 28407
rect 23489 28373 23523 28407
rect 28549 28373 28583 28407
rect 29653 28373 29687 28407
rect 31033 28373 31067 28407
rect 31769 28373 31803 28407
rect 11805 28169 11839 28203
rect 13185 28169 13219 28203
rect 15209 28169 15243 28203
rect 22569 28169 22603 28203
rect 27537 28169 27571 28203
rect 34069 28169 34103 28203
rect 11713 28101 11747 28135
rect 14105 28101 14139 28135
rect 14381 28101 14415 28135
rect 16037 28101 16071 28135
rect 16865 28101 16899 28135
rect 19257 28101 19291 28135
rect 31493 28101 31527 28135
rect 32597 28101 32631 28135
rect 10333 28033 10367 28067
rect 11897 28033 11931 28067
rect 12541 28033 12575 28067
rect 13369 28033 13403 28067
rect 14289 28033 14323 28067
rect 14473 28033 14507 28067
rect 15117 28033 15151 28067
rect 15945 28033 15979 28067
rect 18981 28033 19015 28067
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22385 28033 22419 28067
rect 26985 28033 27019 28067
rect 27353 28033 27387 28067
rect 31309 28033 31343 28067
rect 31585 28033 31619 28067
rect 32321 28033 32355 28067
rect 47593 28033 47627 28067
rect 12081 27965 12115 27999
rect 13553 27965 13587 27999
rect 13645 27965 13679 27999
rect 16681 27965 16715 27999
rect 17141 27965 17175 27999
rect 22109 27965 22143 27999
rect 22201 27965 22235 27999
rect 28549 27965 28583 27999
rect 28825 27965 28859 27999
rect 30297 27965 30331 27999
rect 11529 27897 11563 27931
rect 10517 27829 10551 27863
rect 12633 27829 12667 27863
rect 14657 27829 14691 27863
rect 20729 27829 20763 27863
rect 27353 27829 27387 27863
rect 31309 27829 31343 27863
rect 47685 27829 47719 27863
rect 10872 27625 10906 27659
rect 12357 27625 12391 27659
rect 31585 27625 31619 27659
rect 13461 27557 13495 27591
rect 21465 27557 21499 27591
rect 26525 27557 26559 27591
rect 29561 27557 29595 27591
rect 33609 27557 33643 27591
rect 10609 27489 10643 27523
rect 23213 27489 23247 27523
rect 30021 27489 30055 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 13369 27421 13403 27455
rect 14197 27421 14231 27455
rect 14381 27421 14415 27455
rect 20821 27421 20855 27455
rect 20969 27421 21003 27455
rect 21327 27421 21361 27455
rect 22845 27421 22879 27455
rect 23029 27421 23063 27455
rect 23121 27421 23155 27455
rect 23397 27421 23431 27455
rect 26341 27421 26375 27455
rect 29745 27421 29779 27455
rect 29837 27421 29871 27455
rect 30113 27421 30147 27455
rect 31769 27421 31803 27455
rect 31861 27421 31895 27455
rect 32045 27421 32079 27455
rect 32137 27421 32171 27455
rect 33517 27421 33551 27455
rect 14289 27353 14323 27387
rect 21097 27353 21131 27387
rect 21189 27353 21223 27387
rect 23581 27285 23615 27319
rect 11805 27081 11839 27115
rect 28365 27081 28399 27115
rect 11621 27013 11655 27047
rect 23121 27013 23155 27047
rect 30941 27013 30975 27047
rect 11529 26945 11563 26979
rect 11897 26945 11931 26979
rect 14105 26945 14139 26979
rect 20637 26945 20671 26979
rect 20729 26945 20763 26979
rect 21833 26945 21867 26979
rect 23305 26945 23339 26979
rect 23949 26945 23983 26979
rect 24133 26945 24167 26979
rect 25697 26945 25731 26979
rect 28181 26945 28215 26979
rect 31125 26945 31159 26979
rect 31217 26945 31251 26979
rect 11713 26877 11747 26911
rect 22109 26877 22143 26911
rect 25789 26877 25823 26911
rect 23489 26809 23523 26843
rect 26065 26809 26099 26843
rect 14197 26741 14231 26775
rect 20821 26741 20855 26775
rect 21005 26741 21039 26775
rect 23949 26741 23983 26775
rect 25881 26741 25915 26775
rect 30941 26741 30975 26775
rect 30941 26537 30975 26571
rect 32689 26537 32723 26571
rect 33149 26537 33183 26571
rect 33609 26537 33643 26571
rect 12265 26469 12299 26503
rect 15485 26469 15519 26503
rect 16589 26469 16623 26503
rect 21557 26469 21591 26503
rect 23305 26469 23339 26503
rect 29561 26469 29595 26503
rect 32229 26469 32263 26503
rect 14197 26401 14231 26435
rect 21428 26401 21462 26435
rect 21649 26401 21683 26435
rect 23397 26401 23431 26435
rect 24777 26401 24811 26435
rect 30205 26401 30239 26435
rect 32781 26401 32815 26435
rect 34069 26401 34103 26435
rect 10057 26333 10091 26367
rect 12081 26333 12115 26367
rect 14289 26333 14323 26367
rect 15117 26333 15151 26367
rect 15301 26333 15335 26367
rect 16589 26333 16623 26367
rect 16865 26333 16899 26367
rect 17325 26333 17359 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 20453 26333 20487 26367
rect 23121 26333 23155 26367
rect 24409 26333 24443 26367
rect 24593 26333 24627 26367
rect 26157 26333 26191 26367
rect 26249 26333 26283 26367
rect 26341 26333 26375 26367
rect 26525 26333 26559 26367
rect 27077 26333 27111 26367
rect 27169 26333 27203 26367
rect 28365 26333 28399 26367
rect 28549 26333 28583 26367
rect 28641 26333 28675 26367
rect 29929 26333 29963 26367
rect 31677 26333 31711 26367
rect 31861 26333 31895 26367
rect 32045 26333 32079 26367
rect 32965 26333 32999 26367
rect 33793 26333 33827 26367
rect 33977 26333 34011 26367
rect 47685 26333 47719 26367
rect 20637 26265 20671 26299
rect 20821 26265 20855 26299
rect 21281 26265 21315 26299
rect 22017 26265 22051 26299
rect 25881 26265 25915 26299
rect 28181 26265 28215 26299
rect 30021 26265 30055 26299
rect 30849 26265 30883 26299
rect 31953 26265 31987 26299
rect 32689 26265 32723 26299
rect 10241 26197 10275 26231
rect 14657 26197 14691 26231
rect 16773 26197 16807 26231
rect 17509 26197 17543 26231
rect 18153 26197 18187 26231
rect 22937 26197 22971 26231
rect 27353 26197 27387 26231
rect 18889 25993 18923 26027
rect 19901 25993 19935 26027
rect 27353 25993 27387 26027
rect 29837 25993 29871 26027
rect 31585 25993 31619 26027
rect 32229 25993 32263 26027
rect 33333 25993 33367 26027
rect 13553 25925 13587 25959
rect 16037 25925 16071 25959
rect 20453 25925 20487 25959
rect 26065 25925 26099 25959
rect 28365 25925 28399 25959
rect 10333 25857 10367 25891
rect 12725 25857 12759 25891
rect 16129 25857 16163 25891
rect 17141 25857 17175 25891
rect 19717 25857 19751 25891
rect 20729 25857 20763 25891
rect 20913 25857 20947 25891
rect 21189 25857 21223 25891
rect 25789 25857 25823 25891
rect 26985 25857 27019 25891
rect 27169 25857 27203 25891
rect 28549 25857 28583 25891
rect 28641 25857 28675 25891
rect 29745 25857 29779 25891
rect 30389 25857 30423 25891
rect 31217 25857 31251 25891
rect 31401 25857 31435 25891
rect 32137 25857 32171 25891
rect 32321 25857 32355 25891
rect 32965 25857 32999 25891
rect 33977 25857 34011 25891
rect 34161 25857 34195 25891
rect 34253 25857 34287 25891
rect 10425 25789 10459 25823
rect 12817 25789 12851 25823
rect 13277 25789 13311 25823
rect 15669 25789 15703 25823
rect 17417 25789 17451 25823
rect 19533 25789 19567 25823
rect 21005 25789 21039 25823
rect 22753 25789 22787 25823
rect 23029 25789 23063 25823
rect 24501 25789 24535 25823
rect 26157 25789 26191 25823
rect 26274 25789 26308 25823
rect 33057 25789 33091 25823
rect 20821 25721 20855 25755
rect 30573 25721 30607 25755
rect 10701 25653 10735 25687
rect 15025 25653 15059 25687
rect 15853 25653 15887 25687
rect 26433 25653 26467 25687
rect 28365 25653 28399 25687
rect 33793 25653 33827 25687
rect 47777 25653 47811 25687
rect 18429 25449 18463 25483
rect 19349 25449 19383 25483
rect 23029 25449 23063 25483
rect 24501 25449 24535 25483
rect 34161 25449 34195 25483
rect 15393 25381 15427 25415
rect 23397 25381 23431 25415
rect 29745 25381 29779 25415
rect 10241 25313 10275 25347
rect 10517 25313 10551 25347
rect 12265 25313 12299 25347
rect 16957 25313 16991 25347
rect 20269 25313 20303 25347
rect 32413 25313 32447 25347
rect 32689 25313 32723 25347
rect 46305 25313 46339 25347
rect 14749 25245 14783 25279
rect 15761 25245 15795 25279
rect 16681 25245 16715 25279
rect 19257 25245 19291 25279
rect 20453 25245 20487 25279
rect 20637 25245 20671 25279
rect 21189 25245 21223 25279
rect 21282 25245 21316 25279
rect 21557 25245 21591 25279
rect 21695 25245 21729 25279
rect 23029 25245 23063 25279
rect 23213 25245 23247 25279
rect 24409 25245 24443 25279
rect 25421 25245 25455 25279
rect 25605 25245 25639 25279
rect 25789 25245 25823 25279
rect 26617 25245 26651 25279
rect 26709 25245 26743 25279
rect 26893 25245 26927 25279
rect 26985 25245 27019 25279
rect 29561 25245 29595 25279
rect 30757 25245 30791 25279
rect 31125 25245 31159 25279
rect 1869 25177 1903 25211
rect 14381 25177 14415 25211
rect 14565 25177 14599 25211
rect 15669 25177 15703 25211
rect 21465 25177 21499 25211
rect 25697 25177 25731 25211
rect 30941 25177 30975 25211
rect 31033 25177 31067 25211
rect 35173 25177 35207 25211
rect 46489 25177 46523 25211
rect 48145 25177 48179 25211
rect 1961 25109 1995 25143
rect 14657 25109 14691 25143
rect 14933 25109 14967 25143
rect 15577 25109 15611 25143
rect 15945 25109 15979 25143
rect 21833 25109 21867 25143
rect 25973 25109 26007 25143
rect 26433 25109 26467 25143
rect 31309 25109 31343 25143
rect 35265 25109 35299 25143
rect 14933 24905 14967 24939
rect 15485 24905 15519 24939
rect 17049 24905 17083 24939
rect 21281 24905 21315 24939
rect 26433 24905 26467 24939
rect 16865 24837 16899 24871
rect 16957 24837 16991 24871
rect 31033 24837 31067 24871
rect 10793 24769 10827 24803
rect 10977 24769 11011 24803
rect 11529 24769 11563 24803
rect 11621 24769 11655 24803
rect 14749 24769 14783 24803
rect 15669 24769 15703 24803
rect 15853 24769 15887 24803
rect 15945 24769 15979 24803
rect 16681 24769 16715 24803
rect 18245 24769 18279 24803
rect 18337 24769 18371 24803
rect 20913 24769 20947 24803
rect 21833 24769 21867 24803
rect 26985 24769 27019 24803
rect 28089 24769 28123 24803
rect 30573 24769 30607 24803
rect 31217 24769 31251 24803
rect 32229 24769 32263 24803
rect 32413 24769 32447 24803
rect 32873 24769 32907 24803
rect 32965 24769 32999 24803
rect 35173 24769 35207 24803
rect 39957 24769 39991 24803
rect 47593 24769 47627 24803
rect 47685 24769 47719 24803
rect 14565 24701 14599 24735
rect 17233 24701 17267 24735
rect 21005 24701 21039 24735
rect 22109 24701 22143 24735
rect 24685 24701 24719 24735
rect 24961 24701 24995 24735
rect 27077 24701 27111 24735
rect 28365 24701 28399 24735
rect 29837 24701 29871 24735
rect 31401 24701 31435 24735
rect 35449 24701 35483 24735
rect 45201 24701 45235 24735
rect 45385 24701 45419 24735
rect 46765 24701 46799 24735
rect 10793 24565 10827 24599
rect 23581 24565 23615 24599
rect 30389 24565 30423 24599
rect 40049 24565 40083 24599
rect 16589 24361 16623 24395
rect 23305 24361 23339 24395
rect 26893 24361 26927 24395
rect 29653 24361 29687 24395
rect 31014 24361 31048 24395
rect 32505 24361 32539 24395
rect 45109 24361 45143 24395
rect 19441 24293 19475 24327
rect 10609 24225 10643 24259
rect 25145 24225 25179 24259
rect 25421 24225 25455 24259
rect 30757 24225 30791 24259
rect 34161 24225 34195 24259
rect 36921 24225 36955 24259
rect 40049 24225 40083 24259
rect 40325 24225 40359 24259
rect 46949 24225 46983 24259
rect 10333 24157 10367 24191
rect 12541 24157 12575 24191
rect 16497 24157 16531 24191
rect 17693 24157 17727 24191
rect 19257 24157 19291 24191
rect 19993 24157 20027 24191
rect 23213 24157 23247 24191
rect 29561 24157 29595 24191
rect 35081 24157 35115 24191
rect 39865 24157 39899 24191
rect 45017 24157 45051 24191
rect 45661 24157 45695 24191
rect 46305 24157 46339 24191
rect 12633 24089 12667 24123
rect 33977 24089 34011 24123
rect 35265 24089 35299 24123
rect 45753 24089 45787 24123
rect 46489 24089 46523 24123
rect 12081 24021 12115 24055
rect 17877 24021 17911 24055
rect 20085 24021 20119 24055
rect 17601 23817 17635 23851
rect 23765 23817 23799 23851
rect 25973 23817 26007 23851
rect 32229 23817 32263 23851
rect 34529 23817 34563 23851
rect 41061 23817 41095 23851
rect 10425 23749 10459 23783
rect 14197 23749 14231 23783
rect 19625 23749 19659 23783
rect 1869 23681 1903 23715
rect 10149 23681 10183 23715
rect 14933 23681 14967 23715
rect 15577 23681 15611 23715
rect 17417 23681 17451 23715
rect 18429 23681 18463 23715
rect 23581 23681 23615 23715
rect 24317 23681 24351 23715
rect 25881 23681 25915 23715
rect 32137 23681 32171 23715
rect 34437 23681 34471 23715
rect 35265 23681 35299 23715
rect 39681 23681 39715 23715
rect 40693 23681 40727 23715
rect 43269 23681 43303 23715
rect 43453 23681 43487 23715
rect 44097 23681 44131 23715
rect 44281 23681 44315 23715
rect 45753 23681 45787 23715
rect 47593 23681 47627 23715
rect 11805 23613 11839 23647
rect 11989 23613 12023 23647
rect 13185 23613 13219 23647
rect 15117 23613 15151 23647
rect 18153 23613 18187 23647
rect 19441 23613 19475 23647
rect 20821 23613 20855 23647
rect 36277 23613 36311 23647
rect 39589 23613 39623 23647
rect 40601 23613 40635 23647
rect 43637 23613 43671 23647
rect 46213 23613 46247 23647
rect 46489 23613 46523 23647
rect 2053 23545 2087 23579
rect 40049 23545 40083 23579
rect 14289 23477 14323 23511
rect 15669 23477 15703 23511
rect 24501 23477 24535 23511
rect 44097 23477 44131 23511
rect 45569 23477 45603 23511
rect 47685 23477 47719 23511
rect 11345 23273 11379 23307
rect 12173 23273 12207 23307
rect 13093 23273 13127 23307
rect 13277 23273 13311 23307
rect 20637 23273 20671 23307
rect 25697 23273 25731 23307
rect 42533 23205 42567 23239
rect 14105 23137 14139 23171
rect 15761 23137 15795 23171
rect 16405 23137 16439 23171
rect 30665 23137 30699 23171
rect 35725 23137 35759 23171
rect 40509 23137 40543 23171
rect 43637 23137 43671 23171
rect 46305 23137 46339 23171
rect 46489 23137 46523 23171
rect 48145 23137 48179 23171
rect 9873 23069 9907 23103
rect 10701 23069 10735 23103
rect 11621 23069 11655 23103
rect 12081 23069 12115 23103
rect 19349 23069 19383 23103
rect 20453 23069 20487 23103
rect 22845 23069 22879 23103
rect 23489 23069 23523 23103
rect 25513 23069 25547 23103
rect 28273 23069 28307 23103
rect 30205 23069 30239 23103
rect 33701 23069 33735 23103
rect 35173 23069 35207 23103
rect 39865 23069 39899 23103
rect 42257 23069 42291 23103
rect 43821 23069 43855 23103
rect 45845 23069 45879 23103
rect 11345 23001 11379 23035
rect 12909 23001 12943 23035
rect 14289 23001 14323 23035
rect 16681 23001 16715 23035
rect 19901 23001 19935 23035
rect 30389 23001 30423 23035
rect 40049 23001 40083 23035
rect 44465 23001 44499 23035
rect 9873 22933 9907 22967
rect 10793 22933 10827 22967
rect 11529 22933 11563 22967
rect 13109 22933 13143 22967
rect 18153 22933 18187 22967
rect 22937 22933 22971 22967
rect 23581 22933 23615 22967
rect 28365 22933 28399 22967
rect 33793 22933 33827 22967
rect 45661 22933 45695 22967
rect 10885 22729 10919 22763
rect 11897 22729 11931 22763
rect 13553 22729 13587 22763
rect 14315 22729 14349 22763
rect 32229 22729 32263 22763
rect 39497 22729 39531 22763
rect 47961 22729 47995 22763
rect 11529 22661 11563 22695
rect 11745 22661 11779 22695
rect 14105 22661 14139 22695
rect 21925 22661 21959 22695
rect 23489 22661 23523 22695
rect 25145 22661 25179 22695
rect 33793 22661 33827 22695
rect 41889 22661 41923 22695
rect 43361 22661 43395 22695
rect 45385 22661 45419 22695
rect 47777 22661 47811 22695
rect 8217 22593 8251 22627
rect 10701 22593 10735 22627
rect 12541 22593 12575 22627
rect 13369 22593 13403 22627
rect 15117 22593 15151 22627
rect 16865 22593 16899 22627
rect 21833 22593 21867 22627
rect 25973 22593 26007 22627
rect 27077 22593 27111 22627
rect 27905 22593 27939 22627
rect 28733 22593 28767 22627
rect 32137 22593 32171 22627
rect 39405 22593 39439 22627
rect 40049 22593 40083 22627
rect 42441 22593 42475 22627
rect 43545 22593 43579 22627
rect 43637 22593 43671 22627
rect 44097 22593 44131 22627
rect 44281 22593 44315 22627
rect 47593 22593 47627 22627
rect 47869 22593 47903 22627
rect 8401 22525 8435 22559
rect 8677 22525 8711 22559
rect 15209 22525 15243 22559
rect 15485 22525 15519 22559
rect 17049 22525 17083 22559
rect 18705 22525 18739 22559
rect 19257 22525 19291 22559
rect 19533 22525 19567 22559
rect 21281 22525 21315 22559
rect 23305 22525 23339 22559
rect 27997 22525 28031 22559
rect 28273 22525 28307 22559
rect 29009 22525 29043 22559
rect 33609 22525 33643 22559
rect 35449 22525 35483 22559
rect 40233 22525 40267 22559
rect 42717 22525 42751 22559
rect 45201 22525 45235 22559
rect 46857 22525 46891 22559
rect 43361 22457 43395 22491
rect 44097 22457 44131 22491
rect 11713 22389 11747 22423
rect 12725 22389 12759 22423
rect 14289 22389 14323 22423
rect 14473 22389 14507 22423
rect 25973 22389 26007 22423
rect 27169 22389 27203 22423
rect 30481 22389 30515 22423
rect 48145 22389 48179 22423
rect 8309 22185 8343 22219
rect 9768 22185 9802 22219
rect 11713 22185 11747 22219
rect 15117 22185 15151 22219
rect 16957 22185 16991 22219
rect 40141 22185 40175 22219
rect 40969 22185 41003 22219
rect 43269 22185 43303 22219
rect 11253 22117 11287 22151
rect 12265 22117 12299 22151
rect 20453 22117 20487 22151
rect 28917 22117 28951 22151
rect 9505 22049 9539 22083
rect 19901 22049 19935 22083
rect 21261 22049 21295 22083
rect 26065 22049 26099 22083
rect 29653 22049 29687 22083
rect 32597 22049 32631 22083
rect 8217 21981 8251 22015
rect 11894 21981 11928 22015
rect 12357 21981 12391 22015
rect 14105 21981 14139 22015
rect 15025 21981 15059 22015
rect 16037 21981 16071 22015
rect 16865 21981 16899 22015
rect 17785 21981 17819 22015
rect 19349 21981 19383 22015
rect 20453 21981 20487 22015
rect 20729 21981 20763 22015
rect 21465 21981 21499 22015
rect 22017 21981 22051 22015
rect 22201 21981 22235 22015
rect 22845 21981 22879 22015
rect 23581 21981 23615 22015
rect 25421 21981 25455 22015
rect 28733 21981 28767 22015
rect 29561 21981 29595 22015
rect 34161 21981 34195 22015
rect 40049 21981 40083 22015
rect 41153 21981 41187 22015
rect 43177 21981 43211 22015
rect 43361 21981 43395 22015
rect 45017 21981 45051 22015
rect 45201 21981 45235 22015
rect 45661 21981 45695 22015
rect 48145 21981 48179 22015
rect 12909 21913 12943 21947
rect 18337 21913 18371 21947
rect 21189 21913 21223 21947
rect 26341 21913 26375 21947
rect 28365 21913 28399 21947
rect 28549 21913 28583 21947
rect 32321 21913 32355 21947
rect 32413 21913 32447 21947
rect 34805 21913 34839 21947
rect 34897 21913 34931 21947
rect 35817 21913 35851 21947
rect 43913 21913 43947 21947
rect 44097 21913 44131 21947
rect 45845 21913 45879 21947
rect 47501 21913 47535 21947
rect 11897 21845 11931 21879
rect 13001 21845 13035 21879
rect 14289 21845 14323 21879
rect 16221 21845 16255 21879
rect 20637 21845 20671 21879
rect 21373 21845 21407 21879
rect 22109 21845 22143 21879
rect 23029 21845 23063 21879
rect 23673 21845 23707 21879
rect 25513 21845 25547 21879
rect 27813 21845 27847 21879
rect 28641 21845 28675 21879
rect 33977 21845 34011 21879
rect 40509 21845 40543 21879
rect 44281 21845 44315 21879
rect 45201 21845 45235 21879
rect 47961 21845 47995 21879
rect 11897 21641 11931 21675
rect 12659 21641 12693 21675
rect 16037 21641 16071 21675
rect 19533 21641 19567 21675
rect 20177 21641 20211 21675
rect 21005 21641 21039 21675
rect 33057 21641 33091 21675
rect 33977 21641 34011 21675
rect 48145 21641 48179 21675
rect 12449 21573 12483 21607
rect 20729 21573 20763 21607
rect 22569 21573 22603 21607
rect 27997 21573 28031 21607
rect 28197 21573 28231 21607
rect 30665 21573 30699 21607
rect 31585 21573 31619 21607
rect 35081 21573 35115 21607
rect 45017 21573 45051 21607
rect 8309 21505 8343 21539
rect 11713 21505 11747 21539
rect 11989 21505 12023 21539
rect 13737 21505 13771 21539
rect 14933 21505 14967 21539
rect 15945 21505 15979 21539
rect 17325 21505 17359 21539
rect 18153 21505 18187 21539
rect 19441 21505 19475 21539
rect 20085 21505 20119 21539
rect 20269 21505 20303 21539
rect 20913 21505 20947 21539
rect 21097 21505 21131 21539
rect 27169 21505 27203 21539
rect 28825 21505 28859 21539
rect 29009 21505 29043 21539
rect 29101 21527 29135 21561
rect 29561 21505 29595 21539
rect 29745 21505 29779 21539
rect 32137 21505 32171 21539
rect 33241 21505 33275 21539
rect 34437 21505 34471 21539
rect 39957 21505 39991 21539
rect 40141 21505 40175 21539
rect 43177 21505 43211 21539
rect 43361 21505 43395 21539
rect 44281 21505 44315 21539
rect 46213 21505 46247 21539
rect 47593 21505 47627 21539
rect 8493 21437 8527 21471
rect 9137 21437 9171 21471
rect 17417 21437 17451 21471
rect 18429 21437 18463 21471
rect 22293 21437 22327 21471
rect 24041 21437 24075 21471
rect 24501 21437 24535 21471
rect 24777 21437 24811 21471
rect 27261 21437 27295 21471
rect 30573 21437 30607 21471
rect 32597 21437 32631 21471
rect 34989 21437 35023 21471
rect 35817 21437 35851 21471
rect 46489 21437 46523 21471
rect 47869 21437 47903 21471
rect 12817 21369 12851 21403
rect 27537 21369 27571 21403
rect 28365 21369 28399 21403
rect 28825 21369 28859 21403
rect 11529 21301 11563 21335
rect 12633 21301 12667 21335
rect 13829 21301 13863 21335
rect 15117 21301 15151 21335
rect 17693 21301 17727 21335
rect 21281 21301 21315 21335
rect 26249 21301 26283 21335
rect 28181 21301 28215 21335
rect 29561 21301 29595 21335
rect 32413 21301 32447 21335
rect 33609 21301 33643 21335
rect 34161 21301 34195 21335
rect 40049 21301 40083 21335
rect 43177 21301 43211 21335
rect 47685 21301 47719 21335
rect 9045 21097 9079 21131
rect 20821 21097 20855 21131
rect 21005 21097 21039 21131
rect 22385 21097 22419 21131
rect 25329 21097 25363 21131
rect 11529 21029 11563 21063
rect 43177 21029 43211 21063
rect 11713 20961 11747 20995
rect 14289 20961 14323 20995
rect 14565 20961 14599 20995
rect 16405 20961 16439 20995
rect 17969 20961 18003 20995
rect 21465 20961 21499 20995
rect 21833 20961 21867 20995
rect 24869 20961 24903 20995
rect 43361 20961 43395 20995
rect 43637 20961 43671 20995
rect 46305 20961 46339 20995
rect 48145 20961 48179 20995
rect 8953 20893 8987 20927
rect 10793 20893 10827 20927
rect 14105 20893 14139 20927
rect 19441 20893 19475 20927
rect 21649 20893 21683 20927
rect 22569 20893 22603 20927
rect 23121 20893 23155 20927
rect 24961 20893 24995 20927
rect 28273 20893 28307 20927
rect 29561 20893 29595 20927
rect 30849 20893 30883 20927
rect 33149 20893 33183 20927
rect 42533 20893 42567 20927
rect 42717 20893 42751 20927
rect 43453 20893 43487 20927
rect 43545 20893 43579 20927
rect 44189 20893 44223 20927
rect 44373 20893 44407 20927
rect 45477 20893 45511 20927
rect 45661 20893 45695 20927
rect 11253 20825 11287 20859
rect 16589 20825 16623 20859
rect 20637 20825 20671 20859
rect 20853 20825 20887 20859
rect 28457 20825 28491 20859
rect 31033 20825 31067 20859
rect 32689 20825 32723 20859
rect 46489 20825 46523 20859
rect 10609 20757 10643 20791
rect 19625 20757 19659 20791
rect 23305 20757 23339 20791
rect 29653 20757 29687 20791
rect 33241 20757 33275 20791
rect 42717 20757 42751 20791
rect 44281 20757 44315 20791
rect 45845 20757 45879 20791
rect 16773 20553 16807 20587
rect 23305 20553 23339 20587
rect 45661 20553 45695 20587
rect 48053 20553 48087 20587
rect 11805 20485 11839 20519
rect 18245 20485 18279 20519
rect 24133 20485 24167 20519
rect 28733 20485 28767 20519
rect 32965 20485 32999 20519
rect 44925 20485 44959 20519
rect 16681 20417 16715 20451
rect 17325 20417 17359 20451
rect 20453 20417 20487 20451
rect 21833 20417 21867 20451
rect 23121 20417 23155 20451
rect 23857 20417 23891 20451
rect 28457 20417 28491 20451
rect 32137 20417 32171 20451
rect 43085 20417 43119 20451
rect 43453 20417 43487 20451
rect 44557 20417 44591 20451
rect 44741 20417 44775 20451
rect 45569 20417 45603 20451
rect 46213 20417 46247 20451
rect 47593 20417 47627 20451
rect 11529 20349 11563 20383
rect 13277 20349 13311 20383
rect 14289 20349 14323 20383
rect 14473 20349 14507 20383
rect 16129 20349 16163 20383
rect 17969 20349 18003 20383
rect 20545 20349 20579 20383
rect 30205 20349 30239 20383
rect 32781 20349 32815 20383
rect 34437 20349 34471 20383
rect 44005 20349 44039 20383
rect 46489 20349 46523 20383
rect 19717 20281 19751 20315
rect 17417 20213 17451 20247
rect 20821 20213 20855 20247
rect 21925 20213 21959 20247
rect 32229 20213 32263 20247
rect 47685 20213 47719 20247
rect 28825 20009 28859 20043
rect 30757 20009 30791 20043
rect 42993 20009 43027 20043
rect 43821 20009 43855 20043
rect 48053 20009 48087 20043
rect 10701 19941 10735 19975
rect 12081 19941 12115 19975
rect 15485 19941 15519 19975
rect 23765 19941 23799 19975
rect 43545 19941 43579 19975
rect 16865 19873 16899 19907
rect 17049 19873 17083 19907
rect 19625 19873 19659 19907
rect 19901 19873 19935 19907
rect 31769 19873 31803 19907
rect 45569 19873 45603 19907
rect 45753 19873 45787 19907
rect 46949 19873 46983 19907
rect 2053 19805 2087 19839
rect 10701 19805 10735 19839
rect 11253 19805 11287 19839
rect 11989 19805 12023 19839
rect 12817 19805 12851 19839
rect 14381 19805 14415 19839
rect 15393 19805 15427 19839
rect 22017 19805 22051 19839
rect 26801 19805 26835 19839
rect 28641 19805 28675 19839
rect 30665 19805 30699 19839
rect 31309 19805 31343 19839
rect 42901 19805 42935 19839
rect 43085 19805 43119 19839
rect 43821 19805 43855 19839
rect 44005 19805 44039 19839
rect 18705 19737 18739 19771
rect 22293 19737 22327 19771
rect 31493 19737 31527 19771
rect 11437 19669 11471 19703
rect 13001 19669 13035 19703
rect 14473 19669 14507 19703
rect 21373 19669 21407 19703
rect 26617 19669 26651 19703
rect 14657 19465 14691 19499
rect 18429 19465 18463 19499
rect 19073 19465 19107 19499
rect 22937 19465 22971 19499
rect 26341 19465 26375 19499
rect 31125 19465 31159 19499
rect 43453 19465 43487 19499
rect 44281 19465 44315 19499
rect 46765 19465 46799 19499
rect 15117 19397 15151 19431
rect 15301 19397 15335 19431
rect 46673 19397 46707 19431
rect 46949 19397 46983 19431
rect 1777 19329 1811 19363
rect 10885 19329 10919 19363
rect 11529 19329 11563 19363
rect 12909 19329 12943 19363
rect 15393 19329 15427 19363
rect 15485 19329 15519 19363
rect 18337 19329 18371 19363
rect 18981 19329 19015 19363
rect 22845 19329 22879 19363
rect 26157 19329 26191 19363
rect 26985 19329 27019 19363
rect 28181 19329 28215 19363
rect 28273 19329 28307 19363
rect 28825 19329 28859 19363
rect 31309 19329 31343 19363
rect 32137 19329 32171 19363
rect 43361 19329 43395 19363
rect 43545 19329 43579 19363
rect 44097 19329 44131 19363
rect 44281 19329 44315 19363
rect 46581 19329 46615 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 13185 19261 13219 19295
rect 15669 19261 15703 19295
rect 25973 19261 26007 19295
rect 46397 19193 46431 19227
rect 10701 19125 10735 19159
rect 11621 19125 11655 19159
rect 26985 19125 27019 19159
rect 28917 19125 28951 19159
rect 32229 19125 32263 19159
rect 47777 19125 47811 19159
rect 2237 18921 2271 18955
rect 33793 18921 33827 18955
rect 12909 18853 12943 18887
rect 10425 18785 10459 18819
rect 15025 18785 15059 18819
rect 25881 18785 25915 18819
rect 26801 18785 26835 18819
rect 27077 18785 27111 18819
rect 31401 18785 31435 18819
rect 32321 18785 32355 18819
rect 46305 18785 46339 18819
rect 48145 18785 48179 18819
rect 2145 18717 2179 18751
rect 13093 18717 13127 18751
rect 13369 18717 13403 18751
rect 13553 18717 13587 18751
rect 14657 18717 14691 18751
rect 19441 18717 19475 18751
rect 23213 18717 23247 18751
rect 24409 18717 24443 18751
rect 25973 18717 26007 18751
rect 29929 18717 29963 18751
rect 30113 18717 30147 18751
rect 31217 18717 31251 18751
rect 33517 18717 33551 18751
rect 45845 18717 45879 18751
rect 10701 18649 10735 18683
rect 14473 18649 14507 18683
rect 22017 18649 22051 18683
rect 46489 18649 46523 18683
rect 12173 18581 12207 18615
rect 14749 18581 14783 18615
rect 14841 18581 14875 18615
rect 19533 18581 19567 18615
rect 22109 18581 22143 18615
rect 23397 18581 23431 18615
rect 24593 18581 24627 18615
rect 26341 18581 26375 18615
rect 28549 18581 28583 18615
rect 30113 18581 30147 18615
rect 33977 18581 34011 18615
rect 45661 18581 45695 18615
rect 47685 18377 47719 18411
rect 19625 18309 19659 18343
rect 25605 18309 25639 18343
rect 25973 18309 26007 18343
rect 27261 18309 27295 18343
rect 30021 18309 30055 18343
rect 30205 18309 30239 18343
rect 31217 18309 31251 18343
rect 32505 18309 32539 18343
rect 1409 18241 1443 18275
rect 10609 18241 10643 18275
rect 13277 18241 13311 18275
rect 13921 18241 13955 18275
rect 14105 18241 14139 18275
rect 14749 18241 14783 18275
rect 15945 18241 15979 18275
rect 16773 18241 16807 18275
rect 16957 18241 16991 18275
rect 18797 18241 18831 18275
rect 21833 18241 21867 18275
rect 23305 18241 23339 18275
rect 24225 18241 24259 18275
rect 24777 18241 24811 18275
rect 25789 18241 25823 18275
rect 30389 18241 30423 18275
rect 31033 18241 31067 18275
rect 34805 18241 34839 18275
rect 43361 18241 43395 18275
rect 46029 18241 46063 18275
rect 46397 18241 46431 18275
rect 46765 18241 46799 18275
rect 47041 18241 47075 18275
rect 47593 18241 47627 18275
rect 10517 18173 10551 18207
rect 10977 18173 11011 18207
rect 14657 18173 14691 18207
rect 19441 18173 19475 18207
rect 21281 18173 21315 18207
rect 22109 18173 22143 18207
rect 23949 18173 23983 18207
rect 24041 18173 24075 18207
rect 24133 18173 24167 18207
rect 26985 18173 27019 18207
rect 30849 18173 30883 18207
rect 32321 18173 32355 18207
rect 34069 18173 34103 18207
rect 43545 18173 43579 18207
rect 45201 18173 45235 18207
rect 1593 18105 1627 18139
rect 13369 18105 13403 18139
rect 17141 18105 17175 18139
rect 28733 18105 28767 18139
rect 13921 18037 13955 18071
rect 15117 18037 15151 18071
rect 16037 18037 16071 18071
rect 18797 18037 18831 18071
rect 23121 18037 23155 18071
rect 23765 18037 23799 18071
rect 24869 18037 24903 18071
rect 34621 18037 34655 18071
rect 46305 18037 46339 18071
rect 14565 17833 14599 17867
rect 14749 17833 14783 17867
rect 16957 17833 16991 17867
rect 22109 17833 22143 17867
rect 25605 17833 25639 17867
rect 26525 17833 26559 17867
rect 43453 17833 43487 17867
rect 45661 17833 45695 17867
rect 24685 17765 24719 17799
rect 35909 17765 35943 17799
rect 15209 17697 15243 17731
rect 15485 17697 15519 17731
rect 18429 17697 18463 17731
rect 18705 17697 18739 17731
rect 19533 17697 19567 17731
rect 30297 17697 30331 17731
rect 30573 17697 30607 17731
rect 32229 17697 32263 17731
rect 32413 17697 32447 17731
rect 45385 17697 45419 17731
rect 46305 17697 46339 17731
rect 13185 17629 13219 17663
rect 18337 17629 18371 17663
rect 19257 17629 19291 17663
rect 21741 17629 21775 17663
rect 22753 17629 22787 17663
rect 23305 17629 23339 17663
rect 23489 17629 23523 17663
rect 25513 17629 25547 17663
rect 25697 17629 25731 17663
rect 26525 17629 26559 17663
rect 30205 17629 30239 17663
rect 35173 17629 35207 17663
rect 35357 17629 35391 17663
rect 35449 17629 35483 17663
rect 43361 17629 43395 17663
rect 44281 17629 44315 17663
rect 44465 17629 44499 17663
rect 45477 17629 45511 17663
rect 14381 17561 14415 17595
rect 21557 17561 21591 17595
rect 21925 17561 21959 17595
rect 23581 17561 23615 17595
rect 23857 17561 23891 17595
rect 24409 17561 24443 17595
rect 34069 17561 34103 17595
rect 34805 17561 34839 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 13277 17493 13311 17527
rect 14591 17493 14625 17527
rect 21005 17493 21039 17527
rect 21833 17493 21867 17527
rect 22753 17493 22787 17527
rect 23673 17493 23707 17527
rect 24869 17493 24903 17527
rect 44373 17493 44407 17527
rect 45017 17493 45051 17527
rect 30573 17289 30607 17323
rect 47961 17289 47995 17323
rect 13737 17221 13771 17255
rect 15761 17221 15795 17255
rect 20361 17221 20395 17255
rect 22201 17221 22235 17255
rect 23489 17221 23523 17255
rect 29837 17221 29871 17255
rect 35081 17221 35115 17255
rect 44465 17221 44499 17255
rect 45385 17221 45419 17255
rect 47777 17221 47811 17255
rect 11989 17153 12023 17187
rect 13461 17153 13495 17187
rect 15669 17153 15703 17187
rect 20269 17153 20303 17187
rect 22017 17153 22051 17187
rect 22109 17153 22143 17187
rect 23213 17153 23247 17187
rect 28089 17153 28123 17187
rect 28273 17153 28307 17187
rect 28733 17153 28767 17187
rect 29653 17153 29687 17187
rect 30021 17153 30055 17187
rect 30481 17153 30515 17187
rect 30665 17153 30699 17187
rect 43729 17153 43763 17187
rect 45201 17153 45235 17187
rect 47593 17153 47627 17187
rect 15209 17085 15243 17119
rect 16773 17085 16807 17119
rect 16957 17085 16991 17119
rect 18613 17085 18647 17119
rect 24961 17085 24995 17119
rect 29009 17085 29043 17119
rect 29101 17085 29135 17119
rect 34897 17085 34931 17119
rect 36737 17085 36771 17119
rect 46765 17085 46799 17119
rect 21833 17017 21867 17051
rect 28825 17017 28859 17051
rect 2053 16949 2087 16983
rect 12081 16949 12115 16983
rect 22385 16949 22419 16983
rect 28089 16949 28123 16983
rect 29193 16949 29227 16983
rect 14565 16745 14599 16779
rect 17049 16745 17083 16779
rect 22477 16745 22511 16779
rect 45753 16745 45787 16779
rect 22661 16677 22695 16711
rect 28457 16677 28491 16711
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 11713 16609 11747 16643
rect 11897 16609 11931 16643
rect 29745 16609 29779 16643
rect 30665 16609 30699 16643
rect 46305 16609 46339 16643
rect 11069 16551 11103 16585
rect 14565 16541 14599 16575
rect 14841 16541 14875 16575
rect 16957 16541 16991 16575
rect 21649 16541 21683 16575
rect 21833 16541 21867 16575
rect 24409 16541 24443 16575
rect 27169 16541 27203 16575
rect 27353 16541 27387 16575
rect 27813 16541 27847 16575
rect 27997 16541 28031 16575
rect 29837 16541 29871 16575
rect 45661 16541 45695 16575
rect 45845 16541 45879 16575
rect 1593 16473 1627 16507
rect 13553 16473 13587 16507
rect 22293 16473 22327 16507
rect 22509 16473 22543 16507
rect 28641 16473 28675 16507
rect 29009 16473 29043 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 11161 16405 11195 16439
rect 14749 16405 14783 16439
rect 21741 16405 21775 16439
rect 24501 16405 24535 16439
rect 27353 16405 27387 16439
rect 27997 16405 28031 16439
rect 28733 16405 28767 16439
rect 28825 16405 28859 16439
rect 2145 16201 2179 16235
rect 19901 16201 19935 16235
rect 22293 16201 22327 16235
rect 25605 16201 25639 16235
rect 27261 16201 27295 16235
rect 28549 16201 28583 16235
rect 29469 16201 29503 16235
rect 46949 16201 46983 16235
rect 47685 16201 47719 16235
rect 11713 16133 11747 16167
rect 19533 16133 19567 16167
rect 19733 16133 19767 16167
rect 22109 16133 22143 16167
rect 43913 16133 43947 16167
rect 44649 16133 44683 16167
rect 2053 16065 2087 16099
rect 11529 16065 11563 16099
rect 15117 16065 15151 16099
rect 16865 16065 16899 16099
rect 17417 16065 17451 16099
rect 18889 16065 18923 16099
rect 19073 16065 19107 16099
rect 20545 16065 20579 16099
rect 22385 16065 22419 16099
rect 23029 16065 23063 16099
rect 23857 16065 23891 16099
rect 27169 16065 27203 16099
rect 27353 16065 27387 16099
rect 28457 16065 28491 16099
rect 29285 16065 29319 16099
rect 43821 16065 43855 16099
rect 44465 16065 44499 16099
rect 46857 16065 46891 16099
rect 47593 16065 47627 16099
rect 12449 15997 12483 16031
rect 23121 15997 23155 16031
rect 24133 15997 24167 16031
rect 29101 15997 29135 16031
rect 46121 15997 46155 16031
rect 22109 15929 22143 15963
rect 23397 15929 23431 15963
rect 15209 15861 15243 15895
rect 16865 15861 16899 15895
rect 17509 15861 17543 15895
rect 18981 15861 19015 15895
rect 19717 15861 19751 15895
rect 20637 15861 20671 15895
rect 24777 15657 24811 15691
rect 47685 15657 47719 15691
rect 18613 15589 18647 15623
rect 14565 15521 14599 15555
rect 16865 15521 16899 15555
rect 19349 15521 19383 15555
rect 21557 15521 21591 15555
rect 2053 15453 2087 15487
rect 19441 15453 19475 15487
rect 20545 15453 20579 15487
rect 20821 15453 20855 15487
rect 21281 15453 21315 15487
rect 24685 15453 24719 15487
rect 43545 15453 43579 15487
rect 14841 15385 14875 15419
rect 17141 15385 17175 15419
rect 16313 15317 16347 15351
rect 19809 15317 19843 15351
rect 23029 15317 23063 15351
rect 43637 15317 43671 15351
rect 15577 15113 15611 15147
rect 17325 15113 17359 15147
rect 18797 15113 18831 15147
rect 22385 15113 22419 15147
rect 18429 15045 18463 15079
rect 18645 15045 18679 15079
rect 19533 15045 19567 15079
rect 43821 15045 43855 15079
rect 1777 14977 1811 15011
rect 14289 14977 14323 15011
rect 15485 14977 15519 15011
rect 17509 14977 17543 15011
rect 17785 14977 17819 15011
rect 17969 14977 18003 15011
rect 22293 14977 22327 15011
rect 43637 14977 43671 15011
rect 47777 14977 47811 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 14381 14909 14415 14943
rect 14657 14909 14691 14943
rect 19257 14909 19291 14943
rect 45293 14909 45327 14943
rect 18613 14773 18647 14807
rect 21005 14773 21039 14807
rect 2237 14569 2271 14603
rect 18613 14569 18647 14603
rect 19257 14433 19291 14467
rect 20729 14433 20763 14467
rect 21833 14433 21867 14467
rect 23397 14433 23431 14467
rect 2145 14365 2179 14399
rect 16681 14365 16715 14399
rect 17785 14365 17819 14399
rect 18613 14365 18647 14399
rect 47225 14365 47259 14399
rect 17877 14297 17911 14331
rect 19441 14297 19475 14331
rect 22017 14297 22051 14331
rect 16773 14229 16807 14263
rect 47317 14229 47351 14263
rect 22109 14025 22143 14059
rect 16865 13957 16899 13991
rect 16681 13889 16715 13923
rect 19441 13889 19475 13923
rect 22017 13889 22051 13923
rect 18521 13821 18555 13855
rect 19625 13821 19659 13855
rect 21281 13821 21315 13855
rect 47777 13685 47811 13719
rect 19349 13481 19383 13515
rect 16773 13345 16807 13379
rect 46305 13345 46339 13379
rect 15669 13277 15703 13311
rect 16313 13277 16347 13311
rect 19257 13277 19291 13311
rect 15761 13209 15795 13243
rect 16497 13209 16531 13243
rect 46489 13209 46523 13243
rect 48145 13209 48179 13243
rect 1409 12801 1443 12835
rect 21833 12801 21867 12835
rect 22017 12733 22051 12767
rect 22293 12733 22327 12767
rect 1593 12597 1627 12631
rect 21741 12393 21775 12427
rect 21649 12189 21683 12223
rect 46765 12189 46799 12223
rect 46857 12053 46891 12087
rect 47777 11509 47811 11543
rect 46305 11169 46339 11203
rect 46489 11169 46523 11203
rect 48145 11033 48179 11067
rect 47593 10625 47627 10659
rect 47041 10421 47075 10455
rect 47685 10421 47719 10455
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 47869 9537 47903 9571
rect 48053 9401 48087 9435
rect 47777 8857 47811 8891
rect 47869 8789 47903 8823
rect 48145 8449 48179 8483
rect 47961 8245 47995 8279
rect 45569 7905 45603 7939
rect 47133 7905 47167 7939
rect 47409 7905 47443 7939
rect 45661 7769 45695 7803
rect 46581 7769 46615 7803
rect 47225 7769 47259 7803
rect 47593 7497 47627 7531
rect 46305 7361 46339 7395
rect 47777 7361 47811 7395
rect 46765 7293 46799 7327
rect 46029 7157 46063 7191
rect 46397 7157 46431 7191
rect 38669 6817 38703 6851
rect 47317 6817 47351 6851
rect 47593 6749 47627 6783
rect 37657 6681 37691 6715
rect 37749 6681 37783 6715
rect 37289 6613 37323 6647
rect 37565 6409 37599 6443
rect 48053 6409 48087 6443
rect 38485 6341 38519 6375
rect 39405 6341 39439 6375
rect 37749 6273 37783 6307
rect 47961 6273 47995 6307
rect 38393 6205 38427 6239
rect 37749 5321 37783 5355
rect 37289 5185 37323 5219
rect 39681 5185 39715 5219
rect 47869 5185 47903 5219
rect 48053 5049 48087 5083
rect 37381 4981 37415 5015
rect 39773 4981 39807 5015
rect 41889 4641 41923 4675
rect 42349 4641 42383 4675
rect 43269 4641 43303 4675
rect 47593 4641 47627 4675
rect 14473 4573 14507 4607
rect 15117 4573 15151 4607
rect 15209 4573 15243 4607
rect 15761 4573 15795 4607
rect 15853 4573 15887 4607
rect 16405 4573 16439 4607
rect 16497 4573 16531 4607
rect 17049 4573 17083 4607
rect 20913 4573 20947 4607
rect 21005 4573 21039 4607
rect 21557 4573 21591 4607
rect 39129 4573 39163 4607
rect 39865 4573 39899 4607
rect 40877 4573 40911 4607
rect 46673 4573 46707 4607
rect 47317 4573 47351 4607
rect 26157 4505 26191 4539
rect 26249 4505 26283 4539
rect 27169 4505 27203 4539
rect 40049 4505 40083 4539
rect 42441 4505 42475 4539
rect 14565 4437 14599 4471
rect 17141 4437 17175 4471
rect 21649 4437 21683 4471
rect 39221 4437 39255 4471
rect 40233 4437 40267 4471
rect 40693 4437 40727 4471
rect 46765 4437 46799 4471
rect 14565 4233 14599 4267
rect 21189 4233 21223 4267
rect 46857 4233 46891 4267
rect 42901 4165 42935 4199
rect 43821 4165 43855 4199
rect 46581 4165 46615 4199
rect 47777 4165 47811 4199
rect 2053 4097 2087 4131
rect 10609 4097 10643 4131
rect 13553 4097 13587 4131
rect 14473 4097 14507 4131
rect 15853 4097 15887 4131
rect 16957 4097 16991 4131
rect 17969 4097 18003 4131
rect 19533 4097 19567 4131
rect 20453 4097 20487 4131
rect 21097 4097 21131 4131
rect 22017 4097 22051 4131
rect 38393 4097 38427 4131
rect 39221 4097 39255 4131
rect 39681 4097 39715 4131
rect 44465 4097 44499 4131
rect 7205 4029 7239 4063
rect 7389 4029 7423 4063
rect 8217 4029 8251 4063
rect 38485 4029 38519 4063
rect 39865 4029 39899 4063
rect 41429 4029 41463 4063
rect 42809 4029 42843 4063
rect 22845 3961 22879 3995
rect 2145 3893 2179 3927
rect 2881 3893 2915 3927
rect 10701 3893 10735 3927
rect 13645 3893 13679 3927
rect 15301 3893 15335 3927
rect 15945 3893 15979 3927
rect 17049 3893 17083 3927
rect 18061 3893 18095 3927
rect 19625 3893 19659 3927
rect 20545 3893 20579 3927
rect 22109 3893 22143 3927
rect 39037 3893 39071 3927
rect 44281 3893 44315 3927
rect 46029 3893 46063 3927
rect 47869 3893 47903 3927
rect 8125 3689 8159 3723
rect 17509 3689 17543 3723
rect 21741 3689 21775 3723
rect 39221 3689 39255 3723
rect 40141 3689 40175 3723
rect 40417 3689 40451 3723
rect 33885 3621 33919 3655
rect 3985 3553 4019 3587
rect 10701 3553 10735 3587
rect 10977 3553 11011 3587
rect 15117 3553 15151 3587
rect 15301 3553 15335 3587
rect 16037 3553 16071 3587
rect 23581 3553 23615 3587
rect 26157 3553 26191 3587
rect 27169 3553 27203 3587
rect 41061 3553 41095 3587
rect 41429 3553 41463 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 2697 3485 2731 3519
rect 6745 3485 6779 3519
rect 7389 3485 7423 3519
rect 8033 3485 8067 3519
rect 9321 3485 9355 3519
rect 9873 3485 9907 3519
rect 10517 3485 10551 3519
rect 13369 3485 13403 3519
rect 14289 3485 14323 3519
rect 17417 3485 17451 3519
rect 18061 3485 18095 3519
rect 19257 3485 19291 3519
rect 19901 3485 19935 3519
rect 20545 3485 20579 3519
rect 22017 3485 22051 3519
rect 22845 3485 22879 3519
rect 23489 3485 23523 3519
rect 24777 3485 24811 3519
rect 25605 3485 25639 3519
rect 33057 3485 33091 3519
rect 39129 3485 39163 3519
rect 39865 3485 39899 3519
rect 40233 3485 40267 3519
rect 40877 3485 40911 3519
rect 43177 3485 43211 3519
rect 44005 3485 44039 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 1869 3417 1903 3451
rect 2237 3417 2271 3451
rect 26249 3417 26283 3451
rect 48145 3417 48179 3451
rect 2789 3349 2823 3383
rect 7481 3349 7515 3383
rect 9965 3349 9999 3383
rect 13461 3349 13495 3383
rect 18153 3349 18187 3383
rect 19349 3349 19383 3383
rect 19993 3349 20027 3383
rect 20637 3349 20671 3383
rect 24869 3349 24903 3383
rect 33149 3349 33183 3383
rect 43269 3349 43303 3383
rect 45753 3349 45787 3383
rect 16773 3145 16807 3179
rect 18245 3145 18279 3179
rect 18889 3145 18923 3179
rect 19533 3145 19567 3179
rect 20177 3145 20211 3179
rect 20821 3145 20855 3179
rect 39865 3145 39899 3179
rect 41061 3145 41095 3179
rect 47869 3145 47903 3179
rect 1961 3077 1995 3111
rect 6745 3077 6779 3111
rect 9321 3077 9355 3111
rect 15945 3077 15979 3111
rect 33149 3077 33183 3111
rect 42993 3077 43027 3111
rect 45385 3077 45419 3111
rect 1777 3009 1811 3043
rect 6561 3009 6595 3043
rect 9137 3009 9171 3043
rect 12725 3009 12759 3043
rect 13553 3009 13587 3043
rect 15853 3009 15887 3043
rect 16681 3009 16715 3043
rect 17417 3009 17451 3043
rect 17509 3009 17543 3043
rect 18153 3009 18187 3043
rect 18797 3009 18831 3043
rect 19441 3009 19475 3043
rect 20085 3009 20119 3043
rect 20729 3009 20763 3043
rect 21925 3009 21959 3043
rect 24593 3009 24627 3043
rect 26985 3009 27019 3043
rect 27997 3009 28031 3043
rect 28181 3009 28215 3043
rect 32965 3009 32999 3043
rect 39405 3009 39439 3043
rect 42809 3009 42843 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2237 2941 2271 2975
rect 7021 2941 7055 2975
rect 9597 2941 9631 2975
rect 12633 2941 12667 2975
rect 13737 2941 13771 2975
rect 14197 2941 14231 2975
rect 22109 2941 22143 2975
rect 22569 2941 22603 2975
rect 24777 2941 24811 2975
rect 25145 2941 25179 2975
rect 27445 2941 27479 2975
rect 33517 2941 33551 2975
rect 39221 2941 39255 2975
rect 40417 2941 40451 2975
rect 40601 2941 40635 2975
rect 43269 2941 43303 2975
rect 47041 2941 47075 2975
rect 13093 2805 13127 2839
rect 27261 2805 27295 2839
rect 4537 2601 4571 2635
rect 7481 2601 7515 2635
rect 10793 2601 10827 2635
rect 13461 2601 13495 2635
rect 14197 2601 14231 2635
rect 19901 2601 19935 2635
rect 20913 2601 20947 2635
rect 22385 2601 22419 2635
rect 23397 2601 23431 2635
rect 24961 2601 24995 2635
rect 26249 2601 26283 2635
rect 28641 2601 28675 2635
rect 35541 2601 35575 2635
rect 36369 2601 36403 2635
rect 39129 2601 39163 2635
rect 41705 2601 41739 2635
rect 42533 2601 42567 2635
rect 42901 2601 42935 2635
rect 15853 2533 15887 2567
rect 41245 2533 41279 2567
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2881 2465 2915 2499
rect 9689 2465 9723 2499
rect 27261 2465 27295 2499
rect 38393 2465 38427 2499
rect 40509 2465 40543 2499
rect 46489 2465 46523 2499
rect 47869 2465 47903 2499
rect 5457 2397 5491 2431
rect 13369 2397 13403 2431
rect 14105 2397 14139 2431
rect 16681 2397 16715 2431
rect 19809 2397 19843 2431
rect 23581 2397 23615 2431
rect 26433 2397 26467 2431
rect 26985 2397 27019 2431
rect 28457 2397 28491 2431
rect 29929 2397 29963 2431
rect 35725 2397 35759 2431
rect 39313 2397 39347 2431
rect 41889 2397 41923 2431
rect 42441 2397 42475 2431
rect 43637 2397 43671 2431
rect 43913 2397 43947 2431
rect 46213 2397 46247 2431
rect 47685 2397 47719 2431
rect 4261 2329 4295 2363
rect 9413 2329 9447 2363
rect 15669 2329 15703 2363
rect 20821 2329 20855 2363
rect 22293 2329 22327 2363
rect 24869 2329 24903 2363
rect 36277 2329 36311 2363
rect 38209 2329 38243 2363
rect 40325 2329 40359 2363
rect 41061 2329 41095 2363
rect 45385 2329 45419 2363
rect 5273 2261 5307 2295
rect 16865 2261 16899 2295
rect 29745 2261 29779 2295
rect 45477 2261 45511 2295
<< metal1 >>
rect 44818 47404 44824 47456
rect 44876 47444 44882 47456
rect 45462 47444 45468 47456
rect 44876 47416 45468 47444
rect 44876 47404 44882 47416
rect 45462 47404 45468 47416
rect 45520 47404 45526 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 16899 47175 16957 47181
rect 16899 47141 16911 47175
rect 16945 47172 16957 47175
rect 22278 47172 22284 47184
rect 16945 47144 22284 47172
rect 16945 47141 16957 47144
rect 16899 47135 16957 47141
rect 22278 47132 22284 47144
rect 22336 47132 22342 47184
rect 29917 47175 29975 47181
rect 29917 47141 29929 47175
rect 29963 47172 29975 47175
rect 30190 47172 30196 47184
rect 29963 47144 30196 47172
rect 29963 47141 29975 47144
rect 29917 47135 29975 47141
rect 30190 47132 30196 47144
rect 30248 47132 30254 47184
rect 40126 47172 40132 47184
rect 30576 47144 40132 47172
rect 2041 47107 2099 47113
rect 2041 47073 2053 47107
rect 2087 47104 2099 47107
rect 30576 47104 30604 47144
rect 40126 47132 40132 47144
rect 40184 47132 40190 47184
rect 47949 47175 48007 47181
rect 47949 47141 47961 47175
rect 47995 47172 48007 47175
rect 48038 47172 48044 47184
rect 47995 47144 48044 47172
rect 47995 47141 48007 47144
rect 47949 47135 48007 47141
rect 48038 47132 48044 47144
rect 48096 47132 48102 47184
rect 30742 47104 30748 47116
rect 2087 47076 30604 47104
rect 30703 47076 30748 47104
rect 2087 47073 2099 47076
rect 2041 47067 2099 47073
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 43162 47104 43168 47116
rect 43123 47076 43168 47104
rect 43162 47064 43168 47076
rect 43220 47064 43226 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47036 1823 47039
rect 1946 47036 1952 47048
rect 1811 47008 1952 47036
rect 1811 47005 1823 47008
rect 1765 46999 1823 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4706 47036 4712 47048
rect 4667 47008 4712 47036
rect 3789 46999 3847 47005
rect 4706 46996 4712 47008
rect 4764 46996 4770 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 5868 47008 6377 47036
rect 5868 46996 5874 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 7282 47036 7288 47048
rect 7243 47008 7288 47036
rect 6365 46999 6423 47005
rect 7282 46996 7288 47008
rect 7340 46996 7346 47048
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 9401 46999 9459 47005
rect 11606 46996 11612 47048
rect 11664 47036 11670 47048
rect 11701 47039 11759 47045
rect 11701 47036 11713 47039
rect 11664 47008 11713 47036
rect 11664 46996 11670 47008
rect 11701 47005 11713 47008
rect 11747 47005 11759 47039
rect 11701 46999 11759 47005
rect 12250 46996 12256 47048
rect 12308 47036 12314 47048
rect 12345 47039 12403 47045
rect 12345 47036 12357 47039
rect 12308 47008 12357 47036
rect 12308 46996 12314 47008
rect 12345 47005 12357 47008
rect 12391 47005 12403 47039
rect 12618 47036 12624 47048
rect 12579 47008 12624 47036
rect 12345 46999 12403 47005
rect 12618 46996 12624 47008
rect 12676 46996 12682 47048
rect 13814 46996 13820 47048
rect 13872 47036 13878 47048
rect 15473 47039 15531 47045
rect 15473 47036 15485 47039
rect 13872 47008 15485 47036
rect 13872 46996 13878 47008
rect 15473 47005 15485 47008
rect 15519 47005 15531 47039
rect 15473 46999 15531 47005
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 20714 47036 20720 47048
rect 20675 47008 20720 47036
rect 16669 46999 16727 47005
rect 20714 46996 20720 47008
rect 20772 46996 20778 47048
rect 22005 47039 22063 47045
rect 22005 47036 22017 47039
rect 21008 47008 22017 47036
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 2777 46931 2835 46937
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 2792 46900 2820 46931
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 4982 46968 4988 46980
rect 4943 46940 4988 46968
rect 4982 46928 4988 46940
rect 5040 46928 5046 46980
rect 6638 46968 6644 46980
rect 6599 46940 6644 46968
rect 6638 46928 6644 46940
rect 6696 46928 6702 46980
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 9585 46931 9643 46937
rect 11790 46928 11796 46980
rect 11848 46968 11854 46980
rect 11885 46971 11943 46977
rect 11885 46968 11897 46971
rect 11848 46940 11897 46968
rect 11848 46928 11854 46940
rect 11885 46937 11897 46940
rect 11931 46937 11943 46971
rect 14553 46971 14611 46977
rect 14553 46968 14565 46971
rect 11885 46931 11943 46937
rect 13832 46940 14565 46968
rect 2648 46872 2820 46900
rect 2648 46860 2654 46872
rect 2866 46860 2872 46912
rect 2924 46900 2930 46912
rect 7466 46900 7472 46912
rect 2924 46872 2969 46900
rect 7427 46872 7472 46900
rect 2924 46860 2930 46872
rect 7466 46860 7472 46872
rect 7524 46860 7530 46912
rect 12894 46860 12900 46912
rect 12952 46900 12958 46912
rect 13832 46900 13860 46940
rect 14553 46937 14565 46940
rect 14599 46937 14611 46971
rect 14553 46931 14611 46937
rect 15562 46928 15568 46980
rect 15620 46968 15626 46980
rect 15657 46971 15715 46977
rect 15657 46968 15669 46971
rect 15620 46940 15669 46968
rect 15620 46928 15626 46940
rect 15657 46937 15669 46940
rect 15703 46937 15715 46971
rect 15657 46931 15715 46937
rect 19705 46971 19763 46977
rect 19705 46937 19717 46971
rect 19751 46937 19763 46971
rect 20070 46968 20076 46980
rect 20031 46940 20076 46968
rect 19705 46931 19763 46937
rect 14642 46900 14648 46912
rect 12952 46872 13860 46900
rect 14603 46872 14648 46900
rect 12952 46860 12958 46872
rect 14642 46860 14648 46872
rect 14700 46860 14706 46912
rect 18690 46860 18696 46912
rect 18748 46900 18754 46912
rect 19720 46900 19748 46931
rect 20070 46928 20076 46940
rect 20128 46928 20134 46980
rect 18748 46872 19748 46900
rect 18748 46860 18754 46872
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 21008 46900 21036 47008
rect 22005 47005 22017 47008
rect 22051 47005 22063 47039
rect 22005 46999 22063 47005
rect 28442 46996 28448 47048
rect 28500 47036 28506 47048
rect 28721 47039 28779 47045
rect 28721 47036 28733 47039
rect 28500 47008 28733 47036
rect 28500 46996 28506 47008
rect 28721 47005 28733 47008
rect 28767 47005 28779 47039
rect 28721 46999 28779 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 31021 47039 31079 47045
rect 31021 47005 31033 47039
rect 31067 47036 31079 47039
rect 31570 47036 31576 47048
rect 31067 47008 31576 47036
rect 31067 47005 31079 47008
rect 31021 46999 31079 47005
rect 31570 46996 31576 47008
rect 31628 46996 31634 47048
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 38381 46999 38439 47005
rect 40218 46996 40224 47048
rect 40276 47036 40282 47048
rect 40497 47039 40555 47045
rect 40497 47036 40509 47039
rect 40276 47008 40509 47036
rect 40276 46996 40282 47008
rect 40497 47005 40509 47008
rect 40543 47005 40555 47039
rect 40497 46999 40555 47005
rect 41877 47039 41935 47045
rect 41877 47005 41889 47039
rect 41923 47036 41935 47039
rect 42613 47039 42671 47045
rect 42613 47036 42625 47039
rect 41923 47008 42625 47036
rect 41923 47005 41935 47008
rect 41877 46999 41935 47005
rect 42613 47005 42625 47008
rect 42659 47005 42671 47039
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 42613 46999 42671 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 28350 46928 28356 46980
rect 28408 46968 28414 46980
rect 28537 46971 28595 46977
rect 28537 46968 28549 46971
rect 28408 46940 28549 46968
rect 28408 46928 28414 46940
rect 28537 46937 28549 46940
rect 28583 46937 28595 46971
rect 28537 46931 28595 46937
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 42794 46968 42800 46980
rect 42755 46940 42800 46968
rect 40313 46931 40371 46937
rect 21818 46900 21824 46912
rect 20036 46872 21036 46900
rect 21779 46872 21824 46900
rect 20036 46860 20042 46872
rect 21818 46860 21824 46872
rect 21876 46860 21882 46912
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 42794 46928 42800 46940
rect 42852 46928 42858 46980
rect 45094 46928 45100 46980
rect 45152 46968 45158 46980
rect 45373 46971 45431 46977
rect 45373 46968 45385 46971
rect 45152 46940 45385 46968
rect 45152 46928 45158 46940
rect 45373 46937 45385 46940
rect 45419 46937 45431 46971
rect 45373 46931 45431 46937
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1854 46628 1860 46640
rect 1815 46600 1860 46628
rect 1854 46588 1860 46600
rect 1912 46588 1918 46640
rect 3878 46588 3884 46640
rect 3936 46628 3942 46640
rect 5813 46631 5871 46637
rect 5813 46628 5825 46631
rect 3936 46600 5825 46628
rect 3936 46588 3942 46600
rect 5813 46597 5825 46600
rect 5859 46597 5871 46631
rect 5813 46591 5871 46597
rect 32030 46588 32036 46640
rect 32088 46628 32094 46640
rect 32309 46631 32367 46637
rect 32309 46628 32321 46631
rect 32088 46600 32321 46628
rect 32088 46588 32094 46600
rect 32309 46597 32321 46600
rect 32355 46597 32367 46631
rect 32309 46591 32367 46597
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 47946 46560 47952 46572
rect 47907 46532 47952 46560
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 3970 46492 3976 46504
rect 3931 46464 3976 46492
rect 3970 46452 3976 46464
rect 4028 46452 4034 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46492 4215 46495
rect 5166 46492 5172 46504
rect 4203 46464 5172 46492
rect 4203 46461 4215 46464
rect 4157 46455 4215 46461
rect 5166 46452 5172 46464
rect 5224 46452 5230 46504
rect 13173 46495 13231 46501
rect 13173 46461 13185 46495
rect 13219 46492 13231 46495
rect 13633 46495 13691 46501
rect 13633 46492 13645 46495
rect 13219 46464 13645 46492
rect 13219 46461 13231 46464
rect 13173 46455 13231 46461
rect 13633 46461 13645 46464
rect 13679 46461 13691 46495
rect 13633 46455 13691 46461
rect 13817 46495 13875 46501
rect 13817 46461 13829 46495
rect 13863 46492 13875 46495
rect 14182 46492 14188 46504
rect 13863 46464 14188 46492
rect 13863 46461 13875 46464
rect 13817 46455 13875 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 18969 46495 19027 46501
rect 14332 46464 14377 46492
rect 14332 46452 14338 46464
rect 18969 46461 18981 46495
rect 19015 46492 19027 46495
rect 19429 46495 19487 46501
rect 19429 46492 19441 46495
rect 19015 46464 19441 46492
rect 19015 46461 19027 46464
rect 18969 46455 19027 46461
rect 19429 46461 19441 46464
rect 19475 46461 19487 46495
rect 19610 46492 19616 46504
rect 19571 46464 19616 46492
rect 19429 46455 19487 46461
rect 19610 46452 19616 46464
rect 19668 46452 19674 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 26329 46495 26387 46501
rect 26329 46461 26341 46495
rect 26375 46492 26387 46495
rect 26973 46495 27031 46501
rect 26973 46492 26985 46495
rect 26375 46464 26985 46492
rect 26375 46461 26387 46464
rect 26329 46455 26387 46461
rect 26973 46461 26985 46464
rect 27019 46461 27031 46495
rect 26973 46455 27031 46461
rect 27157 46495 27215 46501
rect 27157 46461 27169 46495
rect 27203 46492 27215 46495
rect 27614 46492 27620 46504
rect 27203 46464 27620 46492
rect 27203 46461 27215 46464
rect 27157 46455 27215 46461
rect 27614 46452 27620 46464
rect 27672 46452 27678 46504
rect 27709 46495 27767 46501
rect 27709 46461 27721 46495
rect 27755 46461 27767 46495
rect 27709 46455 27767 46461
rect 31573 46495 31631 46501
rect 31573 46461 31585 46495
rect 31619 46492 31631 46495
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 31619 46464 32137 46492
rect 31619 46461 31631 46464
rect 31573 46455 31631 46461
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32125 46455 32183 46461
rect 2038 46424 2044 46436
rect 1999 46396 2044 46424
rect 2038 46384 2044 46396
rect 2096 46384 2102 46436
rect 25774 46384 25780 46436
rect 25832 46424 25838 46436
rect 27724 46424 27752 46455
rect 32306 46452 32312 46504
rect 32364 46492 32370 46504
rect 32585 46495 32643 46501
rect 32585 46492 32597 46495
rect 32364 46464 32597 46492
rect 32364 46452 32370 46464
rect 32585 46461 32597 46464
rect 32631 46461 32643 46495
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 32585 46455 32643 46461
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 45186 46492 45192 46504
rect 45147 46464 45192 46492
rect 42889 46455 42947 46461
rect 25832 46396 27752 46424
rect 25832 46384 25838 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 45186 46452 45192 46464
rect 45244 46452 45250 46504
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 45554 46492 45560 46504
rect 45419 46464 45560 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 45554 46452 45560 46464
rect 45612 46452 45618 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 42576 46396 42932 46424
rect 42576 46384 42582 46396
rect 1394 46316 1400 46368
rect 1452 46356 1458 46368
rect 2869 46359 2927 46365
rect 2869 46356 2881 46359
rect 1452 46328 2881 46356
rect 1452 46316 1458 46328
rect 2869 46325 2881 46328
rect 2915 46325 2927 46359
rect 2869 46319 2927 46325
rect 10410 46316 10416 46368
rect 10468 46356 10474 46368
rect 10689 46359 10747 46365
rect 10689 46356 10701 46359
rect 10468 46328 10701 46356
rect 10468 46316 10474 46328
rect 10689 46325 10701 46328
rect 10735 46325 10747 46359
rect 10689 46319 10747 46325
rect 25222 46316 25228 46368
rect 25280 46356 25286 46368
rect 25501 46359 25559 46365
rect 25501 46356 25513 46359
rect 25280 46328 25513 46356
rect 25280 46316 25286 46328
rect 25501 46325 25513 46328
rect 25547 46325 25559 46359
rect 25501 46319 25559 46325
rect 41233 46359 41291 46365
rect 41233 46325 41245 46359
rect 41279 46356 41291 46359
rect 41322 46356 41328 46368
rect 41279 46328 41328 46356
rect 41279 46325 41291 46328
rect 41233 46319 41291 46325
rect 41322 46316 41328 46328
rect 41380 46316 41386 46368
rect 41414 46316 41420 46368
rect 41472 46356 41478 46368
rect 47210 46356 47216 46368
rect 41472 46328 47216 46356
rect 41472 46316 41478 46328
rect 47210 46316 47216 46328
rect 47268 46316 47274 46368
rect 47302 46316 47308 46368
rect 47360 46356 47366 46368
rect 48041 46359 48099 46365
rect 48041 46356 48053 46359
rect 47360 46328 48053 46356
rect 47360 46316 47366 46328
rect 48041 46325 48053 46328
rect 48087 46325 48099 46359
rect 48041 46319 48099 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3970 46112 3976 46164
rect 4028 46152 4034 46164
rect 4433 46155 4491 46161
rect 4433 46152 4445 46155
rect 4028 46124 4445 46152
rect 4028 46112 4034 46124
rect 4433 46121 4445 46124
rect 4479 46121 4491 46155
rect 5166 46152 5172 46164
rect 5127 46124 5172 46152
rect 4433 46115 4491 46121
rect 5166 46112 5172 46124
rect 5224 46112 5230 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 18601 46155 18659 46161
rect 18601 46121 18613 46155
rect 18647 46152 18659 46155
rect 19610 46152 19616 46164
rect 18647 46124 19616 46152
rect 18647 46121 18659 46124
rect 18601 46115 18659 46121
rect 19610 46112 19616 46124
rect 19668 46112 19674 46164
rect 27614 46152 27620 46164
rect 20088 46124 27476 46152
rect 27575 46124 27620 46152
rect 6886 46056 16574 46084
rect 1394 46016 1400 46028
rect 1355 45988 1400 46016
rect 1394 45976 1400 45988
rect 1452 45976 1458 46028
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 5077 45951 5135 45957
rect 5077 45917 5089 45951
rect 5123 45948 5135 45951
rect 6886 45948 6914 46056
rect 10410 46016 10416 46028
rect 10371 45988 10416 46016
rect 10410 45976 10416 45988
rect 10468 45976 10474 46028
rect 10962 45976 10968 46028
rect 11020 46016 11026 46028
rect 11057 46019 11115 46025
rect 11057 46016 11069 46019
rect 11020 45988 11069 46016
rect 11020 45976 11026 45988
rect 11057 45985 11069 45988
rect 11103 45985 11115 46019
rect 16546 46016 16574 46056
rect 20088 46016 20116 46124
rect 20714 46084 20720 46096
rect 16546 45988 20116 46016
rect 20180 46056 20720 46084
rect 11057 45979 11115 45985
rect 14090 45948 14096 45960
rect 5123 45920 6914 45948
rect 14003 45920 14096 45948
rect 5123 45917 5135 45920
rect 5077 45911 5135 45917
rect 14090 45908 14096 45920
rect 14148 45948 14154 45960
rect 18414 45948 18420 45960
rect 14148 45920 18420 45948
rect 14148 45908 14154 45920
rect 18414 45908 18420 45920
rect 18472 45948 18478 45960
rect 18509 45951 18567 45957
rect 18509 45948 18521 45951
rect 18472 45920 18521 45948
rect 18472 45908 18478 45920
rect 18509 45917 18521 45920
rect 18555 45917 18567 45951
rect 18509 45911 18567 45917
rect 18598 45908 18604 45960
rect 18656 45948 18662 45960
rect 20180 45957 20208 46056
rect 20714 46044 20720 46056
rect 20772 46044 20778 46096
rect 26234 45976 26240 46028
rect 26292 46016 26298 46028
rect 26292 45988 26337 46016
rect 26292 45976 26298 45988
rect 19521 45951 19579 45957
rect 19521 45948 19533 45951
rect 18656 45920 19533 45948
rect 18656 45908 18662 45920
rect 19521 45917 19533 45920
rect 19567 45917 19579 45951
rect 19521 45911 19579 45917
rect 20165 45951 20223 45957
rect 20165 45917 20177 45951
rect 20211 45917 20223 45951
rect 20165 45911 20223 45917
rect 21634 45908 21640 45960
rect 21692 45948 21698 45960
rect 22005 45951 22063 45957
rect 22005 45948 22017 45951
rect 21692 45920 22017 45948
rect 21692 45908 21698 45920
rect 22005 45917 22017 45920
rect 22051 45917 22063 45951
rect 25222 45948 25228 45960
rect 25183 45920 25228 45948
rect 22005 45911 22063 45917
rect 25222 45908 25228 45920
rect 25280 45908 25286 45960
rect 1581 45883 1639 45889
rect 1581 45849 1593 45883
rect 1627 45880 1639 45883
rect 2222 45880 2228 45892
rect 1627 45852 2228 45880
rect 1627 45849 1639 45852
rect 1581 45843 1639 45849
rect 2222 45840 2228 45852
rect 2280 45840 2286 45892
rect 10594 45880 10600 45892
rect 10555 45852 10600 45880
rect 10594 45840 10600 45852
rect 10652 45840 10658 45892
rect 19613 45883 19671 45889
rect 19613 45849 19625 45883
rect 19659 45880 19671 45883
rect 20349 45883 20407 45889
rect 20349 45880 20361 45883
rect 19659 45852 20361 45880
rect 19659 45849 19671 45852
rect 19613 45843 19671 45849
rect 20349 45849 20361 45852
rect 20395 45849 20407 45883
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 20349 45843 20407 45849
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 25498 45840 25504 45892
rect 25556 45880 25562 45892
rect 27448 45880 27476 46124
rect 27614 46112 27620 46124
rect 27672 46112 27678 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 42426 46152 42432 46164
rect 39132 46124 42432 46152
rect 39132 46084 39160 46124
rect 42426 46112 42432 46124
rect 42484 46112 42490 46164
rect 41414 46084 41420 46096
rect 27540 46056 39160 46084
rect 40696 46056 41420 46084
rect 27540 45957 27568 46056
rect 40696 46016 40724 46056
rect 41414 46044 41420 46056
rect 41472 46044 41478 46096
rect 41322 46016 41328 46028
rect 35866 45988 40724 46016
rect 41283 45988 41328 46016
rect 27525 45951 27583 45957
rect 27525 45917 27537 45951
rect 27571 45917 27583 45951
rect 27525 45911 27583 45917
rect 35866 45880 35894 45988
rect 41322 45976 41328 45988
rect 41380 45976 41386 46028
rect 41874 46016 41880 46028
rect 41835 45988 41880 46016
rect 41874 45976 41880 45988
rect 41932 45976 41938 46028
rect 46293 46019 46351 46025
rect 46293 45985 46305 46019
rect 46339 46016 46351 46019
rect 46474 46016 46480 46028
rect 46339 45988 46480 46016
rect 46339 45985 46351 45988
rect 46293 45979 46351 45985
rect 46474 45976 46480 45988
rect 46532 45976 46538 46028
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 38194 45948 38200 45960
rect 38155 45920 38200 45948
rect 38194 45908 38200 45920
rect 38252 45908 38258 45960
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43993 45951 44051 45957
rect 43993 45948 44005 45951
rect 43864 45920 44005 45948
rect 43864 45908 43870 45920
rect 43993 45917 44005 45920
rect 44039 45917 44051 45951
rect 43993 45911 44051 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 41506 45880 41512 45892
rect 25556 45852 26740 45880
rect 27448 45852 35894 45880
rect 41467 45852 41512 45880
rect 25556 45840 25562 45852
rect 25130 45772 25136 45824
rect 25188 45812 25194 45824
rect 26234 45812 26240 45824
rect 25188 45784 26240 45812
rect 25188 45772 25194 45784
rect 26234 45772 26240 45784
rect 26292 45772 26298 45824
rect 26712 45812 26740 45852
rect 41506 45840 41512 45852
rect 41564 45840 41570 45892
rect 44174 45880 44180 45892
rect 44135 45852 44180 45880
rect 44174 45840 44180 45852
rect 44232 45840 44238 45892
rect 46477 45883 46535 45889
rect 46477 45849 46489 45883
rect 46523 45880 46535 45883
rect 47670 45880 47676 45892
rect 46523 45852 47676 45880
rect 46523 45849 46535 45852
rect 46477 45843 46535 45849
rect 47670 45840 47676 45852
rect 47728 45840 47734 45892
rect 45741 45815 45799 45821
rect 45741 45812 45753 45815
rect 26712 45784 45753 45812
rect 45741 45781 45753 45784
rect 45787 45781 45799 45815
rect 45741 45775 45799 45781
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 2222 45608 2228 45620
rect 2183 45580 2228 45608
rect 2222 45568 2228 45580
rect 2280 45568 2286 45620
rect 10594 45608 10600 45620
rect 10555 45580 10600 45608
rect 10594 45568 10600 45580
rect 10652 45568 10658 45620
rect 25406 45568 25412 45620
rect 25464 45608 25470 45620
rect 26145 45611 26203 45617
rect 26145 45608 26157 45611
rect 25464 45580 26157 45608
rect 25464 45568 25470 45580
rect 26145 45577 26157 45580
rect 26191 45577 26203 45611
rect 26145 45571 26203 45577
rect 38194 45568 38200 45620
rect 38252 45608 38258 45620
rect 41417 45611 41475 45617
rect 38252 45580 38654 45608
rect 38252 45568 38258 45580
rect 38626 45540 38654 45580
rect 40144 45580 41368 45608
rect 40144 45540 40172 45580
rect 38626 45512 40172 45540
rect 41340 45540 41368 45580
rect 41417 45577 41429 45611
rect 41463 45608 41475 45611
rect 41506 45608 41512 45620
rect 41463 45580 41512 45608
rect 41463 45577 41475 45580
rect 41417 45571 41475 45577
rect 41506 45568 41512 45580
rect 41564 45568 41570 45620
rect 42521 45611 42579 45617
rect 41616 45580 42472 45608
rect 41616 45540 41644 45580
rect 41340 45512 41644 45540
rect 42444 45540 42472 45580
rect 42521 45577 42533 45611
rect 42567 45608 42579 45611
rect 42610 45608 42616 45620
rect 42567 45580 42616 45608
rect 42567 45577 42579 45580
rect 42521 45571 42579 45577
rect 42610 45568 42616 45580
rect 42668 45568 42674 45620
rect 45738 45608 45744 45620
rect 42720 45580 45744 45608
rect 42720 45540 42748 45580
rect 45738 45568 45744 45580
rect 45796 45568 45802 45620
rect 42444 45512 42748 45540
rect 43625 45543 43683 45549
rect 43625 45509 43637 45543
rect 43671 45540 43683 45543
rect 44361 45543 44419 45549
rect 44361 45540 44373 45543
rect 43671 45512 44373 45540
rect 43671 45509 43683 45512
rect 43625 45503 43683 45509
rect 44361 45509 44373 45512
rect 44407 45509 44419 45543
rect 46566 45540 46572 45552
rect 46527 45512 46572 45540
rect 44361 45503 44419 45509
rect 46566 45500 46572 45512
rect 46624 45500 46630 45552
rect 47670 45540 47676 45552
rect 47631 45512 47676 45540
rect 47670 45500 47676 45512
rect 47728 45500 47734 45552
rect 2133 45475 2191 45481
rect 2133 45441 2145 45475
rect 2179 45472 2191 45475
rect 2314 45472 2320 45484
rect 2179 45444 2320 45472
rect 2179 45441 2191 45444
rect 2133 45435 2191 45441
rect 2314 45432 2320 45444
rect 2372 45472 2378 45484
rect 10505 45475 10563 45481
rect 10505 45472 10517 45475
rect 2372 45444 10517 45472
rect 2372 45432 2378 45444
rect 10505 45441 10517 45444
rect 10551 45472 10563 45475
rect 18506 45472 18512 45484
rect 10551 45444 18512 45472
rect 10551 45441 10563 45444
rect 10505 45435 10563 45441
rect 18506 45432 18512 45444
rect 18564 45432 18570 45484
rect 26050 45472 26056 45484
rect 26011 45444 26056 45472
rect 26050 45432 26056 45444
rect 26108 45432 26114 45484
rect 41322 45472 41328 45484
rect 41283 45444 41328 45472
rect 41322 45432 41328 45444
rect 41380 45432 41386 45484
rect 42426 45472 42432 45484
rect 42387 45444 42432 45472
rect 42426 45432 42432 45444
rect 42484 45432 42490 45484
rect 42886 45432 42892 45484
rect 42944 45472 42950 45484
rect 43533 45475 43591 45481
rect 43533 45472 43545 45475
rect 42944 45444 43545 45472
rect 42944 45432 42950 45444
rect 43533 45441 43545 45444
rect 43579 45441 43591 45475
rect 43533 45435 43591 45441
rect 47210 45432 47216 45484
rect 47268 45472 47274 45484
rect 47486 45472 47492 45484
rect 47268 45444 47492 45472
rect 47268 45432 47274 45444
rect 47486 45432 47492 45444
rect 47544 45472 47550 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 47544 45444 47593 45472
rect 47544 45432 47550 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 44177 45407 44235 45413
rect 44177 45373 44189 45407
rect 44223 45404 44235 45407
rect 44450 45404 44456 45416
rect 44223 45376 44456 45404
rect 44223 45373 44235 45376
rect 44177 45367 44235 45373
rect 44450 45364 44456 45376
rect 44508 45364 44514 45416
rect 45370 45404 45376 45416
rect 45331 45376 45376 45404
rect 45370 45364 45376 45376
rect 45428 45364 45434 45416
rect 43254 45228 43260 45280
rect 43312 45268 43318 45280
rect 46661 45271 46719 45277
rect 46661 45268 46673 45271
rect 43312 45240 46673 45268
rect 43312 45228 43318 45240
rect 46661 45237 46673 45240
rect 46707 45237 46719 45271
rect 46661 45231 46719 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 42794 45024 42800 45076
rect 42852 45064 42858 45076
rect 43073 45067 43131 45073
rect 43073 45064 43085 45067
rect 42852 45036 43085 45064
rect 42852 45024 42858 45036
rect 43073 45033 43085 45036
rect 43119 45033 43131 45067
rect 43073 45027 43131 45033
rect 44453 44931 44511 44937
rect 44453 44897 44465 44931
rect 44499 44928 44511 44931
rect 45922 44928 45928 44940
rect 44499 44900 45928 44928
rect 44499 44897 44511 44900
rect 44453 44891 44511 44897
rect 45922 44888 45928 44900
rect 45980 44888 45986 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 38654 44860 38660 44872
rect 38567 44832 38660 44860
rect 38654 44820 38660 44832
rect 38712 44860 38718 44872
rect 42886 44860 42892 44872
rect 38712 44832 42892 44860
rect 38712 44820 38718 44832
rect 42886 44820 42892 44832
rect 42944 44820 42950 44872
rect 42981 44863 43039 44869
rect 42981 44829 42993 44863
rect 43027 44829 43039 44863
rect 45462 44860 45468 44872
rect 45423 44832 45468 44860
rect 42981 44823 43039 44829
rect 38746 44724 38752 44736
rect 38707 44696 38752 44724
rect 38746 44684 38752 44696
rect 38804 44684 38810 44736
rect 42996 44724 43024 44823
rect 45462 44820 45468 44832
rect 45520 44820 45526 44872
rect 46290 44860 46296 44872
rect 46251 44832 46296 44860
rect 46290 44820 46296 44832
rect 46348 44820 46354 44872
rect 45646 44792 45652 44804
rect 45607 44764 45652 44792
rect 45646 44752 45652 44764
rect 45704 44752 45710 44804
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 47670 44792 47676 44804
rect 46523 44764 47676 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 47670 44752 47676 44764
rect 47728 44752 47734 44804
rect 47578 44724 47584 44736
rect 42996 44696 47584 44724
rect 47578 44684 47584 44696
rect 47636 44684 47642 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 45554 44480 45560 44532
rect 45612 44520 45618 44532
rect 45649 44523 45707 44529
rect 45649 44520 45661 44523
rect 45612 44492 45661 44520
rect 45612 44480 45618 44492
rect 45649 44489 45661 44492
rect 45695 44489 45707 44523
rect 47670 44520 47676 44532
rect 47631 44492 47676 44520
rect 45649 44483 45707 44489
rect 47670 44480 47676 44492
rect 47728 44480 47734 44532
rect 38746 44452 38752 44464
rect 38707 44424 38752 44452
rect 38746 44412 38752 44424
rect 38804 44412 38810 44464
rect 46290 44452 46296 44464
rect 45112 44424 46296 44452
rect 44450 44384 44456 44396
rect 44411 44356 44456 44384
rect 44450 44344 44456 44356
rect 44508 44344 44514 44396
rect 45112 44393 45140 44424
rect 46290 44412 46296 44424
rect 46348 44412 46354 44464
rect 45097 44387 45155 44393
rect 45097 44353 45109 44387
rect 45143 44353 45155 44387
rect 45097 44347 45155 44353
rect 45557 44387 45615 44393
rect 45557 44353 45569 44387
rect 45603 44384 45615 44387
rect 45738 44384 45744 44396
rect 45603 44356 45744 44384
rect 45603 44353 45615 44356
rect 45557 44347 45615 44353
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46198 44384 46204 44396
rect 46159 44356 46204 44384
rect 46198 44344 46204 44356
rect 46256 44344 46262 44396
rect 46845 44387 46903 44393
rect 46845 44353 46857 44387
rect 46891 44384 46903 44387
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 46891 44356 47593 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 38562 44316 38568 44328
rect 38523 44288 38568 44316
rect 38562 44276 38568 44288
rect 38620 44276 38626 44328
rect 40034 44316 40040 44328
rect 39995 44288 40040 44316
rect 40034 44276 40040 44288
rect 40092 44276 40098 44328
rect 41322 44276 41328 44328
rect 41380 44316 41386 44328
rect 46860 44316 46888 44347
rect 41380 44288 46888 44316
rect 41380 44276 41386 44288
rect 45094 44208 45100 44260
rect 45152 44248 45158 44260
rect 46293 44251 46351 44257
rect 46293 44248 46305 44251
rect 45152 44220 46305 44248
rect 45152 44208 45158 44220
rect 46293 44217 46305 44220
rect 46339 44217 46351 44251
rect 46293 44211 46351 44217
rect 46934 44180 46940 44192
rect 46895 44152 46940 44180
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 45186 43936 45192 43988
rect 45244 43976 45250 43988
rect 45833 43979 45891 43985
rect 45833 43976 45845 43979
rect 45244 43948 45845 43976
rect 45244 43936 45250 43948
rect 45833 43945 45845 43948
rect 45879 43945 45891 43979
rect 45833 43939 45891 43945
rect 45922 43800 45928 43852
rect 45980 43840 45986 43852
rect 46293 43843 46351 43849
rect 46293 43840 46305 43843
rect 45980 43812 46305 43840
rect 45980 43800 45986 43812
rect 46293 43809 46305 43812
rect 46339 43809 46351 43843
rect 46293 43803 46351 43809
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 46934 43840 46940 43852
rect 46523 43812 46940 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 46934 43800 46940 43812
rect 46992 43800 46998 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 26418 43732 26424 43784
rect 26476 43772 26482 43784
rect 26789 43775 26847 43781
rect 26789 43772 26801 43775
rect 26476 43744 26801 43772
rect 26476 43732 26482 43744
rect 26789 43741 26801 43744
rect 26835 43741 26847 43775
rect 26789 43735 26847 43741
rect 26881 43639 26939 43645
rect 26881 43605 26893 43639
rect 26927 43636 26939 43639
rect 38562 43636 38568 43648
rect 26927 43608 38568 43636
rect 26927 43605 26939 43608
rect 26881 43599 26939 43605
rect 38562 43596 38568 43608
rect 38620 43596 38626 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 45278 43256 45284 43308
rect 45336 43296 45342 43308
rect 45925 43299 45983 43305
rect 45925 43296 45937 43299
rect 45336 43268 45937 43296
rect 45336 43256 45342 43268
rect 45925 43265 45937 43268
rect 45971 43265 45983 43299
rect 45925 43259 45983 43265
rect 46474 43256 46480 43308
rect 46532 43296 46538 43308
rect 46569 43299 46627 43305
rect 46569 43296 46581 43299
rect 46532 43268 46581 43296
rect 46532 43256 46538 43268
rect 46569 43265 46581 43268
rect 46615 43265 46627 43299
rect 46569 43259 46627 43265
rect 1486 43188 1492 43240
rect 1544 43228 1550 43240
rect 1581 43231 1639 43237
rect 1581 43228 1593 43231
rect 1544 43200 1593 43228
rect 1544 43188 1550 43200
rect 1581 43197 1593 43200
rect 1627 43197 1639 43231
rect 1581 43191 1639 43197
rect 47762 43092 47768 43104
rect 47723 43064 47768 43092
rect 47762 43052 47768 43064
rect 47820 43052 47826 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46293 42755 46351 42761
rect 46293 42721 46305 42755
rect 46339 42752 46351 42755
rect 47762 42752 47768 42764
rect 46339 42724 47768 42752
rect 46339 42721 46351 42724
rect 46293 42715 46351 42721
rect 47762 42712 47768 42724
rect 47820 42712 47826 42764
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 47578 42208 47584 42220
rect 47539 42180 47584 42208
rect 47578 42168 47584 42180
rect 47636 42168 47642 42220
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46474 41528 46480 41540
rect 46435 41500 46480 41528
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 2133 41219 2191 41225
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46845 41259 46903 41265
rect 46845 41256 46857 41259
rect 46532 41228 46857 41256
rect 46532 41216 46538 41228
rect 46845 41225 46857 41228
rect 46891 41225 46903 41259
rect 46845 41219 46903 41225
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 42426 41080 42432 41132
rect 42484 41120 42490 41132
rect 46753 41123 46811 41129
rect 46753 41120 46765 41123
rect 42484 41092 46765 41120
rect 42484 41080 42490 41092
rect 46753 41089 46765 41092
rect 46799 41089 46811 41123
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 46753 41083 46811 41089
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 48133 40987 48191 40993
rect 48133 40984 48145 40987
rect 45526 40956 48145 40984
rect 39666 40876 39672 40928
rect 39724 40916 39730 40928
rect 45526 40916 45554 40956
rect 48133 40953 48145 40956
rect 48179 40953 48191 40987
rect 48133 40947 48191 40953
rect 39724 40888 45554 40916
rect 39724 40876 39730 40888
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 1946 40372 1952 40384
rect 1907 40344 1952 40372
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 20162 39516 20168 39568
rect 20220 39556 20226 39568
rect 38654 39556 38660 39568
rect 20220 39528 38660 39556
rect 20220 39516 20226 39528
rect 38654 39516 38660 39528
rect 38712 39516 38718 39568
rect 22646 39448 22652 39500
rect 22704 39488 22710 39500
rect 25409 39491 25467 39497
rect 25409 39488 25421 39491
rect 22704 39460 25421 39488
rect 22704 39448 22710 39460
rect 25409 39457 25421 39460
rect 25455 39457 25467 39491
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 25409 39451 25467 39457
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 22462 39420 22468 39432
rect 22423 39392 22468 39420
rect 22462 39380 22468 39392
rect 22520 39380 22526 39432
rect 25225 39423 25283 39429
rect 25225 39389 25237 39423
rect 25271 39420 25283 39423
rect 25498 39420 25504 39432
rect 25271 39392 25504 39420
rect 25271 39389 25283 39392
rect 25225 39383 25283 39389
rect 25498 39380 25504 39392
rect 25556 39380 25562 39432
rect 22557 39355 22615 39361
rect 22557 39321 22569 39355
rect 22603 39352 22615 39355
rect 46477 39355 46535 39361
rect 46477 39352 46489 39355
rect 22603 39324 46489 39352
rect 22603 39321 22615 39324
rect 22557 39315 22615 39321
rect 46477 39321 46489 39324
rect 46523 39321 46535 39355
rect 46477 39315 46535 39321
rect 23474 39244 23480 39296
rect 23532 39284 23538 39296
rect 24857 39287 24915 39293
rect 24857 39284 24869 39287
rect 23532 39256 24869 39284
rect 23532 39244 23538 39256
rect 24857 39253 24869 39256
rect 24903 39253 24915 39287
rect 24857 39247 24915 39253
rect 25314 39244 25320 39296
rect 25372 39284 25378 39296
rect 25372 39256 25417 39284
rect 25372 39244 25378 39256
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 25041 39083 25099 39089
rect 25041 39049 25053 39083
rect 25087 39080 25099 39083
rect 25314 39080 25320 39092
rect 25087 39052 25320 39080
rect 25087 39049 25099 39052
rect 25041 39043 25099 39049
rect 25314 39040 25320 39052
rect 25372 39040 25378 39092
rect 20073 39015 20131 39021
rect 20073 38981 20085 39015
rect 20119 39012 20131 39015
rect 20162 39012 20168 39024
rect 20119 38984 20168 39012
rect 20119 38981 20131 38984
rect 20073 38975 20131 38981
rect 20162 38972 20168 38984
rect 20220 39012 20226 39024
rect 20438 39012 20444 39024
rect 20220 38984 20444 39012
rect 20220 38972 20226 38984
rect 20438 38972 20444 38984
rect 20496 38972 20502 39024
rect 20717 39015 20775 39021
rect 20717 38981 20729 39015
rect 20763 39012 20775 39015
rect 21818 39012 21824 39024
rect 20763 38984 21824 39012
rect 20763 38981 20775 38984
rect 20717 38975 20775 38981
rect 21818 38972 21824 38984
rect 21876 38972 21882 39024
rect 22646 39012 22652 39024
rect 22066 38984 22652 39012
rect 19426 38944 19432 38956
rect 19387 38916 19432 38944
rect 19426 38904 19432 38916
rect 19484 38904 19490 38956
rect 20901 38947 20959 38953
rect 20901 38913 20913 38947
rect 20947 38944 20959 38947
rect 22066 38944 22094 38984
rect 22646 38972 22652 38984
rect 22704 38972 22710 39024
rect 22830 38972 22836 39024
rect 22888 38972 22894 39024
rect 24673 38947 24731 38953
rect 24673 38944 24685 38947
rect 20947 38916 22094 38944
rect 23860 38916 24685 38944
rect 20947 38913 20959 38916
rect 20901 38907 20959 38913
rect 22094 38836 22100 38888
rect 22152 38876 22158 38888
rect 22370 38876 22376 38888
rect 22152 38848 22197 38876
rect 22331 38848 22376 38876
rect 22152 38836 22158 38848
rect 22370 38836 22376 38848
rect 22428 38836 22434 38888
rect 23860 38885 23888 38916
rect 24673 38913 24685 38916
rect 24719 38944 24731 38947
rect 25498 38944 25504 38956
rect 24719 38916 25504 38944
rect 24719 38913 24731 38916
rect 24673 38907 24731 38913
rect 25498 38904 25504 38916
rect 25556 38904 25562 38956
rect 47670 38944 47676 38956
rect 47631 38916 47676 38944
rect 47670 38904 47676 38916
rect 47728 38904 47734 38956
rect 23845 38879 23903 38885
rect 23845 38845 23857 38879
rect 23891 38845 23903 38879
rect 23845 38839 23903 38845
rect 24394 38836 24400 38888
rect 24452 38876 24458 38888
rect 24581 38879 24639 38885
rect 24581 38876 24593 38879
rect 24452 38848 24593 38876
rect 24452 38836 24458 38848
rect 24581 38845 24593 38848
rect 24627 38845 24639 38879
rect 47854 38876 47860 38888
rect 47815 38848 47860 38876
rect 24581 38839 24639 38845
rect 47854 38836 47860 38848
rect 47912 38836 47918 38888
rect 20530 38700 20536 38752
rect 20588 38740 20594 38752
rect 21085 38743 21143 38749
rect 21085 38740 21097 38743
rect 20588 38712 21097 38740
rect 20588 38700 20594 38712
rect 21085 38709 21097 38712
rect 21131 38709 21143 38743
rect 21085 38703 21143 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 22370 38496 22376 38548
rect 22428 38536 22434 38548
rect 22925 38539 22983 38545
rect 22925 38536 22937 38539
rect 22428 38508 22937 38536
rect 22428 38496 22434 38508
rect 22925 38505 22937 38508
rect 22971 38505 22983 38539
rect 41322 38536 41328 38548
rect 22925 38499 22983 38505
rect 24504 38508 41328 38536
rect 20162 38428 20168 38480
rect 20220 38468 20226 38480
rect 24504 38468 24532 38508
rect 41322 38496 41328 38508
rect 41380 38496 41386 38548
rect 20220 38440 24532 38468
rect 20220 38428 20226 38440
rect 12618 38360 12624 38412
rect 12676 38400 12682 38412
rect 12676 38372 21496 38400
rect 12676 38360 12682 38372
rect 18233 38335 18291 38341
rect 18233 38301 18245 38335
rect 18279 38332 18291 38335
rect 19426 38332 19432 38344
rect 18279 38304 19432 38332
rect 18279 38301 18291 38304
rect 18233 38295 18291 38301
rect 19426 38292 19432 38304
rect 19484 38332 19490 38344
rect 20809 38335 20867 38341
rect 20809 38332 20821 38335
rect 19484 38304 20821 38332
rect 19484 38292 19490 38304
rect 20809 38301 20821 38304
rect 20855 38301 20867 38335
rect 20809 38295 20867 38301
rect 18506 38264 18512 38276
rect 18467 38236 18512 38264
rect 18506 38224 18512 38236
rect 18564 38224 18570 38276
rect 20073 38267 20131 38273
rect 20073 38233 20085 38267
rect 20119 38264 20131 38267
rect 20162 38264 20168 38276
rect 20119 38236 20168 38264
rect 20119 38233 20131 38236
rect 20073 38227 20131 38233
rect 20162 38224 20168 38236
rect 20220 38224 20226 38276
rect 21358 38264 21364 38276
rect 21319 38236 21364 38264
rect 21358 38224 21364 38236
rect 21416 38224 21422 38276
rect 21468 38264 21496 38372
rect 22094 38360 22100 38412
rect 22152 38400 22158 38412
rect 24397 38403 24455 38409
rect 24397 38400 24409 38403
rect 22152 38372 24409 38400
rect 22152 38360 22158 38372
rect 24397 38369 24409 38372
rect 24443 38400 24455 38403
rect 26970 38400 26976 38412
rect 24443 38372 26976 38400
rect 24443 38369 24455 38372
rect 24397 38363 24455 38369
rect 26970 38360 26976 38372
rect 27028 38360 27034 38412
rect 23109 38335 23167 38341
rect 23109 38301 23121 38335
rect 23155 38332 23167 38335
rect 23474 38332 23480 38344
rect 23155 38304 23480 38332
rect 23155 38301 23167 38304
rect 23109 38295 23167 38301
rect 23474 38292 23480 38304
rect 23532 38292 23538 38344
rect 23569 38335 23627 38341
rect 23569 38301 23581 38335
rect 23615 38301 23627 38335
rect 23569 38295 23627 38301
rect 23753 38335 23811 38341
rect 23753 38301 23765 38335
rect 23799 38301 23811 38335
rect 23753 38295 23811 38301
rect 23584 38264 23612 38295
rect 21468 38236 23612 38264
rect 23768 38264 23796 38295
rect 25958 38292 25964 38344
rect 26016 38332 26022 38344
rect 27893 38335 27951 38341
rect 27893 38332 27905 38335
rect 26016 38304 27905 38332
rect 26016 38292 26022 38304
rect 27893 38301 27905 38304
rect 27939 38332 27951 38335
rect 29178 38332 29184 38344
rect 27939 38304 29184 38332
rect 27939 38301 27951 38304
rect 27893 38295 27951 38301
rect 29178 38292 29184 38304
rect 29236 38292 29242 38344
rect 46934 38292 46940 38344
rect 46992 38332 46998 38344
rect 47673 38335 47731 38341
rect 47673 38332 47685 38335
rect 46992 38304 47685 38332
rect 46992 38292 46998 38304
rect 47673 38301 47685 38304
rect 47719 38301 47731 38335
rect 47673 38295 47731 38301
rect 23768 38236 24532 38264
rect 24504 38208 24532 38236
rect 24578 38224 24584 38276
rect 24636 38264 24642 38276
rect 24673 38267 24731 38273
rect 24673 38264 24685 38267
rect 24636 38236 24685 38264
rect 24636 38224 24642 38236
rect 24673 38233 24685 38236
rect 24719 38233 24731 38267
rect 24673 38227 24731 38233
rect 25406 38224 25412 38276
rect 25464 38224 25470 38276
rect 23658 38196 23664 38208
rect 23619 38168 23664 38196
rect 23658 38156 23664 38168
rect 23716 38156 23722 38208
rect 24486 38156 24492 38208
rect 24544 38156 24550 38208
rect 26142 38196 26148 38208
rect 26103 38168 26148 38196
rect 26142 38156 26148 38168
rect 26200 38156 26206 38208
rect 27982 38196 27988 38208
rect 27943 38168 27988 38196
rect 27982 38156 27988 38168
rect 28040 38156 28046 38208
rect 28258 38156 28264 38208
rect 28316 38196 28322 38208
rect 38194 38196 38200 38208
rect 28316 38168 38200 38196
rect 28316 38156 28322 38168
rect 38194 38156 38200 38168
rect 38252 38156 38258 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 18693 37995 18751 38001
rect 18693 37961 18705 37995
rect 18739 37992 18751 37995
rect 19426 37992 19432 38004
rect 18739 37964 19432 37992
rect 18739 37961 18751 37964
rect 18693 37955 18751 37961
rect 19426 37952 19432 37964
rect 19484 37952 19490 38004
rect 20809 37995 20867 38001
rect 20809 37961 20821 37995
rect 20855 37992 20867 37995
rect 22830 37992 22836 38004
rect 20855 37964 22836 37992
rect 20855 37961 20867 37964
rect 20809 37955 20867 37961
rect 22830 37952 22836 37964
rect 22888 37952 22894 38004
rect 24578 37992 24584 38004
rect 24539 37964 24584 37992
rect 24578 37952 24584 37964
rect 24636 37952 24642 38004
rect 25406 37952 25412 38004
rect 25464 37992 25470 38004
rect 25501 37995 25559 38001
rect 25501 37992 25513 37995
rect 25464 37964 25513 37992
rect 25464 37952 25470 37964
rect 25501 37961 25513 37964
rect 25547 37961 25559 37995
rect 25501 37955 25559 37961
rect 23658 37884 23664 37936
rect 23716 37924 23722 37936
rect 23716 37896 24716 37924
rect 23716 37884 23722 37896
rect 18509 37859 18567 37865
rect 18509 37825 18521 37859
rect 18555 37856 18567 37859
rect 19058 37856 19064 37868
rect 18555 37828 19064 37856
rect 18555 37825 18567 37828
rect 18509 37819 18567 37825
rect 19058 37816 19064 37828
rect 19116 37816 19122 37868
rect 19426 37856 19432 37868
rect 19387 37828 19432 37856
rect 19426 37816 19432 37828
rect 19484 37816 19490 37868
rect 19610 37816 19616 37868
rect 19668 37856 19674 37868
rect 20717 37859 20775 37865
rect 20717 37856 20729 37859
rect 19668 37828 20729 37856
rect 19668 37816 19674 37828
rect 20717 37825 20729 37828
rect 20763 37825 20775 37859
rect 20717 37819 20775 37825
rect 24305 37859 24363 37865
rect 24305 37825 24317 37859
rect 24351 37825 24363 37859
rect 24305 37819 24363 37825
rect 19705 37791 19763 37797
rect 19705 37788 19717 37791
rect 19444 37760 19717 37788
rect 19444 37732 19472 37760
rect 19705 37757 19717 37760
rect 19751 37757 19763 37791
rect 19705 37751 19763 37757
rect 19426 37680 19432 37732
rect 19484 37680 19490 37732
rect 24320 37720 24348 37819
rect 24394 37816 24400 37868
rect 24452 37856 24458 37868
rect 24688 37865 24716 37896
rect 27982 37884 27988 37936
rect 28040 37884 28046 37936
rect 24673 37859 24731 37865
rect 24452 37828 24497 37856
rect 24452 37816 24458 37828
rect 24673 37825 24685 37859
rect 24719 37825 24731 37859
rect 24673 37819 24731 37825
rect 24854 37816 24860 37868
rect 24912 37856 24918 37868
rect 25409 37859 25467 37865
rect 25409 37856 25421 37859
rect 24912 37828 25421 37856
rect 24912 37816 24918 37828
rect 25409 37825 25421 37828
rect 25455 37856 25467 37859
rect 25958 37856 25964 37868
rect 25455 37828 25964 37856
rect 25455 37825 25467 37828
rect 25409 37819 25467 37825
rect 25958 37816 25964 37828
rect 26016 37816 26022 37868
rect 26970 37856 26976 37868
rect 26931 37828 26976 37856
rect 26970 37816 26976 37828
rect 27028 37816 27034 37868
rect 29178 37856 29184 37868
rect 29091 37828 29184 37856
rect 29178 37816 29184 37828
rect 29236 37856 29242 37868
rect 31018 37856 31024 37868
rect 29236 37828 31024 37856
rect 29236 37816 29242 37828
rect 31018 37816 31024 37828
rect 31076 37816 31082 37868
rect 47486 37816 47492 37868
rect 47544 37856 47550 37868
rect 47581 37859 47639 37865
rect 47581 37856 47593 37859
rect 47544 37828 47593 37856
rect 47544 37816 47550 37828
rect 47581 37825 47593 37828
rect 47627 37825 47639 37859
rect 47581 37819 47639 37825
rect 24486 37788 24492 37800
rect 24447 37760 24492 37788
rect 24486 37748 24492 37760
rect 24544 37748 24550 37800
rect 27246 37788 27252 37800
rect 27207 37760 27252 37788
rect 27246 37748 27252 37760
rect 27304 37748 27310 37800
rect 24946 37720 24952 37732
rect 24320 37692 24952 37720
rect 24946 37680 24952 37692
rect 25004 37680 25010 37732
rect 21358 37612 21364 37664
rect 21416 37652 21422 37664
rect 28258 37652 28264 37664
rect 21416 37624 28264 37652
rect 21416 37612 21422 37624
rect 28258 37612 28264 37624
rect 28316 37612 28322 37664
rect 28718 37652 28724 37664
rect 28679 37624 28724 37652
rect 28718 37612 28724 37624
rect 28776 37612 28782 37664
rect 29270 37652 29276 37664
rect 29231 37624 29276 37652
rect 29270 37612 29276 37624
rect 29328 37612 29334 37664
rect 47670 37652 47676 37664
rect 47631 37624 47676 37652
rect 47670 37612 47676 37624
rect 47728 37612 47734 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 19610 37448 19616 37460
rect 19571 37420 19616 37448
rect 19610 37408 19616 37420
rect 19668 37448 19674 37460
rect 19978 37448 19984 37460
rect 19668 37420 19984 37448
rect 19668 37408 19674 37420
rect 19978 37408 19984 37420
rect 20036 37408 20042 37460
rect 25501 37451 25559 37457
rect 25501 37417 25513 37451
rect 25547 37448 25559 37451
rect 26142 37448 26148 37460
rect 25547 37420 26148 37448
rect 25547 37417 25559 37420
rect 25501 37411 25559 37417
rect 26142 37408 26148 37420
rect 26200 37408 26206 37460
rect 24394 37340 24400 37392
rect 24452 37380 24458 37392
rect 25774 37380 25780 37392
rect 24452 37352 25780 37380
rect 24452 37340 24458 37352
rect 25774 37340 25780 37352
rect 25832 37340 25838 37392
rect 25409 37315 25467 37321
rect 25409 37281 25421 37315
rect 25455 37312 25467 37315
rect 25455 37284 25636 37312
rect 25455 37281 25467 37284
rect 25409 37275 25467 37281
rect 25608 37256 25636 37284
rect 26970 37272 26976 37324
rect 27028 37312 27034 37324
rect 27249 37315 27307 37321
rect 27249 37312 27261 37315
rect 27028 37284 27261 37312
rect 27028 37272 27034 37284
rect 27249 37281 27261 37284
rect 27295 37281 27307 37315
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 27249 37275 27307 37281
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 2041 37207 2099 37213
rect 14182 37204 14188 37256
rect 14240 37244 14246 37256
rect 14642 37244 14648 37256
rect 14240 37216 14648 37244
rect 14240 37204 14246 37216
rect 14642 37204 14648 37216
rect 14700 37244 14706 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 14700 37216 19441 37244
rect 14700 37204 14706 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 19444 37176 19472 37207
rect 20254 37204 20260 37256
rect 20312 37244 20318 37256
rect 21821 37247 21879 37253
rect 21821 37244 21833 37247
rect 20312 37216 21833 37244
rect 20312 37204 20318 37216
rect 21821 37213 21833 37216
rect 21867 37213 21879 37247
rect 24489 37247 24547 37253
rect 24489 37244 24501 37247
rect 21821 37207 21879 37213
rect 22066 37216 24501 37244
rect 22066 37176 22094 37216
rect 24489 37213 24501 37216
rect 24535 37213 24547 37247
rect 25498 37244 25504 37256
rect 25459 37216 25504 37244
rect 24489 37207 24547 37213
rect 25498 37204 25504 37216
rect 25556 37204 25562 37256
rect 25590 37204 25596 37256
rect 25648 37204 25654 37256
rect 26786 37244 26792 37256
rect 26747 37216 26792 37244
rect 26786 37204 26792 37216
rect 26844 37204 26850 37256
rect 30745 37247 30803 37253
rect 30745 37213 30757 37247
rect 30791 37244 30803 37247
rect 31018 37244 31024 37256
rect 30791 37216 31024 37244
rect 30791 37213 30803 37216
rect 30745 37207 30803 37213
rect 31018 37204 31024 37216
rect 31076 37204 31082 37256
rect 46293 37247 46351 37253
rect 46293 37213 46305 37247
rect 46339 37213 46351 37247
rect 46293 37207 46351 37213
rect 19444 37148 22094 37176
rect 25225 37179 25283 37185
rect 25225 37145 25237 37179
rect 25271 37176 25283 37179
rect 25866 37176 25872 37188
rect 25271 37148 25872 37176
rect 25271 37145 25283 37148
rect 25225 37139 25283 37145
rect 25866 37136 25872 37148
rect 25924 37136 25930 37188
rect 27525 37179 27583 37185
rect 27525 37145 27537 37179
rect 27571 37145 27583 37179
rect 29270 37176 29276 37188
rect 28750 37148 29276 37176
rect 27525 37139 27583 37145
rect 21910 37108 21916 37120
rect 21871 37080 21916 37108
rect 21910 37068 21916 37080
rect 21968 37068 21974 37120
rect 24673 37111 24731 37117
rect 24673 37077 24685 37111
rect 24719 37108 24731 37111
rect 24854 37108 24860 37120
rect 24719 37080 24860 37108
rect 24719 37077 24731 37080
rect 24673 37071 24731 37077
rect 24854 37068 24860 37080
rect 24912 37068 24918 37120
rect 25406 37068 25412 37120
rect 25464 37108 25470 37120
rect 25685 37111 25743 37117
rect 25685 37108 25697 37111
rect 25464 37080 25697 37108
rect 25464 37068 25470 37080
rect 25685 37077 25697 37080
rect 25731 37077 25743 37111
rect 25685 37071 25743 37077
rect 26605 37111 26663 37117
rect 26605 37077 26617 37111
rect 26651 37108 26663 37111
rect 27540 37108 27568 37139
rect 29270 37136 29276 37148
rect 29328 37136 29334 37188
rect 26651 37080 27568 37108
rect 26651 37077 26663 37080
rect 26605 37071 26663 37077
rect 28350 37068 28356 37120
rect 28408 37108 28414 37120
rect 28997 37111 29055 37117
rect 28997 37108 29009 37111
rect 28408 37080 29009 37108
rect 28408 37068 28414 37080
rect 28997 37077 29009 37080
rect 29043 37077 29055 37111
rect 30834 37108 30840 37120
rect 30795 37080 30840 37108
rect 28997 37071 29055 37077
rect 30834 37068 30840 37080
rect 30892 37068 30898 37120
rect 46308 37108 46336 37207
rect 46477 37179 46535 37185
rect 46477 37145 46489 37179
rect 46523 37176 46535 37179
rect 47670 37176 47676 37188
rect 46523 37148 47676 37176
rect 46523 37145 46535 37148
rect 46477 37139 46535 37145
rect 47670 37136 47676 37148
rect 47728 37136 47734 37188
rect 46934 37108 46940 37120
rect 46308 37080 46940 37108
rect 46934 37068 46940 37080
rect 46992 37068 46998 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 24946 36904 24952 36916
rect 24907 36876 24952 36904
rect 24946 36864 24952 36876
rect 25004 36864 25010 36916
rect 25682 36904 25688 36916
rect 25332 36876 25688 36904
rect 11790 36796 11796 36848
rect 11848 36836 11854 36848
rect 25222 36836 25228 36848
rect 11848 36808 22324 36836
rect 11848 36796 11854 36808
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 22296 36777 22324 36808
rect 24504 36808 25228 36836
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 22189 36771 22247 36777
rect 22189 36737 22201 36771
rect 22235 36737 22247 36771
rect 22189 36731 22247 36737
rect 22281 36771 22339 36777
rect 22281 36737 22293 36771
rect 22327 36737 22339 36771
rect 22281 36731 22339 36737
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 22020 36632 22048 36731
rect 22204 36700 22232 36731
rect 24504 36700 24532 36808
rect 25222 36796 25228 36808
rect 25280 36796 25286 36848
rect 24670 36768 24676 36780
rect 24631 36740 24676 36768
rect 24670 36728 24676 36740
rect 24728 36728 24734 36780
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36768 24823 36771
rect 25332 36768 25360 36876
rect 25682 36864 25688 36876
rect 25740 36864 25746 36916
rect 25774 36864 25780 36916
rect 25832 36904 25838 36916
rect 26053 36907 26111 36913
rect 26053 36904 26065 36907
rect 25832 36876 26065 36904
rect 25832 36864 25838 36876
rect 26053 36873 26065 36876
rect 26099 36873 26111 36907
rect 26053 36867 26111 36873
rect 27065 36907 27123 36913
rect 27065 36873 27077 36907
rect 27111 36904 27123 36907
rect 27246 36904 27252 36916
rect 27111 36876 27252 36904
rect 27111 36873 27123 36876
rect 27065 36867 27123 36873
rect 27246 36864 27252 36876
rect 27304 36864 27310 36916
rect 27433 36907 27491 36913
rect 27433 36873 27445 36907
rect 27479 36904 27491 36907
rect 27982 36904 27988 36916
rect 27479 36876 27988 36904
rect 27479 36873 27491 36876
rect 27433 36867 27491 36873
rect 27982 36864 27988 36876
rect 28040 36904 28046 36916
rect 28718 36904 28724 36916
rect 28040 36876 28724 36904
rect 28040 36864 28046 36876
rect 28718 36864 28724 36876
rect 28776 36864 28782 36916
rect 25409 36839 25467 36845
rect 25409 36805 25421 36839
rect 25455 36836 25467 36839
rect 26234 36836 26240 36848
rect 25455 36808 26240 36836
rect 25455 36805 25467 36808
rect 25409 36799 25467 36805
rect 26234 36796 26240 36808
rect 26292 36796 26298 36848
rect 30834 36796 30840 36848
rect 30892 36796 30898 36848
rect 25869 36771 25927 36777
rect 25869 36768 25881 36771
rect 24811 36740 25360 36768
rect 25516 36740 25881 36768
rect 24811 36737 24823 36740
rect 24765 36731 24823 36737
rect 22204 36672 24532 36700
rect 24949 36703 25007 36709
rect 24949 36669 24961 36703
rect 24995 36700 25007 36703
rect 25516 36700 25544 36740
rect 25869 36737 25881 36740
rect 25915 36768 25927 36771
rect 26142 36768 26148 36780
rect 25915 36740 26148 36768
rect 25915 36737 25927 36740
rect 25869 36731 25927 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 27246 36768 27252 36780
rect 27207 36740 27252 36768
rect 27246 36728 27252 36740
rect 27304 36728 27310 36780
rect 27522 36768 27528 36780
rect 27483 36740 27528 36768
rect 27522 36728 27528 36740
rect 27580 36728 27586 36780
rect 24995 36672 25544 36700
rect 24995 36669 25007 36672
rect 24949 36663 25007 36669
rect 25682 36660 25688 36712
rect 25740 36700 25746 36712
rect 25740 36672 25785 36700
rect 25740 36660 25746 36672
rect 25958 36660 25964 36712
rect 26016 36700 26022 36712
rect 26016 36672 28028 36700
rect 26016 36660 26022 36672
rect 24854 36632 24860 36644
rect 22020 36604 24860 36632
rect 24854 36592 24860 36604
rect 24912 36592 24918 36644
rect 27706 36632 27712 36644
rect 25700 36604 27712 36632
rect 21174 36524 21180 36576
rect 21232 36564 21238 36576
rect 21821 36567 21879 36573
rect 21821 36564 21833 36567
rect 21232 36536 21833 36564
rect 21232 36524 21238 36536
rect 21821 36533 21833 36536
rect 21867 36533 21879 36567
rect 21821 36527 21879 36533
rect 22370 36524 22376 36576
rect 22428 36564 22434 36576
rect 25700 36564 25728 36604
rect 27706 36592 27712 36604
rect 27764 36592 27770 36644
rect 22428 36536 25728 36564
rect 25869 36567 25927 36573
rect 22428 36524 22434 36536
rect 25869 36533 25881 36567
rect 25915 36564 25927 36567
rect 27890 36564 27896 36576
rect 25915 36536 27896 36564
rect 25915 36533 25927 36536
rect 25869 36527 25927 36533
rect 27890 36524 27896 36536
rect 27948 36524 27954 36576
rect 28000 36564 28028 36672
rect 28994 36660 29000 36712
rect 29052 36700 29058 36712
rect 29549 36703 29607 36709
rect 29549 36700 29561 36703
rect 29052 36672 29561 36700
rect 29052 36660 29058 36672
rect 29549 36669 29561 36672
rect 29595 36669 29607 36703
rect 29822 36700 29828 36712
rect 29783 36672 29828 36700
rect 29549 36663 29607 36669
rect 29822 36660 29828 36672
rect 29880 36660 29886 36712
rect 31110 36564 31116 36576
rect 28000 36536 31116 36564
rect 31110 36524 31116 36536
rect 31168 36524 31174 36576
rect 31294 36564 31300 36576
rect 31255 36536 31300 36564
rect 31294 36524 31300 36536
rect 31352 36524 31358 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 9490 36320 9496 36372
rect 9548 36360 9554 36372
rect 26418 36360 26424 36372
rect 9548 36332 26096 36360
rect 26379 36332 26424 36360
rect 9548 36320 9554 36332
rect 23661 36295 23719 36301
rect 23661 36261 23673 36295
rect 23707 36261 23719 36295
rect 23661 36255 23719 36261
rect 19150 36184 19156 36236
rect 19208 36224 19214 36236
rect 20901 36227 20959 36233
rect 20901 36224 20913 36227
rect 19208 36196 20913 36224
rect 19208 36184 19214 36196
rect 20901 36193 20913 36196
rect 20947 36224 20959 36227
rect 22186 36224 22192 36236
rect 20947 36196 22192 36224
rect 20947 36193 20959 36196
rect 20901 36187 20959 36193
rect 22186 36184 22192 36196
rect 22244 36184 22250 36236
rect 23382 36224 23388 36236
rect 23343 36196 23388 36224
rect 23382 36184 23388 36196
rect 23440 36184 23446 36236
rect 2130 36156 2136 36168
rect 2043 36128 2136 36156
rect 2130 36116 2136 36128
rect 2188 36156 2194 36168
rect 2188 36128 6914 36156
rect 2188 36116 2194 36128
rect 6886 36088 6914 36128
rect 19334 36116 19340 36168
rect 19392 36156 19398 36168
rect 19889 36159 19947 36165
rect 19889 36156 19901 36159
rect 19392 36128 19901 36156
rect 19392 36116 19398 36128
rect 19889 36125 19901 36128
rect 19935 36156 19947 36159
rect 19978 36156 19984 36168
rect 19935 36128 19984 36156
rect 19935 36125 19947 36128
rect 19889 36119 19947 36125
rect 19978 36116 19984 36128
rect 20036 36116 20042 36168
rect 23293 36159 23351 36165
rect 23293 36125 23305 36159
rect 23339 36125 23351 36159
rect 23676 36156 23704 36255
rect 24670 36252 24676 36304
rect 24728 36252 24734 36304
rect 24854 36252 24860 36304
rect 24912 36292 24918 36304
rect 24949 36295 25007 36301
rect 24949 36292 24961 36295
rect 24912 36264 24961 36292
rect 24912 36252 24918 36264
rect 24949 36261 24961 36264
rect 24995 36261 25007 36295
rect 25958 36292 25964 36304
rect 24949 36255 25007 36261
rect 25056 36264 25964 36292
rect 24688 36224 24716 36252
rect 24688 36196 24808 36224
rect 24780 36165 24808 36196
rect 24397 36159 24455 36165
rect 24397 36156 24409 36159
rect 23676 36128 24409 36156
rect 23293 36119 23351 36125
rect 24397 36125 24409 36128
rect 24443 36125 24455 36159
rect 24673 36159 24731 36165
rect 24673 36156 24685 36159
rect 24397 36119 24455 36125
rect 24504 36128 24685 36156
rect 19426 36088 19432 36100
rect 6886 36060 19432 36088
rect 19426 36048 19432 36060
rect 19484 36048 19490 36100
rect 21174 36088 21180 36100
rect 21135 36060 21180 36088
rect 21174 36048 21180 36060
rect 21232 36048 21238 36100
rect 21910 36048 21916 36100
rect 21968 36048 21974 36100
rect 22922 36088 22928 36100
rect 22664 36060 22928 36088
rect 19978 36020 19984 36032
rect 19939 35992 19984 36020
rect 19978 35980 19984 35992
rect 20036 35980 20042 36032
rect 22664 36029 22692 36060
rect 22922 36048 22928 36060
rect 22980 36088 22986 36100
rect 23308 36088 23336 36119
rect 24504 36088 24532 36128
rect 24673 36125 24685 36128
rect 24719 36125 24731 36159
rect 24673 36119 24731 36125
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36156 24823 36159
rect 25056 36156 25084 36264
rect 25958 36252 25964 36264
rect 26016 36252 26022 36304
rect 25222 36184 25228 36236
rect 25280 36224 25286 36236
rect 26068 36224 26096 36332
rect 26418 36320 26424 36332
rect 26476 36320 26482 36372
rect 26786 36320 26792 36372
rect 26844 36360 26850 36372
rect 27617 36363 27675 36369
rect 27617 36360 27629 36363
rect 26844 36332 27629 36360
rect 26844 36320 26850 36332
rect 27617 36329 27629 36332
rect 27663 36329 27675 36363
rect 27617 36323 27675 36329
rect 27706 36320 27712 36372
rect 27764 36360 27770 36372
rect 29549 36363 29607 36369
rect 27764 36332 28212 36360
rect 27764 36320 27770 36332
rect 27525 36295 27583 36301
rect 27525 36261 27537 36295
rect 27571 36292 27583 36295
rect 28074 36292 28080 36304
rect 27571 36264 28080 36292
rect 27571 36261 27583 36264
rect 27525 36255 27583 36261
rect 28074 36252 28080 36264
rect 28132 36252 28138 36304
rect 28184 36292 28212 36332
rect 29549 36329 29561 36363
rect 29595 36360 29607 36363
rect 29822 36360 29828 36372
rect 29595 36332 29828 36360
rect 29595 36329 29607 36332
rect 29549 36323 29607 36329
rect 29822 36320 29828 36332
rect 29880 36320 29886 36372
rect 28184 36264 30144 36292
rect 30009 36227 30067 36233
rect 30009 36224 30021 36227
rect 25280 36196 26004 36224
rect 26068 36196 30021 36224
rect 25280 36184 25286 36196
rect 25406 36156 25412 36168
rect 24811 36128 25084 36156
rect 25367 36128 25412 36156
rect 24811 36125 24823 36128
rect 24765 36119 24823 36125
rect 25406 36116 25412 36128
rect 25464 36116 25470 36168
rect 22980 36060 24532 36088
rect 24581 36091 24639 36097
rect 22980 36048 22986 36060
rect 24581 36057 24593 36091
rect 24627 36088 24639 36091
rect 25498 36088 25504 36100
rect 24627 36060 25504 36088
rect 24627 36057 24639 36060
rect 24581 36051 24639 36057
rect 25498 36048 25504 36060
rect 25556 36048 25562 36100
rect 25593 36091 25651 36097
rect 25593 36057 25605 36091
rect 25639 36088 25651 36091
rect 25682 36088 25688 36100
rect 25639 36060 25688 36088
rect 25639 36057 25651 36060
rect 25593 36051 25651 36057
rect 25682 36048 25688 36060
rect 25740 36048 25746 36100
rect 25976 36088 26004 36196
rect 30009 36193 30021 36196
rect 30055 36193 30067 36227
rect 30009 36187 30067 36193
rect 26234 36156 26240 36168
rect 26195 36128 26240 36156
rect 26234 36116 26240 36128
rect 26292 36116 26298 36168
rect 27982 36156 27988 36168
rect 26988 36128 27988 36156
rect 26878 36088 26884 36100
rect 25976 36060 26884 36088
rect 26878 36048 26884 36060
rect 26936 36048 26942 36100
rect 22649 36023 22707 36029
rect 22649 35989 22661 36023
rect 22695 35989 22707 36023
rect 22649 35983 22707 35989
rect 23566 35980 23572 36032
rect 23624 36020 23630 36032
rect 25777 36023 25835 36029
rect 25777 36020 25789 36023
rect 23624 35992 25789 36020
rect 23624 35980 23630 35992
rect 25777 35989 25789 35992
rect 25823 35989 25835 36023
rect 25777 35983 25835 35989
rect 25866 35980 25872 36032
rect 25924 36020 25930 36032
rect 26988 36020 27016 36128
rect 27982 36116 27988 36128
rect 28040 36156 28046 36168
rect 28077 36159 28135 36165
rect 28077 36156 28089 36159
rect 28040 36128 28089 36156
rect 28040 36116 28046 36128
rect 28077 36125 28089 36128
rect 28123 36125 28135 36159
rect 28077 36119 28135 36125
rect 29733 36159 29791 36165
rect 29733 36125 29745 36159
rect 29779 36125 29791 36159
rect 29733 36119 29791 36125
rect 27157 36091 27215 36097
rect 27157 36057 27169 36091
rect 27203 36088 27215 36091
rect 28534 36088 28540 36100
rect 27203 36060 28540 36088
rect 27203 36057 27215 36060
rect 27157 36051 27215 36057
rect 28534 36048 28540 36060
rect 28592 36048 28598 36100
rect 29748 36088 29776 36119
rect 29822 36116 29828 36168
rect 29880 36156 29886 36168
rect 30116 36165 30144 36264
rect 30561 36227 30619 36233
rect 30561 36193 30573 36227
rect 30607 36224 30619 36227
rect 31294 36224 31300 36236
rect 30607 36196 31300 36224
rect 30607 36193 30619 36196
rect 30561 36187 30619 36193
rect 31294 36184 31300 36196
rect 31352 36184 31358 36236
rect 30101 36159 30159 36165
rect 29880 36128 29925 36156
rect 29880 36116 29886 36128
rect 30101 36125 30113 36159
rect 30147 36125 30159 36159
rect 30101 36119 30159 36125
rect 30745 36159 30803 36165
rect 30745 36125 30757 36159
rect 30791 36156 30803 36159
rect 30834 36156 30840 36168
rect 30791 36128 30840 36156
rect 30791 36125 30803 36128
rect 30745 36119 30803 36125
rect 30834 36116 30840 36128
rect 30892 36116 30898 36168
rect 31018 36116 31024 36168
rect 31076 36156 31082 36168
rect 32033 36159 32091 36165
rect 32033 36156 32045 36159
rect 31076 36128 32045 36156
rect 31076 36116 31082 36128
rect 32033 36125 32045 36128
rect 32079 36125 32091 36159
rect 32033 36119 32091 36125
rect 30929 36091 30987 36097
rect 30929 36088 30941 36091
rect 29748 36060 30941 36088
rect 30929 36057 30941 36060
rect 30975 36057 30987 36091
rect 30929 36051 30987 36057
rect 25924 35992 27016 36020
rect 25924 35980 25930 35992
rect 27430 35980 27436 36032
rect 27488 36020 27494 36032
rect 28169 36023 28227 36029
rect 28169 36020 28181 36023
rect 27488 35992 28181 36020
rect 27488 35980 27494 35992
rect 28169 35989 28181 35992
rect 28215 35989 28227 36023
rect 28169 35983 28227 35989
rect 32125 36023 32183 36029
rect 32125 35989 32137 36023
rect 32171 36020 32183 36023
rect 33134 36020 33140 36032
rect 32171 35992 33140 36020
rect 32171 35989 32183 35992
rect 32125 35983 32183 35989
rect 33134 35980 33140 35992
rect 33192 35980 33198 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 22557 35819 22615 35825
rect 22557 35816 22569 35819
rect 19444 35788 22569 35816
rect 19444 35757 19472 35788
rect 22557 35785 22569 35788
rect 22603 35785 22615 35819
rect 22557 35779 22615 35785
rect 27709 35819 27767 35825
rect 27709 35785 27721 35819
rect 27755 35816 27767 35819
rect 28369 35819 28427 35825
rect 28369 35816 28381 35819
rect 27755 35788 28381 35816
rect 27755 35785 27767 35788
rect 27709 35779 27767 35785
rect 28369 35785 28381 35788
rect 28415 35785 28427 35819
rect 28534 35816 28540 35828
rect 28495 35788 28540 35816
rect 28369 35779 28427 35785
rect 28534 35776 28540 35788
rect 28592 35776 28598 35828
rect 29733 35819 29791 35825
rect 29733 35785 29745 35819
rect 29779 35816 29791 35819
rect 29822 35816 29828 35828
rect 29779 35788 29828 35816
rect 29779 35785 29791 35788
rect 29733 35779 29791 35785
rect 29822 35776 29828 35788
rect 29880 35776 29886 35828
rect 29917 35819 29975 35825
rect 29917 35785 29929 35819
rect 29963 35816 29975 35819
rect 30926 35816 30932 35828
rect 29963 35788 30932 35816
rect 29963 35785 29975 35788
rect 29917 35779 29975 35785
rect 30926 35776 30932 35788
rect 30984 35816 30990 35828
rect 31205 35819 31263 35825
rect 31205 35816 31217 35819
rect 30984 35788 31217 35816
rect 30984 35776 30990 35788
rect 31205 35785 31217 35788
rect 31251 35785 31263 35819
rect 31205 35779 31263 35785
rect 19429 35751 19487 35757
rect 19429 35717 19441 35751
rect 19475 35717 19487 35751
rect 19429 35711 19487 35717
rect 19978 35708 19984 35760
rect 20036 35708 20042 35760
rect 21542 35708 21548 35760
rect 21600 35748 21606 35760
rect 26970 35748 26976 35760
rect 21600 35720 26976 35748
rect 21600 35708 21606 35720
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 21818 35680 21824 35692
rect 21779 35652 21824 35680
rect 21818 35640 21824 35652
rect 21876 35640 21882 35692
rect 22020 35689 22048 35720
rect 26970 35708 26976 35720
rect 27028 35708 27034 35760
rect 27065 35751 27123 35757
rect 27065 35717 27077 35751
rect 27111 35748 27123 35751
rect 28166 35748 28172 35760
rect 27111 35720 27844 35748
rect 28127 35720 28172 35748
rect 27111 35717 27123 35720
rect 27065 35711 27123 35717
rect 22005 35683 22063 35689
rect 22005 35649 22017 35683
rect 22051 35649 22063 35683
rect 22005 35643 22063 35649
rect 22189 35683 22247 35689
rect 22189 35649 22201 35683
rect 22235 35680 22247 35683
rect 22278 35680 22284 35692
rect 22235 35652 22284 35680
rect 22235 35649 22247 35652
rect 22189 35643 22247 35649
rect 22278 35640 22284 35652
rect 22336 35640 22342 35692
rect 22370 35640 22376 35692
rect 22428 35680 22434 35692
rect 22830 35680 22836 35692
rect 22428 35652 22836 35680
rect 22428 35640 22434 35652
rect 22830 35640 22836 35652
rect 22888 35640 22894 35692
rect 23201 35683 23259 35689
rect 23201 35649 23213 35683
rect 23247 35649 23259 35683
rect 23201 35643 23259 35649
rect 23385 35683 23443 35689
rect 23385 35649 23397 35683
rect 23431 35680 23443 35683
rect 23566 35680 23572 35692
rect 23431 35652 23572 35680
rect 23431 35649 23443 35652
rect 23385 35643 23443 35649
rect 18598 35572 18604 35624
rect 18656 35612 18662 35624
rect 19150 35612 19156 35624
rect 18656 35584 19156 35612
rect 18656 35572 18662 35584
rect 19150 35572 19156 35584
rect 19208 35572 19214 35624
rect 20901 35615 20959 35621
rect 20901 35581 20913 35615
rect 20947 35612 20959 35615
rect 22097 35615 22155 35621
rect 22097 35612 22109 35615
rect 20947 35584 22109 35612
rect 20947 35581 20959 35584
rect 20901 35575 20959 35581
rect 22097 35581 22109 35584
rect 22143 35612 22155 35615
rect 22646 35612 22652 35624
rect 22143 35584 22652 35612
rect 22143 35581 22155 35584
rect 22097 35575 22155 35581
rect 22646 35572 22652 35584
rect 22704 35612 22710 35624
rect 23216 35612 23244 35643
rect 23566 35640 23572 35652
rect 23624 35640 23630 35692
rect 24581 35683 24639 35689
rect 24581 35649 24593 35683
rect 24627 35649 24639 35683
rect 24581 35643 24639 35649
rect 25225 35683 25283 35689
rect 25225 35649 25237 35683
rect 25271 35680 25283 35683
rect 25501 35683 25559 35689
rect 25271 35652 25452 35680
rect 25271 35649 25283 35652
rect 25225 35643 25283 35649
rect 22704 35584 23244 35612
rect 23477 35615 23535 35621
rect 22704 35572 22710 35584
rect 23477 35581 23489 35615
rect 23523 35581 23535 35615
rect 24596 35612 24624 35643
rect 24762 35612 24768 35624
rect 24596 35584 24768 35612
rect 23477 35575 23535 35581
rect 21634 35504 21640 35556
rect 21692 35544 21698 35556
rect 23017 35547 23075 35553
rect 23017 35544 23029 35547
rect 21692 35516 23029 35544
rect 21692 35504 21698 35516
rect 23017 35513 23029 35516
rect 23063 35513 23075 35547
rect 23492 35544 23520 35575
rect 24762 35572 24768 35584
rect 24820 35612 24826 35624
rect 25317 35615 25375 35621
rect 25317 35612 25329 35615
rect 24820 35584 25329 35612
rect 24820 35572 24826 35584
rect 25317 35581 25329 35584
rect 25363 35581 25375 35615
rect 25424 35612 25452 35652
rect 25501 35649 25513 35683
rect 25547 35680 25559 35683
rect 25590 35680 25596 35692
rect 25547 35652 25596 35680
rect 25547 35649 25559 35652
rect 25501 35643 25559 35649
rect 25590 35640 25596 35652
rect 25648 35680 25654 35692
rect 27080 35680 27108 35711
rect 27430 35680 27436 35692
rect 25648 35652 27108 35680
rect 27391 35652 27436 35680
rect 25648 35640 25654 35652
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 27816 35680 27844 35720
rect 28166 35708 28172 35720
rect 28224 35708 28230 35760
rect 31021 35751 31079 35757
rect 31021 35748 31033 35751
rect 30392 35720 31033 35748
rect 30392 35692 30420 35720
rect 31021 35717 31033 35720
rect 31067 35748 31079 35751
rect 31294 35748 31300 35760
rect 31067 35720 31300 35748
rect 31067 35717 31079 35720
rect 31021 35711 31079 35717
rect 31294 35708 31300 35720
rect 31352 35708 31358 35760
rect 33134 35708 33140 35760
rect 33192 35708 33198 35760
rect 28350 35680 28356 35692
rect 27816 35652 28356 35680
rect 28350 35640 28356 35652
rect 28408 35640 28414 35692
rect 29454 35640 29460 35692
rect 29512 35680 29518 35692
rect 29858 35683 29916 35689
rect 29858 35680 29870 35683
rect 29512 35652 29870 35680
rect 29512 35640 29518 35652
rect 29858 35649 29870 35652
rect 29904 35649 29916 35683
rect 30374 35680 30380 35692
rect 30287 35652 30380 35680
rect 29858 35643 29916 35649
rect 30374 35640 30380 35652
rect 30432 35640 30438 35692
rect 30834 35680 30840 35692
rect 30795 35652 30840 35680
rect 30834 35640 30840 35652
rect 30892 35640 30898 35692
rect 48130 35680 48136 35692
rect 48091 35652 48136 35680
rect 48130 35640 48136 35652
rect 48188 35640 48194 35692
rect 25682 35612 25688 35624
rect 25424 35584 25688 35612
rect 25317 35575 25375 35581
rect 25682 35572 25688 35584
rect 25740 35612 25746 35624
rect 25740 35584 26004 35612
rect 25740 35572 25746 35584
rect 25866 35544 25872 35556
rect 23492 35516 24716 35544
rect 23017 35507 23075 35513
rect 24688 35488 24716 35516
rect 25516 35516 25872 35544
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 2222 35476 2228 35488
rect 1443 35448 2228 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 2222 35436 2228 35448
rect 2280 35436 2286 35488
rect 24670 35476 24676 35488
rect 24631 35448 24676 35476
rect 24670 35436 24676 35448
rect 24728 35436 24734 35488
rect 25516 35485 25544 35516
rect 25866 35504 25872 35516
rect 25924 35504 25930 35556
rect 25976 35544 26004 35584
rect 27154 35572 27160 35624
rect 27212 35612 27218 35624
rect 27525 35615 27583 35621
rect 27525 35612 27537 35615
rect 27212 35584 27537 35612
rect 27212 35572 27218 35584
rect 27525 35581 27537 35584
rect 27571 35581 27583 35615
rect 29086 35612 29092 35624
rect 27525 35575 27583 35581
rect 27724 35584 29092 35612
rect 27724 35544 27752 35584
rect 29086 35572 29092 35584
rect 29144 35572 29150 35624
rect 32122 35612 32128 35624
rect 32083 35584 32128 35612
rect 32122 35572 32128 35584
rect 32180 35572 32186 35624
rect 32401 35615 32459 35621
rect 32401 35581 32413 35615
rect 32447 35612 32459 35615
rect 32490 35612 32496 35624
rect 32447 35584 32496 35612
rect 32447 35581 32459 35584
rect 32401 35575 32459 35581
rect 32490 35572 32496 35584
rect 32548 35572 32554 35624
rect 25976 35516 27752 35544
rect 28258 35504 28264 35556
rect 28316 35544 28322 35556
rect 30285 35547 30343 35553
rect 30285 35544 30297 35547
rect 28316 35516 30297 35544
rect 28316 35504 28322 35516
rect 30285 35513 30297 35516
rect 30331 35513 30343 35547
rect 30285 35507 30343 35513
rect 25501 35479 25559 35485
rect 25501 35445 25513 35479
rect 25547 35445 25559 35479
rect 25501 35439 25559 35445
rect 25685 35479 25743 35485
rect 25685 35445 25697 35479
rect 25731 35476 25743 35479
rect 25774 35476 25780 35488
rect 25731 35448 25780 35476
rect 25731 35445 25743 35448
rect 25685 35439 25743 35445
rect 25774 35436 25780 35448
rect 25832 35476 25838 35488
rect 28353 35479 28411 35485
rect 28353 35476 28365 35479
rect 25832 35448 28365 35476
rect 25832 35436 25838 35448
rect 28353 35445 28365 35448
rect 28399 35445 28411 35479
rect 28353 35439 28411 35445
rect 31018 35436 31024 35488
rect 31076 35476 31082 35488
rect 32030 35476 32036 35488
rect 31076 35448 32036 35476
rect 31076 35436 31082 35448
rect 32030 35436 32036 35448
rect 32088 35476 32094 35488
rect 33873 35479 33931 35485
rect 33873 35476 33885 35479
rect 32088 35448 33885 35476
rect 32088 35436 32094 35448
rect 33873 35445 33885 35448
rect 33919 35445 33931 35479
rect 33873 35439 33931 35445
rect 47118 35436 47124 35488
rect 47176 35476 47182 35488
rect 47949 35479 48007 35485
rect 47949 35476 47961 35479
rect 47176 35448 47961 35476
rect 47176 35436 47182 35448
rect 47949 35445 47961 35448
rect 47995 35445 48007 35479
rect 47949 35439 48007 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 21634 35272 21640 35284
rect 21595 35244 21640 35272
rect 21634 35232 21640 35244
rect 21692 35232 21698 35284
rect 21818 35272 21824 35284
rect 21779 35244 21824 35272
rect 21818 35232 21824 35244
rect 21876 35232 21882 35284
rect 22554 35232 22560 35284
rect 22612 35272 22618 35284
rect 22649 35275 22707 35281
rect 22649 35272 22661 35275
rect 22612 35244 22661 35272
rect 22612 35232 22618 35244
rect 22649 35241 22661 35244
rect 22695 35272 22707 35275
rect 23382 35272 23388 35284
rect 22695 35244 23388 35272
rect 22695 35241 22707 35244
rect 22649 35235 22707 35241
rect 23382 35232 23388 35244
rect 23440 35272 23446 35284
rect 24578 35272 24584 35284
rect 23440 35244 24584 35272
rect 23440 35232 23446 35244
rect 24578 35232 24584 35244
rect 24636 35232 24642 35284
rect 24762 35272 24768 35284
rect 24723 35244 24768 35272
rect 24762 35232 24768 35244
rect 24820 35232 24826 35284
rect 26973 35275 27031 35281
rect 26973 35241 26985 35275
rect 27019 35272 27031 35275
rect 27246 35272 27252 35284
rect 27019 35244 27252 35272
rect 27019 35241 27031 35244
rect 26973 35235 27031 35241
rect 27246 35232 27252 35244
rect 27304 35232 27310 35284
rect 28074 35272 28080 35284
rect 28035 35244 28080 35272
rect 28074 35232 28080 35244
rect 28132 35232 28138 35284
rect 28534 35272 28540 35284
rect 28495 35244 28540 35272
rect 28534 35232 28540 35244
rect 28592 35232 28598 35284
rect 28902 35232 28908 35284
rect 28960 35272 28966 35284
rect 31846 35272 31852 35284
rect 28960 35244 31852 35272
rect 28960 35232 28966 35244
rect 31846 35232 31852 35244
rect 31904 35232 31910 35284
rect 32490 35272 32496 35284
rect 32451 35244 32496 35272
rect 32490 35232 32496 35244
rect 32548 35232 32554 35284
rect 25498 35164 25504 35216
rect 25556 35204 25562 35216
rect 26421 35207 26479 35213
rect 26421 35204 26433 35207
rect 25556 35176 26433 35204
rect 25556 35164 25562 35176
rect 26421 35173 26433 35176
rect 26467 35204 26479 35207
rect 26467 35176 27292 35204
rect 26467 35173 26479 35176
rect 26421 35167 26479 35173
rect 22557 35139 22615 35145
rect 22557 35105 22569 35139
rect 22603 35136 22615 35139
rect 23474 35136 23480 35148
rect 22603 35108 23480 35136
rect 22603 35105 22615 35108
rect 22557 35099 22615 35105
rect 23474 35096 23480 35108
rect 23532 35136 23538 35148
rect 27264 35136 27292 35176
rect 28718 35164 28724 35216
rect 28776 35204 28782 35216
rect 31938 35204 31944 35216
rect 28776 35176 31944 35204
rect 28776 35164 28782 35176
rect 31938 35164 31944 35176
rect 31996 35164 32002 35216
rect 27798 35136 27804 35148
rect 23532 35108 24440 35136
rect 23532 35096 23538 35108
rect 20346 35028 20352 35080
rect 20404 35068 20410 35080
rect 21269 35071 21327 35077
rect 21269 35068 21281 35071
rect 20404 35040 21281 35068
rect 20404 35028 20410 35040
rect 21269 35037 21281 35040
rect 21315 35037 21327 35071
rect 21269 35031 21327 35037
rect 21637 35071 21695 35077
rect 21637 35037 21649 35071
rect 21683 35068 21695 35071
rect 22094 35068 22100 35080
rect 21683 35040 22100 35068
rect 21683 35037 21695 35040
rect 21637 35031 21695 35037
rect 22094 35028 22100 35040
rect 22152 35028 22158 35080
rect 22646 35068 22652 35080
rect 22607 35040 22652 35068
rect 22646 35028 22652 35040
rect 22704 35028 22710 35080
rect 24412 35077 24440 35108
rect 27264 35108 27804 35136
rect 24397 35071 24455 35077
rect 24397 35037 24409 35071
rect 24443 35037 24455 35071
rect 24397 35031 24455 35037
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35068 26295 35071
rect 26326 35068 26332 35080
rect 26283 35040 26332 35068
rect 26283 35037 26295 35040
rect 26237 35031 26295 35037
rect 26326 35028 26332 35040
rect 26384 35028 26390 35080
rect 27154 35068 27160 35080
rect 27115 35040 27160 35068
rect 27154 35028 27160 35040
rect 27212 35028 27218 35080
rect 27264 35077 27292 35108
rect 27798 35096 27804 35108
rect 27856 35096 27862 35148
rect 30745 35139 30803 35145
rect 30745 35105 30757 35139
rect 30791 35136 30803 35139
rect 32030 35136 32036 35148
rect 30791 35108 31800 35136
rect 31991 35108 32036 35136
rect 30791 35105 30803 35108
rect 30745 35099 30803 35105
rect 27249 35071 27307 35077
rect 27249 35037 27261 35071
rect 27295 35037 27307 35071
rect 27249 35031 27307 35037
rect 27617 35071 27675 35077
rect 27617 35037 27629 35071
rect 27663 35068 27675 35071
rect 27890 35068 27896 35080
rect 27663 35040 27896 35068
rect 27663 35037 27675 35040
rect 27617 35031 27675 35037
rect 27890 35028 27896 35040
rect 27948 35028 27954 35080
rect 28258 35068 28264 35080
rect 28219 35040 28264 35068
rect 28258 35028 28264 35040
rect 28316 35028 28322 35080
rect 28350 35028 28356 35080
rect 28408 35068 28414 35080
rect 28626 35068 28632 35080
rect 28408 35040 28453 35068
rect 28587 35040 28632 35068
rect 28408 35028 28414 35040
rect 28626 35028 28632 35040
rect 28684 35028 28690 35080
rect 29086 35028 29092 35080
rect 29144 35068 29150 35080
rect 29917 35071 29975 35077
rect 29917 35068 29929 35071
rect 29144 35040 29929 35068
rect 29144 35028 29150 35040
rect 29917 35037 29929 35040
rect 29963 35037 29975 35071
rect 30098 35068 30104 35080
rect 30059 35040 30104 35068
rect 29917 35031 29975 35037
rect 22373 35003 22431 35009
rect 22373 34969 22385 35003
rect 22419 35000 22431 35003
rect 23566 35000 23572 35012
rect 22419 34972 23572 35000
rect 22419 34969 22431 34972
rect 22373 34963 22431 34969
rect 23566 34960 23572 34972
rect 23624 34960 23630 35012
rect 24578 35000 24584 35012
rect 24539 34972 24584 35000
rect 24578 34960 24584 34972
rect 24636 34960 24642 35012
rect 27338 35000 27344 35012
rect 27300 34972 27344 35000
rect 27338 34960 27344 34972
rect 27396 34960 27402 35012
rect 27430 34960 27436 35012
rect 27488 35009 27494 35012
rect 27488 35003 27517 35009
rect 27505 34969 27517 35003
rect 29932 35000 29960 35031
rect 30098 35028 30104 35040
rect 30156 35028 30162 35080
rect 30926 35068 30932 35080
rect 30887 35040 30932 35068
rect 30926 35028 30932 35040
rect 30984 35028 30990 35080
rect 31018 35028 31024 35080
rect 31076 35068 31082 35080
rect 31205 35071 31263 35077
rect 31076 35040 31121 35068
rect 31076 35028 31082 35040
rect 31205 35037 31217 35071
rect 31251 35037 31263 35071
rect 31205 35031 31263 35037
rect 31297 35071 31355 35077
rect 31297 35037 31309 35071
rect 31343 35068 31355 35071
rect 31662 35068 31668 35080
rect 31343 35040 31668 35068
rect 31343 35037 31355 35040
rect 31297 35031 31355 35037
rect 30558 35000 30564 35012
rect 29932 34972 30564 35000
rect 27488 34963 27517 34969
rect 27488 34960 27494 34963
rect 30558 34960 30564 34972
rect 30616 34960 30622 35012
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22833 34935 22891 34941
rect 22833 34932 22845 34935
rect 22520 34904 22845 34932
rect 22520 34892 22526 34904
rect 22833 34901 22845 34904
rect 22879 34901 22891 34935
rect 22833 34895 22891 34901
rect 27706 34892 27712 34944
rect 27764 34932 27770 34944
rect 30009 34935 30067 34941
rect 30009 34932 30021 34935
rect 27764 34904 30021 34932
rect 27764 34892 27770 34904
rect 30009 34901 30021 34904
rect 30055 34932 30067 34935
rect 31220 34932 31248 35031
rect 31662 35028 31668 35040
rect 31720 35028 31726 35080
rect 31772 35077 31800 35108
rect 32030 35096 32036 35108
rect 32088 35096 32094 35148
rect 32125 35139 32183 35145
rect 32125 35105 32137 35139
rect 32171 35136 32183 35139
rect 32858 35136 32864 35148
rect 32171 35108 32864 35136
rect 32171 35105 32183 35108
rect 32125 35099 32183 35105
rect 32858 35096 32864 35108
rect 32916 35096 32922 35148
rect 31757 35071 31815 35077
rect 31757 35037 31769 35071
rect 31803 35037 31815 35071
rect 31757 35031 31815 35037
rect 31846 35028 31852 35080
rect 31904 35068 31910 35080
rect 31941 35071 31999 35077
rect 31941 35068 31953 35071
rect 31904 35040 31953 35068
rect 31904 35028 31910 35040
rect 31941 35037 31953 35040
rect 31987 35037 31999 35071
rect 32306 35068 32312 35080
rect 32267 35040 32312 35068
rect 31941 35031 31999 35037
rect 32306 35028 32312 35040
rect 32364 35028 32370 35080
rect 48133 35071 48191 35077
rect 48133 35037 48145 35071
rect 48179 35068 48191 35071
rect 48222 35068 48228 35080
rect 48179 35040 48228 35068
rect 48179 35037 48191 35040
rect 48133 35031 48191 35037
rect 48222 35028 48228 35040
rect 48280 35028 48286 35080
rect 30055 34904 31248 34932
rect 30055 34901 30067 34904
rect 30009 34895 30067 34901
rect 47854 34892 47860 34944
rect 47912 34932 47918 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47912 34904 47961 34932
rect 47912 34892 47918 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 20254 34688 20260 34740
rect 20312 34728 20318 34740
rect 20530 34728 20536 34740
rect 20312 34700 20536 34728
rect 20312 34688 20318 34700
rect 20530 34688 20536 34700
rect 20588 34728 20594 34740
rect 20588 34700 24624 34728
rect 20588 34688 20594 34700
rect 19610 34620 19616 34672
rect 19668 34620 19674 34672
rect 23109 34663 23167 34669
rect 23109 34660 23121 34663
rect 22204 34632 23121 34660
rect 22204 34601 22232 34632
rect 23109 34629 23121 34632
rect 23155 34629 23167 34663
rect 23109 34623 23167 34629
rect 24596 34604 24624 34700
rect 26970 34688 26976 34740
rect 27028 34728 27034 34740
rect 28902 34728 28908 34740
rect 27028 34700 28908 34728
rect 27028 34688 27034 34700
rect 28902 34688 28908 34700
rect 28960 34688 28966 34740
rect 29917 34731 29975 34737
rect 29917 34697 29929 34731
rect 29963 34728 29975 34731
rect 30834 34728 30840 34740
rect 29963 34700 30840 34728
rect 29963 34697 29975 34700
rect 29917 34691 29975 34697
rect 30834 34688 30840 34700
rect 30892 34728 30898 34740
rect 31202 34728 31208 34740
rect 30892 34700 31208 34728
rect 30892 34688 30898 34700
rect 31202 34688 31208 34700
rect 31260 34688 31266 34740
rect 26326 34620 26332 34672
rect 26384 34660 26390 34672
rect 28166 34660 28172 34672
rect 26384 34632 28172 34660
rect 26384 34620 26390 34632
rect 28166 34620 28172 34632
rect 28224 34620 28230 34672
rect 30282 34660 30288 34672
rect 28276 34632 30288 34660
rect 22189 34595 22247 34601
rect 22189 34592 22201 34595
rect 22066 34564 22201 34592
rect 18598 34524 18604 34536
rect 18559 34496 18604 34524
rect 18598 34484 18604 34496
rect 18656 34484 18662 34536
rect 20349 34527 20407 34533
rect 20349 34493 20361 34527
rect 20395 34524 20407 34527
rect 21082 34524 21088 34536
rect 20395 34496 21088 34524
rect 20395 34493 20407 34496
rect 20349 34487 20407 34493
rect 21082 34484 21088 34496
rect 21140 34524 21146 34536
rect 22066 34524 22094 34564
rect 22189 34561 22201 34564
rect 22235 34561 22247 34595
rect 22189 34555 22247 34561
rect 22465 34595 22523 34601
rect 22465 34561 22477 34595
rect 22511 34592 22523 34595
rect 22922 34592 22928 34604
rect 22511 34564 22928 34592
rect 22511 34561 22523 34564
rect 22465 34555 22523 34561
rect 22922 34552 22928 34564
rect 22980 34552 22986 34604
rect 24578 34592 24584 34604
rect 24539 34564 24584 34592
rect 24578 34552 24584 34564
rect 24636 34552 24642 34604
rect 27430 34552 27436 34604
rect 27488 34592 27494 34604
rect 27525 34595 27583 34601
rect 27525 34592 27537 34595
rect 27488 34564 27537 34592
rect 27488 34552 27494 34564
rect 27525 34561 27537 34564
rect 27571 34592 27583 34595
rect 28276 34592 28304 34632
rect 30282 34620 30288 34632
rect 30340 34620 30346 34672
rect 30377 34663 30435 34669
rect 30377 34629 30389 34663
rect 30423 34660 30435 34663
rect 30466 34660 30472 34672
rect 30423 34632 30472 34660
rect 30423 34629 30435 34632
rect 30377 34623 30435 34629
rect 30466 34620 30472 34632
rect 30524 34660 30530 34672
rect 30524 34632 30880 34660
rect 30524 34620 30530 34632
rect 30852 34604 30880 34632
rect 27571 34564 28304 34592
rect 28721 34595 28779 34601
rect 27571 34561 27583 34564
rect 27525 34555 27583 34561
rect 28721 34561 28733 34595
rect 28767 34592 28779 34595
rect 28810 34592 28816 34604
rect 28767 34564 28816 34592
rect 28767 34561 28779 34564
rect 28721 34555 28779 34561
rect 28810 34552 28816 34564
rect 28868 34552 28874 34604
rect 29549 34595 29607 34601
rect 29549 34561 29561 34595
rect 29595 34592 29607 34595
rect 30098 34592 30104 34604
rect 29595 34564 30104 34592
rect 29595 34561 29607 34564
rect 29549 34555 29607 34561
rect 21140 34496 22094 34524
rect 22373 34527 22431 34533
rect 21140 34484 21146 34496
rect 22373 34493 22385 34527
rect 22419 34524 22431 34527
rect 22554 34524 22560 34536
rect 22419 34496 22560 34524
rect 22419 34493 22431 34496
rect 22373 34487 22431 34493
rect 22554 34484 22560 34496
rect 22612 34484 22618 34536
rect 24673 34527 24731 34533
rect 24673 34493 24685 34527
rect 24719 34524 24731 34527
rect 25130 34524 25136 34536
rect 24719 34496 25136 34524
rect 24719 34493 24731 34496
rect 24673 34487 24731 34493
rect 25130 34484 25136 34496
rect 25188 34484 25194 34536
rect 27154 34484 27160 34536
rect 27212 34524 27218 34536
rect 27617 34527 27675 34533
rect 27617 34524 27629 34527
rect 27212 34496 27629 34524
rect 27212 34484 27218 34496
rect 27617 34493 27629 34496
rect 27663 34524 27675 34527
rect 27706 34524 27712 34536
rect 27663 34496 27712 34524
rect 27663 34493 27675 34496
rect 27617 34487 27675 34493
rect 27706 34484 27712 34496
rect 27764 34484 27770 34536
rect 27801 34527 27859 34533
rect 27801 34493 27813 34527
rect 27847 34524 27859 34527
rect 27847 34496 27936 34524
rect 27847 34493 27859 34496
rect 27801 34487 27859 34493
rect 27522 34416 27528 34468
rect 27580 34456 27586 34468
rect 27908 34456 27936 34496
rect 28074 34484 28080 34536
rect 28132 34524 28138 34536
rect 29362 34524 29368 34536
rect 28132 34496 29368 34524
rect 28132 34484 28138 34496
rect 29362 34484 29368 34496
rect 29420 34524 29426 34536
rect 29564 34524 29592 34555
rect 30098 34552 30104 34564
rect 30156 34552 30162 34604
rect 30653 34595 30711 34601
rect 30653 34561 30665 34595
rect 30699 34561 30711 34595
rect 30653 34555 30711 34561
rect 29420 34496 29592 34524
rect 29641 34527 29699 34533
rect 29420 34484 29426 34496
rect 29641 34493 29653 34527
rect 29687 34524 29699 34527
rect 30561 34527 30619 34533
rect 30561 34524 30573 34527
rect 29687 34496 30573 34524
rect 29687 34493 29699 34496
rect 29641 34487 29699 34493
rect 30561 34493 30573 34496
rect 30607 34493 30619 34527
rect 30668 34524 30696 34555
rect 30834 34552 30840 34604
rect 30892 34552 30898 34604
rect 47762 34592 47768 34604
rect 47723 34564 47768 34592
rect 47762 34552 47768 34564
rect 47820 34552 47826 34604
rect 31018 34524 31024 34536
rect 30668 34496 31024 34524
rect 30561 34487 30619 34493
rect 28810 34456 28816 34468
rect 27580 34428 27752 34456
rect 27908 34428 28816 34456
rect 27580 34416 27586 34428
rect 18864 34391 18922 34397
rect 18864 34357 18876 34391
rect 18910 34388 18922 34391
rect 20254 34388 20260 34400
rect 18910 34360 20260 34388
rect 18910 34357 18922 34360
rect 18864 34351 18922 34357
rect 20254 34348 20260 34360
rect 20312 34348 20318 34400
rect 22005 34391 22063 34397
rect 22005 34357 22017 34391
rect 22051 34388 22063 34391
rect 22554 34388 22560 34400
rect 22051 34360 22560 34388
rect 22051 34357 22063 34360
rect 22005 34351 22063 34357
rect 22554 34348 22560 34360
rect 22612 34348 22618 34400
rect 23198 34348 23204 34400
rect 23256 34388 23262 34400
rect 27724 34397 27752 34428
rect 28810 34416 28816 34428
rect 28868 34416 28874 34468
rect 30466 34456 30472 34468
rect 29748 34428 30472 34456
rect 29748 34397 29776 34428
rect 30466 34416 30472 34428
rect 30524 34416 30530 34468
rect 30576 34456 30604 34487
rect 31018 34484 31024 34496
rect 31076 34484 31082 34536
rect 30650 34456 30656 34468
rect 30576 34428 30656 34456
rect 30650 34416 30656 34428
rect 30708 34416 30714 34468
rect 23293 34391 23351 34397
rect 23293 34388 23305 34391
rect 23256 34360 23305 34388
rect 23256 34348 23262 34360
rect 23293 34357 23305 34360
rect 23339 34357 23351 34391
rect 23293 34351 23351 34357
rect 27709 34391 27767 34397
rect 27709 34357 27721 34391
rect 27755 34357 27767 34391
rect 27709 34351 27767 34357
rect 29733 34391 29791 34397
rect 29733 34357 29745 34391
rect 29779 34357 29791 34391
rect 30374 34388 30380 34400
rect 30335 34360 30380 34388
rect 29733 34351 29791 34357
rect 30374 34348 30380 34360
rect 30432 34348 30438 34400
rect 30558 34348 30564 34400
rect 30616 34388 30622 34400
rect 30837 34391 30895 34397
rect 30837 34388 30849 34391
rect 30616 34360 30849 34388
rect 30616 34348 30622 34360
rect 30837 34357 30849 34360
rect 30883 34357 30895 34391
rect 30837 34351 30895 34357
rect 47210 34348 47216 34400
rect 47268 34388 47274 34400
rect 47581 34391 47639 34397
rect 47581 34388 47593 34391
rect 47268 34360 47593 34388
rect 47268 34348 47274 34360
rect 47581 34357 47593 34360
rect 47627 34357 47639 34391
rect 47581 34351 47639 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 19610 34184 19616 34196
rect 19571 34156 19616 34184
rect 19610 34144 19616 34156
rect 19668 34144 19674 34196
rect 20254 34144 20260 34196
rect 20312 34184 20318 34196
rect 21545 34187 21603 34193
rect 21545 34184 21557 34187
rect 20312 34156 21557 34184
rect 20312 34144 20318 34156
rect 21545 34153 21557 34156
rect 21591 34153 21603 34187
rect 21545 34147 21603 34153
rect 22094 34144 22100 34196
rect 22152 34184 22158 34196
rect 22373 34187 22431 34193
rect 22373 34184 22385 34187
rect 22152 34156 22385 34184
rect 22152 34144 22158 34156
rect 22373 34153 22385 34156
rect 22419 34184 22431 34187
rect 23842 34184 23848 34196
rect 22419 34156 23848 34184
rect 22419 34153 22431 34156
rect 22373 34147 22431 34153
rect 23842 34144 23848 34156
rect 23900 34144 23906 34196
rect 25222 34144 25228 34196
rect 25280 34184 25286 34196
rect 28721 34187 28779 34193
rect 28721 34184 28733 34187
rect 25280 34156 28733 34184
rect 25280 34144 25286 34156
rect 28721 34153 28733 34156
rect 28767 34184 28779 34187
rect 28810 34184 28816 34196
rect 28767 34156 28816 34184
rect 28767 34153 28779 34156
rect 28721 34147 28779 34153
rect 28810 34144 28816 34156
rect 28868 34144 28874 34196
rect 30098 34144 30104 34196
rect 30156 34184 30162 34196
rect 31297 34187 31355 34193
rect 31297 34184 31309 34187
rect 30156 34156 31309 34184
rect 30156 34144 30162 34156
rect 31297 34153 31309 34156
rect 31343 34153 31355 34187
rect 31297 34147 31355 34153
rect 30650 34076 30656 34128
rect 30708 34116 30714 34128
rect 30708 34088 31524 34116
rect 30708 34076 30714 34088
rect 1946 34008 1952 34060
rect 2004 34048 2010 34060
rect 21177 34051 21235 34057
rect 21177 34048 21189 34051
rect 2004 34020 21189 34048
rect 2004 34008 2010 34020
rect 21177 34017 21189 34020
rect 21223 34017 21235 34051
rect 21177 34011 21235 34017
rect 21376 34020 22140 34048
rect 19521 33983 19579 33989
rect 19521 33949 19533 33983
rect 19567 33980 19579 33983
rect 20530 33980 20536 33992
rect 19567 33952 20536 33980
rect 19567 33949 19579 33952
rect 19521 33943 19579 33949
rect 20530 33940 20536 33952
rect 20588 33940 20594 33992
rect 20809 33983 20867 33989
rect 20809 33949 20821 33983
rect 20855 33949 20867 33983
rect 20990 33980 20996 33992
rect 20951 33952 20996 33980
rect 20809 33943 20867 33949
rect 20824 33912 20852 33943
rect 20990 33940 20996 33952
rect 21048 33940 21054 33992
rect 21082 33940 21088 33992
rect 21140 33980 21146 33992
rect 21376 33989 21404 34020
rect 21361 33983 21419 33989
rect 21140 33952 21185 33980
rect 21140 33940 21146 33952
rect 21361 33949 21373 33983
rect 21407 33949 21419 33983
rect 22002 33980 22008 33992
rect 21963 33952 22008 33980
rect 21361 33943 21419 33949
rect 22002 33940 22008 33952
rect 22060 33940 22066 33992
rect 22112 33980 22140 34020
rect 22186 34008 22192 34060
rect 22244 34048 22250 34060
rect 23290 34048 23296 34060
rect 22244 34020 23296 34048
rect 22244 34008 22250 34020
rect 23290 34008 23296 34020
rect 23348 34048 23354 34060
rect 24397 34051 24455 34057
rect 24397 34048 24409 34051
rect 23348 34020 24409 34048
rect 23348 34008 23354 34020
rect 24397 34017 24409 34020
rect 24443 34017 24455 34051
rect 28626 34048 28632 34060
rect 24397 34011 24455 34017
rect 27264 34020 28632 34048
rect 22373 33983 22431 33989
rect 22112 33952 22232 33980
rect 22204 33912 22232 33952
rect 22373 33949 22385 33983
rect 22419 33980 22431 33983
rect 22554 33980 22560 33992
rect 22419 33952 22560 33980
rect 22419 33949 22431 33952
rect 22373 33943 22431 33949
rect 22554 33940 22560 33952
rect 22612 33940 22618 33992
rect 22738 33940 22744 33992
rect 22796 33980 22802 33992
rect 23014 33980 23020 33992
rect 22796 33952 23020 33980
rect 22796 33940 22802 33952
rect 23014 33940 23020 33952
rect 23072 33940 23078 33992
rect 27264 33924 27292 34020
rect 28626 34008 28632 34020
rect 28684 34008 28690 34060
rect 29917 34051 29975 34057
rect 29917 34017 29929 34051
rect 29963 34048 29975 34051
rect 31386 34048 31392 34060
rect 29963 34020 31392 34048
rect 29963 34017 29975 34020
rect 29917 34011 29975 34017
rect 31386 34008 31392 34020
rect 31444 34008 31450 34060
rect 31496 34057 31524 34088
rect 31481 34051 31539 34057
rect 31481 34017 31493 34051
rect 31527 34017 31539 34051
rect 47118 34048 47124 34060
rect 47079 34020 47124 34048
rect 31481 34011 31539 34017
rect 47118 34008 47124 34020
rect 47176 34008 47182 34060
rect 47670 34048 47676 34060
rect 47631 34020 47676 34048
rect 47670 34008 47676 34020
rect 47728 34008 47734 34060
rect 29546 33940 29552 33992
rect 29604 33980 29610 33992
rect 29733 33983 29791 33989
rect 29733 33980 29745 33983
rect 29604 33952 29745 33980
rect 29604 33940 29610 33952
rect 29733 33949 29745 33952
rect 29779 33949 29791 33983
rect 30006 33980 30012 33992
rect 29967 33952 30012 33980
rect 29733 33943 29791 33949
rect 30006 33940 30012 33952
rect 30064 33940 30070 33992
rect 30469 33983 30527 33989
rect 30469 33949 30481 33983
rect 30515 33949 30527 33983
rect 30469 33943 30527 33949
rect 24670 33912 24676 33924
rect 20824 33884 22094 33912
rect 22204 33884 23244 33912
rect 24631 33884 24676 33912
rect 22066 33844 22094 33884
rect 23216 33853 23244 33884
rect 24670 33872 24676 33884
rect 24728 33872 24734 33924
rect 25130 33872 25136 33924
rect 25188 33872 25194 33924
rect 27246 33912 27252 33924
rect 27207 33884 27252 33912
rect 27246 33872 27252 33884
rect 27304 33872 27310 33924
rect 28258 33872 28264 33924
rect 28316 33912 28322 33924
rect 28629 33915 28687 33921
rect 28629 33912 28641 33915
rect 28316 33884 28641 33912
rect 28316 33872 28322 33884
rect 28629 33881 28641 33884
rect 28675 33912 28687 33915
rect 28902 33912 28908 33924
rect 28675 33884 28908 33912
rect 28675 33881 28687 33884
rect 28629 33875 28687 33881
rect 28902 33872 28908 33884
rect 28960 33912 28966 33924
rect 30484 33912 30512 33943
rect 30834 33940 30840 33992
rect 30892 33980 30898 33992
rect 31205 33983 31263 33989
rect 31205 33980 31217 33983
rect 30892 33952 31217 33980
rect 30892 33940 30898 33952
rect 31205 33949 31217 33952
rect 31251 33949 31263 33983
rect 31205 33943 31263 33949
rect 28960 33884 30512 33912
rect 28960 33872 28966 33884
rect 47210 33872 47216 33924
rect 47268 33912 47274 33924
rect 47268 33884 47313 33912
rect 47268 33872 47274 33884
rect 22557 33847 22615 33853
rect 22557 33844 22569 33847
rect 22066 33816 22569 33844
rect 22557 33813 22569 33816
rect 22603 33813 22615 33847
rect 22557 33807 22615 33813
rect 23201 33847 23259 33853
rect 23201 33813 23213 33847
rect 23247 33844 23259 33847
rect 23566 33844 23572 33856
rect 23247 33816 23572 33844
rect 23247 33813 23259 33816
rect 23201 33807 23259 33813
rect 23566 33804 23572 33816
rect 23624 33804 23630 33856
rect 25314 33804 25320 33856
rect 25372 33844 25378 33856
rect 26145 33847 26203 33853
rect 26145 33844 26157 33847
rect 25372 33816 26157 33844
rect 25372 33804 25378 33816
rect 26145 33813 26157 33816
rect 26191 33813 26203 33847
rect 27338 33844 27344 33856
rect 27251 33816 27344 33844
rect 26145 33807 26203 33813
rect 27338 33804 27344 33816
rect 27396 33844 27402 33856
rect 28718 33844 28724 33856
rect 27396 33816 28724 33844
rect 27396 33804 27402 33816
rect 28718 33804 28724 33816
rect 28776 33804 28782 33856
rect 29270 33804 29276 33856
rect 29328 33844 29334 33856
rect 29549 33847 29607 33853
rect 29549 33844 29561 33847
rect 29328 33816 29561 33844
rect 29328 33804 29334 33816
rect 29549 33813 29561 33816
rect 29595 33813 29607 33847
rect 29549 33807 29607 33813
rect 30558 33804 30564 33856
rect 30616 33844 30622 33856
rect 30653 33847 30711 33853
rect 30653 33844 30665 33847
rect 30616 33816 30665 33844
rect 30616 33804 30622 33816
rect 30653 33813 30665 33816
rect 30699 33813 30711 33847
rect 30653 33807 30711 33813
rect 31294 33804 31300 33856
rect 31352 33844 31358 33856
rect 31481 33847 31539 33853
rect 31481 33844 31493 33847
rect 31352 33816 31493 33844
rect 31352 33804 31358 33816
rect 31481 33813 31493 33816
rect 31527 33813 31539 33847
rect 31481 33807 31539 33813
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 23290 33640 23296 33652
rect 23251 33612 23296 33640
rect 23290 33600 23296 33612
rect 23348 33600 23354 33652
rect 47762 33600 47768 33652
rect 47820 33640 47826 33652
rect 48041 33643 48099 33649
rect 48041 33640 48053 33643
rect 47820 33612 48053 33640
rect 47820 33600 47826 33612
rect 48041 33609 48053 33612
rect 48087 33609 48099 33643
rect 48041 33603 48099 33609
rect 23201 33575 23259 33581
rect 23201 33541 23213 33575
rect 23247 33572 23259 33575
rect 25038 33572 25044 33584
rect 23247 33544 25044 33572
rect 23247 33541 23259 33544
rect 23201 33535 23259 33541
rect 25038 33532 25044 33544
rect 25096 33532 25102 33584
rect 29270 33572 29276 33584
rect 29231 33544 29276 33572
rect 29270 33532 29276 33544
rect 29328 33532 29334 33584
rect 1578 33504 1584 33516
rect 1539 33476 1584 33504
rect 1578 33464 1584 33476
rect 1636 33464 1642 33516
rect 2222 33504 2228 33516
rect 2183 33476 2228 33504
rect 2222 33464 2228 33476
rect 2280 33464 2286 33516
rect 19797 33507 19855 33513
rect 19797 33473 19809 33507
rect 19843 33504 19855 33507
rect 20530 33504 20536 33516
rect 19843 33476 20536 33504
rect 19843 33473 19855 33476
rect 19797 33467 19855 33473
rect 20530 33464 20536 33476
rect 20588 33464 20594 33516
rect 22002 33504 22008 33516
rect 21963 33476 22008 33504
rect 22002 33464 22008 33476
rect 22060 33464 22066 33516
rect 24118 33513 24124 33516
rect 24107 33507 24124 33513
rect 24107 33473 24119 33507
rect 24176 33504 24182 33516
rect 25222 33504 25228 33516
rect 24176 33476 24716 33504
rect 25183 33476 25228 33504
rect 24107 33467 24124 33473
rect 24118 33464 24124 33467
rect 24176 33464 24182 33476
rect 2409 33439 2467 33445
rect 2409 33405 2421 33439
rect 2455 33436 2467 33439
rect 3786 33436 3792 33448
rect 2455 33408 3792 33436
rect 2455 33405 2467 33408
rect 2409 33399 2467 33405
rect 3786 33396 3792 33408
rect 3844 33396 3850 33448
rect 4065 33439 4123 33445
rect 4065 33405 4077 33439
rect 4111 33436 4123 33439
rect 4614 33436 4620 33448
rect 4111 33408 4620 33436
rect 4111 33405 4123 33408
rect 4065 33399 4123 33405
rect 4614 33396 4620 33408
rect 4672 33396 4678 33448
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 23658 33436 23664 33448
rect 22327 33408 23664 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 23658 33396 23664 33408
rect 23716 33396 23722 33448
rect 23934 33436 23940 33448
rect 23895 33408 23940 33436
rect 23934 33396 23940 33408
rect 23992 33396 23998 33448
rect 24688 33436 24716 33476
rect 25222 33464 25228 33476
rect 25280 33464 25286 33516
rect 25314 33464 25320 33516
rect 25372 33504 25378 33516
rect 25593 33507 25651 33513
rect 25372 33476 25417 33504
rect 25372 33464 25378 33476
rect 25593 33473 25605 33507
rect 25639 33504 25651 33507
rect 27338 33504 27344 33516
rect 25639 33476 27344 33504
rect 25639 33473 25651 33476
rect 25593 33467 25651 33473
rect 25332 33436 25360 33464
rect 24688 33408 25360 33436
rect 24394 33368 24400 33380
rect 24355 33340 24400 33368
rect 24394 33328 24400 33340
rect 24452 33328 24458 33380
rect 24486 33328 24492 33380
rect 24544 33368 24550 33380
rect 25608 33368 25636 33467
rect 27338 33464 27344 33476
rect 27396 33464 27402 33516
rect 30374 33464 30380 33516
rect 30432 33464 30438 33516
rect 46842 33504 46848 33516
rect 46803 33476 46848 33504
rect 46842 33464 46848 33476
rect 46900 33464 46906 33516
rect 47302 33464 47308 33516
rect 47360 33504 47366 33516
rect 47581 33507 47639 33513
rect 47581 33504 47593 33507
rect 47360 33476 47593 33504
rect 47360 33464 47366 33476
rect 47581 33473 47593 33476
rect 47627 33473 47639 33507
rect 47581 33467 47639 33473
rect 28994 33436 29000 33448
rect 28955 33408 29000 33436
rect 28994 33396 29000 33408
rect 29052 33396 29058 33448
rect 29270 33396 29276 33448
rect 29328 33436 29334 33448
rect 30006 33436 30012 33448
rect 29328 33408 30012 33436
rect 29328 33396 29334 33408
rect 30006 33396 30012 33408
rect 30064 33396 30070 33448
rect 44174 33368 44180 33380
rect 24544 33340 25636 33368
rect 30300 33340 44180 33368
rect 24544 33328 24550 33340
rect 1397 33303 1455 33309
rect 1397 33269 1409 33303
rect 1443 33300 1455 33303
rect 2774 33300 2780 33312
rect 1443 33272 2780 33300
rect 1443 33269 1455 33272
rect 1397 33263 1455 33269
rect 2774 33260 2780 33272
rect 2832 33260 2838 33312
rect 19889 33303 19947 33309
rect 19889 33269 19901 33303
rect 19935 33300 19947 33303
rect 19978 33300 19984 33312
rect 19935 33272 19984 33300
rect 19935 33269 19947 33272
rect 19889 33263 19947 33269
rect 19978 33260 19984 33272
rect 20036 33260 20042 33312
rect 21818 33300 21824 33312
rect 21779 33272 21824 33300
rect 21818 33260 21824 33272
rect 21876 33260 21882 33312
rect 22186 33300 22192 33312
rect 22147 33272 22192 33300
rect 22186 33260 22192 33272
rect 22244 33260 22250 33312
rect 22554 33260 22560 33312
rect 22612 33300 22618 33312
rect 24504 33300 24532 33328
rect 22612 33272 24532 33300
rect 22612 33260 22618 33272
rect 24946 33260 24952 33312
rect 25004 33300 25010 33312
rect 25041 33303 25099 33309
rect 25041 33300 25053 33303
rect 25004 33272 25053 33300
rect 25004 33260 25010 33272
rect 25041 33269 25053 33272
rect 25087 33269 25099 33303
rect 25041 33263 25099 33269
rect 25501 33303 25559 33309
rect 25501 33269 25513 33303
rect 25547 33300 25559 33303
rect 30300 33300 30328 33340
rect 44174 33328 44180 33340
rect 44232 33328 44238 33380
rect 25547 33272 30328 33300
rect 25547 33269 25559 33272
rect 25501 33263 25559 33269
rect 30650 33260 30656 33312
rect 30708 33300 30714 33312
rect 30745 33303 30803 33309
rect 30745 33300 30757 33303
rect 30708 33272 30757 33300
rect 30708 33260 30714 33272
rect 30745 33269 30757 33272
rect 30791 33269 30803 33303
rect 46934 33300 46940 33312
rect 46895 33272 46940 33300
rect 30745 33263 30803 33269
rect 46934 33260 46940 33272
rect 46992 33260 46998 33312
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 2774 33096 2780 33108
rect 2735 33068 2780 33096
rect 2774 33056 2780 33068
rect 2832 33056 2838 33108
rect 3786 33096 3792 33108
rect 3747 33068 3792 33096
rect 3786 33056 3792 33068
rect 3844 33056 3850 33108
rect 21913 33099 21971 33105
rect 21913 33065 21925 33099
rect 21959 33096 21971 33099
rect 22002 33096 22008 33108
rect 21959 33068 22008 33096
rect 21959 33065 21971 33068
rect 21913 33059 21971 33065
rect 22002 33056 22008 33068
rect 22060 33056 22066 33108
rect 22186 33056 22192 33108
rect 22244 33096 22250 33108
rect 23017 33099 23075 33105
rect 23017 33096 23029 33099
rect 22244 33068 23029 33096
rect 22244 33056 22250 33068
rect 23017 33065 23029 33068
rect 23063 33065 23075 33099
rect 23017 33059 23075 33065
rect 24394 33056 24400 33108
rect 24452 33096 24458 33108
rect 24765 33099 24823 33105
rect 24765 33096 24777 33099
rect 24452 33068 24777 33096
rect 24452 33056 24458 33068
rect 24765 33065 24777 33068
rect 24811 33065 24823 33099
rect 24765 33059 24823 33065
rect 27982 33056 27988 33108
rect 28040 33096 28046 33108
rect 28261 33099 28319 33105
rect 28261 33096 28273 33099
rect 28040 33068 28273 33096
rect 28040 33056 28046 33068
rect 28261 33065 28273 33068
rect 28307 33096 28319 33099
rect 28350 33096 28356 33108
rect 28307 33068 28356 33096
rect 28307 33065 28319 33068
rect 28261 33059 28319 33065
rect 28350 33056 28356 33068
rect 28408 33056 28414 33108
rect 28994 33056 29000 33108
rect 29052 33096 29058 33108
rect 30745 33099 30803 33105
rect 30745 33096 30757 33099
rect 29052 33068 30757 33096
rect 29052 33056 29058 33068
rect 30745 33065 30757 33068
rect 30791 33096 30803 33099
rect 32122 33096 32128 33108
rect 30791 33068 32128 33096
rect 30791 33065 30803 33068
rect 30745 33059 30803 33065
rect 32122 33056 32128 33068
rect 32180 33056 32186 33108
rect 46198 33096 46204 33108
rect 41386 33068 46204 33096
rect 25222 33028 25228 33040
rect 22112 33000 25228 33028
rect 1394 32960 1400 32972
rect 1355 32932 1400 32960
rect 1394 32920 1400 32932
rect 1452 32920 1458 32972
rect 3145 32963 3203 32969
rect 3145 32929 3157 32963
rect 3191 32960 3203 32963
rect 19521 32963 19579 32969
rect 3191 32932 4016 32960
rect 3191 32929 3203 32932
rect 3145 32923 3203 32929
rect 1673 32895 1731 32901
rect 1673 32861 1685 32895
rect 1719 32892 1731 32895
rect 2682 32892 2688 32904
rect 1719 32864 2688 32892
rect 1719 32861 1731 32864
rect 1673 32855 1731 32861
rect 2682 32852 2688 32864
rect 2740 32852 2746 32904
rect 3988 32901 4016 32932
rect 19521 32929 19533 32963
rect 19567 32960 19579 32963
rect 21818 32960 21824 32972
rect 19567 32932 21824 32960
rect 19567 32929 19579 32932
rect 19521 32923 19579 32929
rect 21818 32920 21824 32932
rect 21876 32920 21882 32972
rect 3973 32895 4031 32901
rect 3973 32861 3985 32895
rect 4019 32861 4031 32895
rect 3973 32855 4031 32861
rect 18138 32852 18144 32904
rect 18196 32892 18202 32904
rect 18598 32892 18604 32904
rect 18196 32864 18604 32892
rect 18196 32852 18202 32864
rect 18598 32852 18604 32864
rect 18656 32892 18662 32904
rect 22112 32901 22140 33000
rect 25222 32988 25228 33000
rect 25280 32988 25286 33040
rect 29270 33028 29276 33040
rect 26206 33000 29276 33028
rect 22278 32920 22284 32972
rect 22336 32960 22342 32972
rect 22373 32963 22431 32969
rect 22373 32960 22385 32963
rect 22336 32932 22385 32960
rect 22336 32920 22342 32932
rect 22373 32929 22385 32932
rect 22419 32929 22431 32963
rect 22373 32923 22431 32929
rect 24397 32963 24455 32969
rect 24397 32929 24409 32963
rect 24443 32960 24455 32963
rect 24670 32960 24676 32972
rect 24443 32932 24676 32960
rect 24443 32929 24455 32932
rect 24397 32923 24455 32929
rect 24670 32920 24676 32932
rect 24728 32920 24734 32972
rect 24946 32960 24952 32972
rect 24780 32932 24952 32960
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18656 32864 19257 32892
rect 18656 32852 18662 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 22097 32895 22155 32901
rect 22097 32861 22109 32895
rect 22143 32861 22155 32895
rect 22097 32855 22155 32861
rect 22189 32895 22247 32901
rect 22189 32861 22201 32895
rect 22235 32861 22247 32895
rect 22189 32855 22247 32861
rect 22465 32895 22523 32901
rect 22465 32861 22477 32895
rect 22511 32892 22523 32895
rect 22554 32892 22560 32904
rect 22511 32864 22560 32892
rect 22511 32861 22523 32864
rect 22465 32855 22523 32861
rect 19978 32784 19984 32836
rect 20036 32784 20042 32836
rect 22204 32824 22232 32855
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 22922 32892 22928 32904
rect 22883 32864 22928 32892
rect 22922 32852 22928 32864
rect 22980 32852 22986 32904
rect 23109 32895 23167 32901
rect 23109 32861 23121 32895
rect 23155 32892 23167 32895
rect 23934 32892 23940 32904
rect 23155 32864 23940 32892
rect 23155 32861 23167 32864
rect 23109 32855 23167 32861
rect 23934 32852 23940 32864
rect 23992 32852 23998 32904
rect 24581 32895 24639 32901
rect 24581 32861 24593 32895
rect 24627 32892 24639 32895
rect 24780 32892 24808 32932
rect 24946 32920 24952 32932
rect 25004 32920 25010 32972
rect 24627 32864 24808 32892
rect 24857 32895 24915 32901
rect 24627 32861 24639 32864
rect 24581 32855 24639 32861
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 26206 32892 26234 33000
rect 29270 32988 29276 33000
rect 29328 32988 29334 33040
rect 29546 33028 29552 33040
rect 29507 33000 29552 33028
rect 29546 32988 29552 33000
rect 29604 32988 29610 33040
rect 30650 33028 30656 33040
rect 29840 33000 30656 33028
rect 27246 32920 27252 32972
rect 27304 32960 27310 32972
rect 27525 32963 27583 32969
rect 27525 32960 27537 32963
rect 27304 32932 27537 32960
rect 27304 32920 27310 32932
rect 27525 32929 27537 32932
rect 27571 32929 27583 32963
rect 27525 32923 27583 32929
rect 28166 32892 28172 32904
rect 24903 32864 26234 32892
rect 28079 32864 28172 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 21284 32796 22232 32824
rect 21284 32768 21312 32796
rect 23658 32784 23664 32836
rect 23716 32824 23722 32836
rect 24872 32824 24900 32855
rect 28166 32852 28172 32864
rect 28224 32892 28230 32904
rect 28224 32864 28672 32892
rect 28224 32852 28230 32864
rect 23716 32796 24900 32824
rect 26697 32827 26755 32833
rect 23716 32784 23722 32796
rect 26697 32793 26709 32827
rect 26743 32824 26755 32827
rect 27341 32827 27399 32833
rect 27341 32824 27353 32827
rect 26743 32796 27353 32824
rect 26743 32793 26755 32796
rect 26697 32787 26755 32793
rect 27341 32793 27353 32796
rect 27387 32824 27399 32827
rect 27982 32824 27988 32836
rect 27387 32796 27988 32824
rect 27387 32793 27399 32796
rect 27341 32787 27399 32793
rect 27982 32784 27988 32796
rect 28040 32784 28046 32836
rect 19426 32716 19432 32768
rect 19484 32756 19490 32768
rect 20254 32756 20260 32768
rect 19484 32728 20260 32756
rect 19484 32716 19490 32728
rect 20254 32716 20260 32728
rect 20312 32716 20318 32768
rect 20993 32759 21051 32765
rect 20993 32725 21005 32759
rect 21039 32756 21051 32759
rect 21266 32756 21272 32768
rect 21039 32728 21272 32756
rect 21039 32725 21051 32728
rect 20993 32719 21051 32725
rect 21266 32716 21272 32728
rect 21324 32716 21330 32768
rect 26973 32759 27031 32765
rect 26973 32725 26985 32759
rect 27019 32756 27031 32759
rect 27154 32756 27160 32768
rect 27019 32728 27160 32756
rect 27019 32725 27031 32728
rect 26973 32719 27031 32725
rect 27154 32716 27160 32728
rect 27212 32716 27218 32768
rect 27430 32716 27436 32768
rect 27488 32756 27494 32768
rect 28644 32756 28672 32864
rect 28810 32852 28816 32904
rect 28868 32892 28874 32904
rect 29840 32901 29868 33000
rect 30650 32988 30656 33000
rect 30708 32988 30714 33040
rect 31386 33028 31392 33040
rect 31347 33000 31392 33028
rect 31386 32988 31392 33000
rect 31444 32988 31450 33040
rect 32030 32988 32036 33040
rect 32088 33028 32094 33040
rect 41386 33028 41414 33068
rect 46198 33056 46204 33068
rect 46256 33096 46262 33108
rect 46474 33096 46480 33108
rect 46256 33068 46480 33096
rect 46256 33056 46262 33068
rect 46474 33056 46480 33068
rect 46532 33056 46538 33108
rect 32088 33000 41414 33028
rect 32088 32988 32094 33000
rect 30009 32963 30067 32969
rect 30009 32929 30021 32963
rect 30055 32960 30067 32963
rect 47581 32963 47639 32969
rect 47581 32960 47593 32963
rect 30055 32932 47593 32960
rect 30055 32929 30067 32932
rect 30009 32923 30067 32929
rect 47581 32929 47593 32932
rect 47627 32929 47639 32963
rect 47581 32923 47639 32929
rect 29733 32895 29791 32901
rect 29733 32892 29745 32895
rect 28868 32864 29745 32892
rect 28868 32852 28874 32864
rect 29733 32861 29745 32864
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 29825 32895 29883 32901
rect 29825 32861 29837 32895
rect 29871 32861 29883 32895
rect 29825 32855 29883 32861
rect 30101 32895 30159 32901
rect 30101 32861 30113 32895
rect 30147 32861 30159 32895
rect 31294 32892 31300 32904
rect 31255 32864 31300 32892
rect 30101 32855 30159 32861
rect 28718 32784 28724 32836
rect 28776 32824 28782 32836
rect 30116 32824 30144 32855
rect 31294 32852 31300 32864
rect 31352 32852 31358 32904
rect 31386 32852 31392 32904
rect 31444 32892 31450 32904
rect 31481 32895 31539 32901
rect 31481 32892 31493 32895
rect 31444 32864 31493 32892
rect 31444 32852 31450 32864
rect 31481 32861 31493 32864
rect 31527 32861 31539 32895
rect 31481 32855 31539 32861
rect 31570 32852 31576 32904
rect 31628 32892 31634 32904
rect 32309 32895 32367 32901
rect 32309 32892 32321 32895
rect 31628 32864 32321 32892
rect 31628 32852 31634 32864
rect 32309 32861 32321 32864
rect 32355 32861 32367 32895
rect 32582 32892 32588 32904
rect 32543 32864 32588 32892
rect 32309 32855 32367 32861
rect 32582 32852 32588 32864
rect 32640 32852 32646 32904
rect 46290 32852 46296 32904
rect 46348 32892 46354 32904
rect 46845 32895 46903 32901
rect 46845 32892 46857 32895
rect 46348 32864 46857 32892
rect 46348 32852 46354 32864
rect 46845 32861 46857 32864
rect 46891 32861 46903 32895
rect 46845 32855 46903 32861
rect 47305 32895 47363 32901
rect 47305 32861 47317 32895
rect 47351 32861 47363 32895
rect 47305 32855 47363 32861
rect 30650 32824 30656 32836
rect 28776 32796 30144 32824
rect 30611 32796 30656 32824
rect 28776 32784 28782 32796
rect 30650 32784 30656 32796
rect 30708 32784 30714 32836
rect 30742 32784 30748 32836
rect 30800 32824 30806 32836
rect 32030 32824 32036 32836
rect 30800 32796 32036 32824
rect 30800 32784 30806 32796
rect 32030 32784 32036 32796
rect 32088 32784 32094 32836
rect 32125 32827 32183 32833
rect 32125 32793 32137 32827
rect 32171 32824 32183 32827
rect 32398 32824 32404 32836
rect 32171 32796 32404 32824
rect 32171 32793 32183 32796
rect 32125 32787 32183 32793
rect 32398 32784 32404 32796
rect 32456 32784 32462 32836
rect 47320 32824 47348 32855
rect 46860 32796 47348 32824
rect 46860 32768 46888 32796
rect 31018 32756 31024 32768
rect 27488 32728 27533 32756
rect 28644 32728 31024 32756
rect 27488 32716 27494 32728
rect 31018 32716 31024 32728
rect 31076 32716 31082 32768
rect 32490 32756 32496 32768
rect 32451 32728 32496 32756
rect 32490 32716 32496 32728
rect 32548 32716 32554 32768
rect 46842 32716 46848 32768
rect 46900 32716 46906 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 19978 32512 19984 32564
rect 20036 32552 20042 32564
rect 20530 32552 20536 32564
rect 20036 32524 20536 32552
rect 20036 32512 20042 32524
rect 20530 32512 20536 32524
rect 20588 32512 20594 32564
rect 21269 32555 21327 32561
rect 21269 32521 21281 32555
rect 21315 32552 21327 32555
rect 22922 32552 22928 32564
rect 21315 32524 22928 32552
rect 21315 32521 21327 32524
rect 21269 32515 21327 32521
rect 22922 32512 22928 32524
rect 22980 32512 22986 32564
rect 23474 32512 23480 32564
rect 23532 32552 23538 32564
rect 23569 32555 23627 32561
rect 23569 32552 23581 32555
rect 23532 32524 23581 32552
rect 23532 32512 23538 32524
rect 23569 32521 23581 32524
rect 23615 32521 23627 32555
rect 25038 32552 25044 32564
rect 24999 32524 25044 32552
rect 23569 32515 23627 32521
rect 25038 32512 25044 32524
rect 25096 32512 25102 32564
rect 30101 32555 30159 32561
rect 30101 32521 30113 32555
rect 30147 32552 30159 32555
rect 30374 32552 30380 32564
rect 30147 32524 30380 32552
rect 30147 32521 30159 32524
rect 30101 32515 30159 32521
rect 30374 32512 30380 32524
rect 30432 32512 30438 32564
rect 30466 32512 30472 32564
rect 30524 32552 30530 32564
rect 30524 32524 30972 32552
rect 30524 32512 30530 32524
rect 30944 32496 30972 32524
rect 31018 32512 31024 32564
rect 31076 32552 31082 32564
rect 31570 32552 31576 32564
rect 31076 32524 31432 32552
rect 31531 32524 31576 32552
rect 31076 32512 31082 32524
rect 19426 32444 19432 32496
rect 19484 32444 19490 32496
rect 20254 32444 20260 32496
rect 20312 32484 20318 32496
rect 30742 32484 30748 32496
rect 20312 32456 30748 32484
rect 20312 32444 20318 32456
rect 30742 32444 30748 32456
rect 30800 32444 30806 32496
rect 30926 32444 30932 32496
rect 30984 32484 30990 32496
rect 31297 32487 31355 32493
rect 31297 32484 31309 32487
rect 30984 32456 31309 32484
rect 30984 32444 30990 32456
rect 31297 32453 31309 32456
rect 31343 32453 31355 32487
rect 31404 32484 31432 32524
rect 31570 32512 31576 32524
rect 31628 32512 31634 32564
rect 46934 32552 46940 32564
rect 31726 32524 46940 32552
rect 31726 32484 31754 32524
rect 46934 32512 46940 32524
rect 46992 32512 46998 32564
rect 32398 32484 32404 32496
rect 31404 32456 31754 32484
rect 32359 32456 32404 32484
rect 31297 32447 31355 32453
rect 32398 32444 32404 32456
rect 32456 32444 32462 32496
rect 33410 32444 33416 32496
rect 33468 32444 33474 32496
rect 18138 32416 18144 32428
rect 18099 32388 18144 32416
rect 18138 32376 18144 32388
rect 18196 32376 18202 32428
rect 20993 32419 21051 32425
rect 20993 32385 21005 32419
rect 21039 32416 21051 32419
rect 21910 32416 21916 32428
rect 21039 32388 21916 32416
rect 21039 32385 21051 32388
rect 20993 32379 21051 32385
rect 21910 32376 21916 32388
rect 21968 32416 21974 32428
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 21968 32388 22109 32416
rect 21968 32376 21974 32388
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 23109 32419 23167 32425
rect 23109 32385 23121 32419
rect 23155 32416 23167 32419
rect 23155 32388 23336 32416
rect 23155 32385 23167 32388
rect 23109 32379 23167 32385
rect 1670 32308 1676 32360
rect 1728 32348 1734 32360
rect 1765 32351 1823 32357
rect 1765 32348 1777 32351
rect 1728 32320 1777 32348
rect 1728 32308 1734 32320
rect 1765 32317 1777 32320
rect 1811 32317 1823 32351
rect 1765 32311 1823 32317
rect 1949 32351 2007 32357
rect 1949 32317 1961 32351
rect 1995 32348 2007 32351
rect 2222 32348 2228 32360
rect 1995 32320 2228 32348
rect 1995 32317 2007 32320
rect 1949 32311 2007 32317
rect 2222 32308 2228 32320
rect 2280 32308 2286 32360
rect 2774 32348 2780 32360
rect 2735 32320 2780 32348
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 18417 32351 18475 32357
rect 18417 32317 18429 32351
rect 18463 32348 18475 32351
rect 20530 32348 20536 32360
rect 18463 32320 20536 32348
rect 18463 32317 18475 32320
rect 18417 32311 18475 32317
rect 20530 32308 20536 32320
rect 20588 32308 20594 32360
rect 21266 32348 21272 32360
rect 21227 32320 21272 32348
rect 21266 32308 21272 32320
rect 21324 32308 21330 32360
rect 21821 32351 21879 32357
rect 21821 32317 21833 32351
rect 21867 32317 21879 32351
rect 23198 32348 23204 32360
rect 23111 32320 23204 32348
rect 21821 32311 21879 32317
rect 19889 32283 19947 32289
rect 19889 32249 19901 32283
rect 19935 32280 19947 32283
rect 21836 32280 21864 32311
rect 23198 32308 23204 32320
rect 23256 32308 23262 32360
rect 23308 32348 23336 32388
rect 23382 32376 23388 32428
rect 23440 32416 23446 32428
rect 24029 32419 24087 32425
rect 23440 32388 23485 32416
rect 23440 32376 23446 32388
rect 24029 32385 24041 32419
rect 24075 32416 24087 32419
rect 24118 32416 24124 32428
rect 24075 32388 24124 32416
rect 24075 32385 24087 32388
rect 24029 32379 24087 32385
rect 24118 32376 24124 32388
rect 24176 32376 24182 32428
rect 24213 32419 24271 32425
rect 24213 32385 24225 32419
rect 24259 32416 24271 32419
rect 24854 32416 24860 32428
rect 24259 32388 24860 32416
rect 24259 32385 24271 32388
rect 24213 32379 24271 32385
rect 24854 32376 24860 32388
rect 24912 32376 24918 32428
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32416 25007 32419
rect 27062 32416 27068 32428
rect 24995 32388 27068 32416
rect 24995 32385 25007 32388
rect 24949 32379 25007 32385
rect 27062 32376 27068 32388
rect 27120 32376 27126 32428
rect 27154 32376 27160 32428
rect 27212 32416 27218 32428
rect 27893 32419 27951 32425
rect 27212 32388 27257 32416
rect 27212 32376 27218 32388
rect 27893 32385 27905 32419
rect 27939 32416 27951 32419
rect 28166 32416 28172 32428
rect 27939 32388 28172 32416
rect 27939 32385 27951 32388
rect 27893 32379 27951 32385
rect 28166 32376 28172 32388
rect 28224 32376 28230 32428
rect 29086 32376 29092 32428
rect 29144 32416 29150 32428
rect 29181 32419 29239 32425
rect 29181 32416 29193 32419
rect 29144 32388 29193 32416
rect 29144 32376 29150 32388
rect 29181 32385 29193 32388
rect 29227 32385 29239 32419
rect 29181 32379 29239 32385
rect 30009 32419 30067 32425
rect 30009 32385 30021 32419
rect 30055 32385 30067 32419
rect 30009 32379 30067 32385
rect 31021 32419 31079 32425
rect 31021 32385 31033 32419
rect 31067 32385 31079 32419
rect 31021 32379 31079 32385
rect 25222 32348 25228 32360
rect 23308 32320 25228 32348
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 29273 32351 29331 32357
rect 29273 32317 29285 32351
rect 29319 32348 29331 32351
rect 29362 32348 29368 32360
rect 29319 32320 29368 32348
rect 29319 32317 29331 32320
rect 29273 32311 29331 32317
rect 29362 32308 29368 32320
rect 29420 32308 29426 32360
rect 23216 32280 23244 32308
rect 27614 32280 27620 32292
rect 19935 32252 22094 32280
rect 23216 32252 27620 32280
rect 19935 32249 19947 32252
rect 19889 32243 19947 32249
rect 21082 32212 21088 32224
rect 21043 32184 21088 32212
rect 21082 32172 21088 32184
rect 21140 32172 21146 32224
rect 22066 32212 22094 32252
rect 27614 32240 27620 32252
rect 27672 32240 27678 32292
rect 28258 32240 28264 32292
rect 28316 32280 28322 32292
rect 30024 32280 30052 32379
rect 28316 32252 30052 32280
rect 28316 32240 28322 32252
rect 23109 32215 23167 32221
rect 23109 32212 23121 32215
rect 22066 32184 23121 32212
rect 23109 32181 23121 32184
rect 23155 32181 23167 32215
rect 24394 32212 24400 32224
rect 24355 32184 24400 32212
rect 23109 32175 23167 32181
rect 24394 32172 24400 32184
rect 24452 32172 24458 32224
rect 26326 32172 26332 32224
rect 26384 32212 26390 32224
rect 26973 32215 27031 32221
rect 26973 32212 26985 32215
rect 26384 32184 26985 32212
rect 26384 32172 26390 32184
rect 26973 32181 26985 32184
rect 27019 32181 27031 32215
rect 26973 32175 27031 32181
rect 27154 32172 27160 32224
rect 27212 32212 27218 32224
rect 27985 32215 28043 32221
rect 27985 32212 27997 32215
rect 27212 32184 27997 32212
rect 27212 32172 27218 32184
rect 27985 32181 27997 32184
rect 28031 32181 28043 32215
rect 27985 32175 28043 32181
rect 29549 32215 29607 32221
rect 29549 32181 29561 32215
rect 29595 32212 29607 32215
rect 29914 32212 29920 32224
rect 29595 32184 29920 32212
rect 29595 32181 29607 32184
rect 29549 32175 29607 32181
rect 29914 32172 29920 32184
rect 29972 32172 29978 32224
rect 31036 32212 31064 32379
rect 31110 32376 31116 32428
rect 31168 32416 31174 32428
rect 31205 32419 31263 32425
rect 31205 32416 31217 32419
rect 31168 32388 31217 32416
rect 31168 32376 31174 32388
rect 31205 32385 31217 32388
rect 31251 32385 31263 32419
rect 31205 32379 31263 32385
rect 31389 32419 31447 32425
rect 31389 32385 31401 32419
rect 31435 32416 31447 32419
rect 31478 32416 31484 32428
rect 31435 32388 31484 32416
rect 31435 32385 31447 32388
rect 31389 32379 31447 32385
rect 31478 32376 31484 32388
rect 31536 32376 31542 32428
rect 32122 32416 32128 32428
rect 32083 32388 32128 32416
rect 32122 32376 32128 32388
rect 32180 32376 32186 32428
rect 46474 32376 46480 32428
rect 46532 32416 46538 32428
rect 47581 32419 47639 32425
rect 47581 32416 47593 32419
rect 46532 32388 47593 32416
rect 46532 32376 46538 32388
rect 47581 32385 47593 32388
rect 47627 32385 47639 32419
rect 47581 32379 47639 32385
rect 32766 32212 32772 32224
rect 31036 32184 32772 32212
rect 32766 32172 32772 32184
rect 32824 32212 32830 32224
rect 33873 32215 33931 32221
rect 33873 32212 33885 32215
rect 32824 32184 33885 32212
rect 32824 32172 32830 32184
rect 33873 32181 33885 32184
rect 33919 32181 33931 32215
rect 33873 32175 33931 32181
rect 46474 32172 46480 32224
rect 46532 32212 46538 32224
rect 47673 32215 47731 32221
rect 47673 32212 47685 32215
rect 46532 32184 47685 32212
rect 46532 32172 46538 32184
rect 47673 32181 47685 32184
rect 47719 32181 47731 32215
rect 47673 32175 47731 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1670 32008 1676 32020
rect 1631 31980 1676 32008
rect 1670 31968 1676 31980
rect 1728 31968 1734 32020
rect 2222 32008 2228 32020
rect 2183 31980 2228 32008
rect 2222 31968 2228 31980
rect 2280 31968 2286 32020
rect 19426 32008 19432 32020
rect 19387 31980 19432 32008
rect 19426 31968 19432 31980
rect 19484 31968 19490 32020
rect 21910 32008 21916 32020
rect 21871 31980 21916 32008
rect 21910 31968 21916 31980
rect 21968 32008 21974 32020
rect 22649 32011 22707 32017
rect 22649 32008 22661 32011
rect 21968 31980 22661 32008
rect 21968 31968 21974 31980
rect 22649 31977 22661 31980
rect 22695 31977 22707 32011
rect 24762 32008 24768 32020
rect 24723 31980 24768 32008
rect 22649 31971 22707 31977
rect 24762 31968 24768 31980
rect 24820 31968 24826 32020
rect 25222 32008 25228 32020
rect 25183 31980 25228 32008
rect 25222 31968 25228 31980
rect 25280 31968 25286 32020
rect 28994 32008 29000 32020
rect 26068 31980 29000 32008
rect 22189 31943 22247 31949
rect 22189 31909 22201 31943
rect 22235 31940 22247 31943
rect 23934 31940 23940 31952
rect 22235 31912 23940 31940
rect 22235 31909 22247 31912
rect 22189 31903 22247 31909
rect 23934 31900 23940 31912
rect 23992 31900 23998 31952
rect 2682 31832 2688 31884
rect 2740 31872 2746 31884
rect 3973 31875 4031 31881
rect 3973 31872 3985 31875
rect 2740 31844 3985 31872
rect 2740 31832 2746 31844
rect 3973 31841 3985 31844
rect 4019 31841 4031 31875
rect 4614 31872 4620 31884
rect 4575 31844 4620 31872
rect 3973 31835 4031 31841
rect 4614 31832 4620 31844
rect 4672 31872 4678 31884
rect 5442 31872 5448 31884
rect 4672 31844 5448 31872
rect 4672 31832 4678 31844
rect 5442 31832 5448 31844
rect 5500 31832 5506 31884
rect 21266 31832 21272 31884
rect 21324 31872 21330 31884
rect 21913 31875 21971 31881
rect 21913 31872 21925 31875
rect 21324 31844 21925 31872
rect 21324 31832 21330 31844
rect 21913 31841 21925 31844
rect 21959 31841 21971 31875
rect 21913 31835 21971 31841
rect 22833 31875 22891 31881
rect 22833 31841 22845 31875
rect 22879 31872 22891 31875
rect 24394 31872 24400 31884
rect 22879 31844 24400 31872
rect 22879 31841 22891 31844
rect 22833 31835 22891 31841
rect 2133 31807 2191 31813
rect 2133 31773 2145 31807
rect 2179 31804 2191 31807
rect 2314 31804 2320 31816
rect 2179 31776 2320 31804
rect 2179 31773 2191 31776
rect 2133 31767 2191 31773
rect 2314 31764 2320 31776
rect 2372 31764 2378 31816
rect 3786 31804 3792 31816
rect 3747 31776 3792 31804
rect 3786 31764 3792 31776
rect 3844 31764 3850 31816
rect 17773 31807 17831 31813
rect 17773 31773 17785 31807
rect 17819 31804 17831 31807
rect 18138 31804 18144 31816
rect 17819 31776 18144 31804
rect 17819 31773 17831 31776
rect 17773 31767 17831 31773
rect 18138 31764 18144 31776
rect 18196 31764 18202 31816
rect 18233 31807 18291 31813
rect 18233 31773 18245 31807
rect 18279 31804 18291 31807
rect 18506 31804 18512 31816
rect 18279 31776 18512 31804
rect 18279 31773 18291 31776
rect 18233 31767 18291 31773
rect 18506 31764 18512 31776
rect 18564 31764 18570 31816
rect 19337 31807 19395 31813
rect 19337 31773 19349 31807
rect 19383 31804 19395 31807
rect 19978 31804 19984 31816
rect 19383 31776 19984 31804
rect 19383 31773 19395 31776
rect 19337 31767 19395 31773
rect 19978 31764 19984 31776
rect 20036 31764 20042 31816
rect 21082 31764 21088 31816
rect 21140 31804 21146 31816
rect 21821 31807 21879 31813
rect 21821 31804 21833 31807
rect 21140 31776 21833 31804
rect 21140 31764 21146 31776
rect 21821 31773 21833 31776
rect 21867 31773 21879 31807
rect 21928 31804 21956 31835
rect 24394 31832 24400 31844
rect 24452 31832 24458 31884
rect 24854 31872 24860 31884
rect 24815 31844 24860 31872
rect 24854 31832 24860 31844
rect 24912 31832 24918 31884
rect 26068 31881 26096 31980
rect 28994 31968 29000 31980
rect 29052 31968 29058 32020
rect 32493 32011 32551 32017
rect 32493 31977 32505 32011
rect 32539 32008 32551 32011
rect 32582 32008 32588 32020
rect 32539 31980 32588 32008
rect 32539 31977 32551 31980
rect 32493 31971 32551 31977
rect 32582 31968 32588 31980
rect 32640 31968 32646 32020
rect 33321 32011 33379 32017
rect 33321 31977 33333 32011
rect 33367 32008 33379 32011
rect 33410 32008 33416 32020
rect 33367 31980 33416 32008
rect 33367 31977 33379 31980
rect 33321 31971 33379 31977
rect 33410 31968 33416 31980
rect 33468 31968 33474 32020
rect 48038 32008 48044 32020
rect 41386 31980 48044 32008
rect 41386 31940 41414 31980
rect 48038 31968 48044 31980
rect 48096 31968 48102 32020
rect 31726 31912 41414 31940
rect 26053 31875 26111 31881
rect 26053 31841 26065 31875
rect 26099 31841 26111 31875
rect 26326 31872 26332 31884
rect 26287 31844 26332 31872
rect 26053 31835 26111 31841
rect 26326 31832 26332 31844
rect 26384 31832 26390 31884
rect 27338 31832 27344 31884
rect 27396 31872 27402 31884
rect 27522 31872 27528 31884
rect 27396 31844 27528 31872
rect 27396 31832 27402 31844
rect 27522 31832 27528 31844
rect 27580 31872 27586 31884
rect 27801 31875 27859 31881
rect 27801 31872 27813 31875
rect 27580 31844 27813 31872
rect 27580 31832 27586 31844
rect 27801 31841 27813 31844
rect 27847 31841 27859 31875
rect 27801 31835 27859 31841
rect 27982 31832 27988 31884
rect 28040 31872 28046 31884
rect 31726 31872 31754 31912
rect 28040 31844 31754 31872
rect 32125 31875 32183 31881
rect 28040 31832 28046 31844
rect 32125 31841 32137 31875
rect 32171 31841 32183 31875
rect 46290 31872 46296 31884
rect 46251 31844 46296 31872
rect 32125 31835 32183 31841
rect 22925 31807 22983 31813
rect 22925 31804 22937 31807
rect 21928 31776 22937 31804
rect 21821 31767 21879 31773
rect 22925 31773 22937 31776
rect 22971 31804 22983 31807
rect 23382 31804 23388 31816
rect 22971 31776 23388 31804
rect 22971 31773 22983 31776
rect 22925 31767 22983 31773
rect 21836 31736 21864 31767
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 24118 31764 24124 31816
rect 24176 31804 24182 31816
rect 24765 31807 24823 31813
rect 24765 31804 24777 31807
rect 24176 31776 24777 31804
rect 24176 31764 24182 31776
rect 24765 31773 24777 31776
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 25041 31807 25099 31813
rect 25041 31773 25053 31807
rect 25087 31804 25099 31807
rect 25087 31776 26096 31804
rect 27462 31776 28212 31804
rect 25087 31773 25099 31776
rect 25041 31767 25099 31773
rect 22094 31736 22100 31748
rect 21836 31708 22100 31736
rect 22094 31696 22100 31708
rect 22152 31736 22158 31748
rect 22649 31739 22707 31745
rect 22649 31736 22661 31739
rect 22152 31708 22661 31736
rect 22152 31696 22158 31708
rect 22649 31705 22661 31708
rect 22695 31736 22707 31739
rect 23290 31736 23296 31748
rect 22695 31708 23296 31736
rect 22695 31705 22707 31708
rect 22649 31699 22707 31705
rect 23290 31696 23296 31708
rect 23348 31696 23354 31748
rect 26068 31736 26096 31776
rect 28184 31736 28212 31776
rect 28258 31764 28264 31816
rect 28316 31804 28322 31816
rect 29914 31804 29920 31816
rect 28316 31776 28361 31804
rect 29875 31776 29920 31804
rect 28316 31764 28322 31776
rect 29914 31764 29920 31776
rect 29972 31764 29978 31816
rect 30006 31764 30012 31816
rect 30064 31804 30070 31816
rect 30101 31807 30159 31813
rect 30101 31804 30113 31807
rect 30064 31776 30113 31804
rect 30064 31764 30070 31776
rect 30101 31773 30113 31776
rect 30147 31773 30159 31807
rect 30101 31767 30159 31773
rect 31478 31764 31484 31816
rect 31536 31804 31542 31816
rect 32140 31804 32168 31835
rect 46290 31832 46296 31844
rect 46348 31832 46354 31884
rect 46474 31872 46480 31884
rect 46435 31844 46480 31872
rect 46474 31832 46480 31844
rect 46532 31832 46538 31884
rect 48130 31872 48136 31884
rect 48091 31844 48136 31872
rect 48130 31832 48136 31844
rect 48188 31832 48194 31884
rect 31536 31776 32168 31804
rect 32217 31807 32275 31813
rect 31536 31764 31542 31776
rect 32217 31773 32229 31807
rect 32263 31804 32275 31807
rect 32582 31804 32588 31816
rect 32263 31776 32588 31804
rect 32263 31773 32275 31776
rect 32217 31767 32275 31773
rect 32582 31764 32588 31776
rect 32640 31804 32646 31816
rect 32766 31804 32772 31816
rect 32640 31776 32772 31804
rect 32640 31764 32646 31776
rect 32766 31764 32772 31776
rect 32824 31764 32830 31816
rect 33229 31807 33287 31813
rect 33229 31773 33241 31807
rect 33275 31804 33287 31807
rect 34606 31804 34612 31816
rect 33275 31776 34612 31804
rect 33275 31773 33287 31776
rect 33229 31767 33287 31773
rect 34606 31764 34612 31776
rect 34664 31764 34670 31816
rect 28353 31739 28411 31745
rect 28353 31736 28365 31739
rect 26068 31708 26280 31736
rect 28184 31708 28365 31736
rect 18325 31671 18383 31677
rect 18325 31637 18337 31671
rect 18371 31668 18383 31671
rect 18506 31668 18512 31680
rect 18371 31640 18512 31668
rect 18371 31637 18383 31640
rect 18325 31631 18383 31637
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 23109 31671 23167 31677
rect 23109 31637 23121 31671
rect 23155 31668 23167 31671
rect 23198 31668 23204 31680
rect 23155 31640 23204 31668
rect 23155 31637 23167 31640
rect 23109 31631 23167 31637
rect 23198 31628 23204 31640
rect 23256 31628 23262 31680
rect 26252 31668 26280 31708
rect 28353 31705 28365 31708
rect 28399 31705 28411 31739
rect 28353 31699 28411 31705
rect 27338 31668 27344 31680
rect 26252 31640 27344 31668
rect 27338 31628 27344 31640
rect 27396 31628 27402 31680
rect 28718 31628 28724 31680
rect 28776 31668 28782 31680
rect 30009 31671 30067 31677
rect 30009 31668 30021 31671
rect 28776 31640 30021 31668
rect 28776 31628 28782 31640
rect 30009 31637 30021 31640
rect 30055 31637 30067 31671
rect 30009 31631 30067 31637
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 24578 31424 24584 31476
rect 24636 31464 24642 31476
rect 24673 31467 24731 31473
rect 24673 31464 24685 31467
rect 24636 31436 24685 31464
rect 24636 31424 24642 31436
rect 24673 31433 24685 31436
rect 24719 31433 24731 31467
rect 24673 31427 24731 31433
rect 27062 31424 27068 31476
rect 27120 31464 27126 31476
rect 28629 31467 28687 31473
rect 28629 31464 28641 31467
rect 27120 31436 28641 31464
rect 27120 31424 27126 31436
rect 28629 31433 28641 31436
rect 28675 31464 28687 31467
rect 28675 31436 29684 31464
rect 28675 31433 28687 31436
rect 28629 31427 28687 31433
rect 18506 31396 18512 31408
rect 18467 31368 18512 31396
rect 18506 31356 18512 31368
rect 18564 31356 18570 31408
rect 24854 31396 24860 31408
rect 23768 31368 24860 31396
rect 18138 31288 18144 31340
rect 18196 31328 18202 31340
rect 18325 31331 18383 31337
rect 18325 31328 18337 31331
rect 18196 31300 18337 31328
rect 18196 31288 18202 31300
rect 18325 31297 18337 31300
rect 18371 31297 18383 31331
rect 18325 31291 18383 31297
rect 21910 31288 21916 31340
rect 21968 31328 21974 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21968 31300 22017 31328
rect 21968 31288 21974 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22833 31331 22891 31337
rect 22833 31328 22845 31331
rect 22005 31291 22063 31297
rect 22388 31300 22845 31328
rect 20165 31263 20223 31269
rect 20165 31229 20177 31263
rect 20211 31260 20223 31263
rect 20254 31260 20260 31272
rect 20211 31232 20260 31260
rect 20211 31229 20223 31232
rect 20165 31223 20223 31229
rect 20254 31220 20260 31232
rect 20312 31220 20318 31272
rect 22094 31260 22100 31272
rect 22055 31232 22100 31260
rect 22094 31220 22100 31232
rect 22152 31220 22158 31272
rect 22388 31269 22416 31300
rect 22833 31297 22845 31300
rect 22879 31297 22891 31331
rect 22833 31291 22891 31297
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31328 23075 31331
rect 23106 31328 23112 31340
rect 23063 31300 23112 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 23106 31288 23112 31300
rect 23164 31288 23170 31340
rect 23768 31337 23796 31368
rect 24854 31356 24860 31368
rect 24912 31356 24918 31408
rect 26053 31399 26111 31405
rect 26053 31365 26065 31399
rect 26099 31365 26111 31399
rect 26053 31359 26111 31365
rect 23753 31331 23811 31337
rect 23753 31297 23765 31331
rect 23799 31297 23811 31331
rect 23934 31328 23940 31340
rect 23895 31300 23940 31328
rect 23753 31291 23811 31297
rect 23934 31288 23940 31300
rect 23992 31288 23998 31340
rect 24029 31331 24087 31337
rect 24029 31297 24041 31331
rect 24075 31328 24087 31331
rect 24118 31328 24124 31340
rect 24075 31300 24124 31328
rect 24075 31297 24087 31300
rect 24029 31291 24087 31297
rect 24118 31288 24124 31300
rect 24176 31288 24182 31340
rect 24578 31328 24584 31340
rect 24539 31300 24584 31328
rect 24578 31288 24584 31300
rect 24636 31288 24642 31340
rect 26068 31328 26096 31359
rect 26142 31356 26148 31408
rect 26200 31396 26206 31408
rect 29656 31405 29684 31436
rect 26253 31399 26311 31405
rect 26253 31396 26265 31399
rect 26200 31368 26265 31396
rect 26200 31356 26206 31368
rect 26253 31365 26265 31368
rect 26299 31365 26311 31399
rect 26253 31359 26311 31365
rect 29641 31399 29699 31405
rect 29641 31365 29653 31399
rect 29687 31365 29699 31399
rect 29641 31359 29699 31365
rect 26694 31328 26700 31340
rect 26068 31300 26700 31328
rect 26694 31288 26700 31300
rect 26752 31328 26758 31340
rect 27154 31328 27160 31340
rect 26752 31300 27160 31328
rect 26752 31288 26758 31300
rect 27154 31288 27160 31300
rect 27212 31288 27218 31340
rect 27338 31328 27344 31340
rect 27299 31300 27344 31328
rect 27338 31288 27344 31300
rect 27396 31288 27402 31340
rect 27614 31288 27620 31340
rect 27672 31328 27678 31340
rect 30837 31331 30895 31337
rect 30837 31328 30849 31331
rect 27672 31300 30849 31328
rect 27672 31288 27678 31300
rect 30837 31297 30849 31300
rect 30883 31297 30895 31331
rect 30837 31291 30895 31297
rect 22373 31263 22431 31269
rect 22373 31229 22385 31263
rect 22419 31229 22431 31263
rect 22373 31223 22431 31229
rect 31205 31263 31263 31269
rect 31205 31229 31217 31263
rect 31251 31260 31263 31263
rect 31478 31260 31484 31272
rect 31251 31232 31484 31260
rect 31251 31229 31263 31232
rect 31205 31223 31263 31229
rect 31478 31220 31484 31232
rect 31536 31220 31542 31272
rect 22833 31195 22891 31201
rect 22833 31192 22845 31195
rect 22296 31164 22845 31192
rect 21818 31084 21824 31136
rect 21876 31124 21882 31136
rect 22296 31124 22324 31164
rect 22833 31161 22845 31164
rect 22879 31161 22891 31195
rect 22833 31155 22891 31161
rect 23290 31152 23296 31204
rect 23348 31192 23354 31204
rect 29825 31195 29883 31201
rect 23348 31164 28994 31192
rect 23348 31152 23354 31164
rect 21876 31096 22324 31124
rect 21876 31084 21882 31096
rect 23474 31084 23480 31136
rect 23532 31124 23538 31136
rect 23569 31127 23627 31133
rect 23569 31124 23581 31127
rect 23532 31096 23581 31124
rect 23532 31084 23538 31096
rect 23569 31093 23581 31096
rect 23615 31093 23627 31127
rect 26234 31124 26240 31136
rect 26195 31096 26240 31124
rect 23569 31087 23627 31093
rect 26234 31084 26240 31096
rect 26292 31084 26298 31136
rect 26421 31127 26479 31133
rect 26421 31093 26433 31127
rect 26467 31124 26479 31127
rect 27062 31124 27068 31136
rect 26467 31096 27068 31124
rect 26467 31093 26479 31096
rect 26421 31087 26479 31093
rect 27062 31084 27068 31096
rect 27120 31084 27126 31136
rect 28966 31124 28994 31164
rect 29825 31161 29837 31195
rect 29871 31192 29883 31195
rect 30558 31192 30564 31204
rect 29871 31164 30564 31192
rect 29871 31161 29883 31164
rect 29825 31155 29883 31161
rect 30558 31152 30564 31164
rect 30616 31152 30622 31204
rect 31297 31195 31355 31201
rect 31297 31192 31309 31195
rect 30668 31164 31309 31192
rect 30668 31124 30696 31164
rect 31297 31161 31309 31164
rect 31343 31161 31355 31195
rect 31297 31155 31355 31161
rect 31018 31133 31024 31136
rect 28966 31096 30696 31124
rect 31002 31127 31024 31133
rect 31002 31093 31014 31127
rect 31002 31087 31024 31093
rect 31018 31084 31024 31087
rect 31076 31084 31082 31136
rect 31110 31084 31116 31136
rect 31168 31124 31174 31136
rect 31168 31096 31213 31124
rect 31168 31084 31174 31096
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 20530 30880 20536 30932
rect 20588 30920 20594 30932
rect 22465 30923 22523 30929
rect 22465 30920 22477 30923
rect 20588 30892 22477 30920
rect 20588 30880 20594 30892
rect 22465 30889 22477 30892
rect 22511 30889 22523 30923
rect 22465 30883 22523 30889
rect 23569 30923 23627 30929
rect 23569 30889 23581 30923
rect 23615 30920 23627 30923
rect 23934 30920 23940 30932
rect 23615 30892 23940 30920
rect 23615 30889 23627 30892
rect 23569 30883 23627 30889
rect 23934 30880 23940 30892
rect 23992 30880 23998 30932
rect 25314 30880 25320 30932
rect 25372 30920 25378 30932
rect 25777 30923 25835 30929
rect 25777 30920 25789 30923
rect 25372 30892 25789 30920
rect 25372 30880 25378 30892
rect 25777 30889 25789 30892
rect 25823 30920 25835 30923
rect 26142 30920 26148 30932
rect 25823 30892 26148 30920
rect 25823 30889 25835 30892
rect 25777 30883 25835 30889
rect 26142 30880 26148 30892
rect 26200 30880 26206 30932
rect 27430 30880 27436 30932
rect 27488 30920 27494 30932
rect 27525 30923 27583 30929
rect 27525 30920 27537 30923
rect 27488 30892 27537 30920
rect 27488 30880 27494 30892
rect 27525 30889 27537 30892
rect 27571 30889 27583 30923
rect 27525 30883 27583 30889
rect 28169 30923 28227 30929
rect 28169 30889 28181 30923
rect 28215 30920 28227 30923
rect 31754 30920 31760 30932
rect 28215 30892 31760 30920
rect 28215 30889 28227 30892
rect 28169 30883 28227 30889
rect 31754 30880 31760 30892
rect 31812 30920 31818 30932
rect 32490 30920 32496 30932
rect 31812 30892 32496 30920
rect 31812 30880 31818 30892
rect 32490 30880 32496 30892
rect 32548 30880 32554 30932
rect 29086 30812 29092 30864
rect 29144 30852 29150 30864
rect 29144 30824 29684 30852
rect 29144 30812 29150 30824
rect 20441 30787 20499 30793
rect 20441 30753 20453 30787
rect 20487 30784 20499 30787
rect 21082 30784 21088 30796
rect 20487 30756 21088 30784
rect 20487 30753 20499 30756
rect 20441 30747 20499 30753
rect 21082 30744 21088 30756
rect 21140 30744 21146 30796
rect 23474 30784 23480 30796
rect 22204 30756 23336 30784
rect 23435 30756 23480 30784
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30716 20407 30719
rect 21174 30716 21180 30728
rect 20395 30688 21180 30716
rect 20395 30685 20407 30688
rect 20349 30679 20407 30685
rect 21174 30676 21180 30688
rect 21232 30676 21238 30728
rect 21818 30716 21824 30728
rect 21779 30688 21824 30716
rect 21818 30676 21824 30688
rect 21876 30676 21882 30728
rect 21910 30676 21916 30728
rect 21968 30716 21974 30728
rect 22204 30725 22232 30756
rect 22189 30719 22247 30725
rect 21968 30688 22013 30716
rect 21968 30676 21974 30688
rect 22189 30685 22201 30719
rect 22235 30685 22247 30719
rect 22189 30679 22247 30685
rect 22286 30719 22344 30725
rect 22286 30685 22298 30719
rect 22332 30685 22344 30719
rect 23198 30716 23204 30728
rect 23159 30688 23204 30716
rect 22286 30679 22344 30685
rect 22002 30608 22008 30660
rect 22060 30648 22066 30660
rect 22097 30651 22155 30657
rect 22097 30648 22109 30651
rect 22060 30620 22109 30648
rect 22060 30608 22066 30620
rect 22097 30617 22109 30620
rect 22143 30617 22155 30651
rect 22097 30611 22155 30617
rect 20717 30583 20775 30589
rect 20717 30549 20729 30583
rect 20763 30580 20775 30583
rect 20806 30580 20812 30592
rect 20763 30552 20812 30580
rect 20763 30549 20775 30552
rect 20717 30543 20775 30549
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 20898 30540 20904 30592
rect 20956 30580 20962 30592
rect 22296 30580 22324 30679
rect 23198 30676 23204 30688
rect 23256 30676 23262 30728
rect 23308 30716 23336 30756
rect 23474 30744 23480 30756
rect 23532 30744 23538 30796
rect 24762 30744 24768 30796
rect 24820 30784 24826 30796
rect 24949 30787 25007 30793
rect 24949 30784 24961 30787
rect 24820 30756 24961 30784
rect 24820 30744 24826 30756
rect 24949 30753 24961 30756
rect 24995 30784 25007 30787
rect 27062 30784 27068 30796
rect 24995 30756 26004 30784
rect 27023 30756 27068 30784
rect 24995 30753 25007 30756
rect 24949 30747 25007 30753
rect 23842 30716 23848 30728
rect 23308 30688 23848 30716
rect 23842 30676 23848 30688
rect 23900 30676 23906 30728
rect 25976 30725 26004 30756
rect 27062 30744 27068 30756
rect 27120 30744 27126 30796
rect 28994 30744 29000 30796
rect 29052 30784 29058 30796
rect 29549 30787 29607 30793
rect 29549 30784 29561 30787
rect 29052 30756 29561 30784
rect 29052 30744 29058 30756
rect 29549 30753 29561 30756
rect 29595 30753 29607 30787
rect 29656 30784 29684 30824
rect 31018 30812 31024 30864
rect 31076 30852 31082 30864
rect 33321 30855 33379 30861
rect 33321 30852 33333 30855
rect 31076 30824 33333 30852
rect 31076 30812 31082 30824
rect 30834 30784 30840 30796
rect 29656 30756 30840 30784
rect 29549 30747 29607 30753
rect 30834 30744 30840 30756
rect 30892 30784 30898 30796
rect 31297 30787 31355 30793
rect 31297 30784 31309 30787
rect 30892 30756 31309 30784
rect 30892 30744 30898 30756
rect 31297 30753 31309 30756
rect 31343 30753 31355 30787
rect 31726 30784 31754 30824
rect 33321 30821 33333 30824
rect 33367 30821 33379 30855
rect 33321 30815 33379 30821
rect 31726 30756 31800 30784
rect 31297 30747 31355 30753
rect 25133 30719 25191 30725
rect 25133 30685 25145 30719
rect 25179 30716 25191 30719
rect 25777 30719 25835 30725
rect 25777 30716 25789 30719
rect 25179 30688 25789 30716
rect 25179 30685 25191 30688
rect 25133 30679 25191 30685
rect 25777 30685 25789 30688
rect 25823 30685 25835 30719
rect 25777 30679 25835 30685
rect 25961 30719 26019 30725
rect 25961 30685 25973 30719
rect 26007 30716 26019 30719
rect 26050 30716 26056 30728
rect 26007 30688 26056 30716
rect 26007 30685 26019 30688
rect 25961 30679 26019 30685
rect 23216 30648 23244 30676
rect 25148 30648 25176 30679
rect 26050 30676 26056 30688
rect 26108 30676 26114 30728
rect 27157 30719 27215 30725
rect 27157 30685 27169 30719
rect 27203 30716 27215 30719
rect 27522 30716 27528 30728
rect 27203 30688 27528 30716
rect 27203 30685 27215 30688
rect 27157 30679 27215 30685
rect 27522 30676 27528 30688
rect 27580 30676 27586 30728
rect 27706 30676 27712 30728
rect 27764 30716 27770 30728
rect 27985 30719 28043 30725
rect 27985 30716 27997 30719
rect 27764 30688 27997 30716
rect 27764 30676 27770 30688
rect 27985 30685 27997 30688
rect 28031 30716 28043 30719
rect 28074 30716 28080 30728
rect 28031 30688 28080 30716
rect 28031 30685 28043 30688
rect 27985 30679 28043 30685
rect 28074 30676 28080 30688
rect 28132 30676 28138 30728
rect 28258 30676 28264 30728
rect 28316 30716 28322 30728
rect 28626 30716 28632 30728
rect 28316 30688 28632 30716
rect 28316 30676 28322 30688
rect 28626 30676 28632 30688
rect 28684 30716 28690 30728
rect 31772 30725 31800 30756
rect 31938 30744 31944 30796
rect 31996 30784 32002 30796
rect 32217 30787 32275 30793
rect 32217 30784 32229 30787
rect 31996 30756 32229 30784
rect 31996 30744 32002 30756
rect 32217 30753 32229 30756
rect 32263 30784 32275 30787
rect 32582 30784 32588 30796
rect 32263 30756 32588 30784
rect 32263 30753 32275 30756
rect 32217 30747 32275 30753
rect 32582 30744 32588 30756
rect 32640 30744 32646 30796
rect 33042 30744 33048 30796
rect 33100 30784 33106 30796
rect 34701 30787 34759 30793
rect 34701 30784 34713 30787
rect 33100 30756 34713 30784
rect 33100 30744 33106 30756
rect 34701 30753 34713 30756
rect 34747 30753 34759 30787
rect 47670 30784 47676 30796
rect 47631 30756 47676 30784
rect 34701 30747 34759 30753
rect 47670 30744 47676 30756
rect 47728 30784 47734 30796
rect 48038 30784 48044 30796
rect 47728 30756 48044 30784
rect 47728 30744 47734 30756
rect 48038 30744 48044 30756
rect 48096 30744 48102 30796
rect 28813 30719 28871 30725
rect 28813 30716 28825 30719
rect 28684 30688 28825 30716
rect 28684 30676 28690 30688
rect 28813 30685 28825 30688
rect 28859 30685 28871 30719
rect 28813 30679 28871 30685
rect 31757 30719 31815 30725
rect 31757 30685 31769 30719
rect 31803 30685 31815 30719
rect 31757 30679 31815 30685
rect 31849 30719 31907 30725
rect 31849 30685 31861 30719
rect 31895 30685 31907 30719
rect 32030 30716 32036 30728
rect 31991 30688 32036 30716
rect 31849 30679 31907 30685
rect 23216 30620 25176 30648
rect 25590 30608 25596 30660
rect 25648 30648 25654 30660
rect 28276 30648 28304 30676
rect 29822 30648 29828 30660
rect 25648 30620 28304 30648
rect 29783 30620 29828 30648
rect 25648 30608 25654 30620
rect 29822 30608 29828 30620
rect 29880 30608 29886 30660
rect 29932 30620 30314 30648
rect 23750 30580 23756 30592
rect 20956 30552 22324 30580
rect 23711 30552 23756 30580
rect 20956 30540 20962 30552
rect 23750 30540 23756 30552
rect 23808 30540 23814 30592
rect 25222 30540 25228 30592
rect 25280 30580 25286 30592
rect 25317 30583 25375 30589
rect 25317 30580 25329 30583
rect 25280 30552 25329 30580
rect 25280 30540 25286 30552
rect 25317 30549 25329 30552
rect 25363 30549 25375 30583
rect 25317 30543 25375 30549
rect 28905 30583 28963 30589
rect 28905 30549 28917 30583
rect 28951 30580 28963 30583
rect 29932 30580 29960 30620
rect 31110 30608 31116 30660
rect 31168 30648 31174 30660
rect 31570 30648 31576 30660
rect 31168 30620 31576 30648
rect 31168 30608 31174 30620
rect 31570 30608 31576 30620
rect 31628 30648 31634 30660
rect 31864 30648 31892 30679
rect 32030 30676 32036 30688
rect 32088 30676 32094 30728
rect 33137 30719 33195 30725
rect 33137 30685 33149 30719
rect 33183 30716 33195 30719
rect 33686 30716 33692 30728
rect 33183 30688 33692 30716
rect 33183 30685 33195 30688
rect 33137 30679 33195 30685
rect 33686 30676 33692 30688
rect 33744 30716 33750 30728
rect 33781 30719 33839 30725
rect 33781 30716 33793 30719
rect 33744 30688 33793 30716
rect 33744 30676 33750 30688
rect 33781 30685 33793 30688
rect 33827 30716 33839 30719
rect 33827 30688 34284 30716
rect 33827 30685 33839 30688
rect 33781 30679 33839 30685
rect 31628 30620 31892 30648
rect 31628 30608 31634 30620
rect 32674 30608 32680 30660
rect 32732 30648 32738 30660
rect 32953 30651 33011 30657
rect 32953 30648 32965 30651
rect 32732 30620 32965 30648
rect 32732 30608 32738 30620
rect 32953 30617 32965 30620
rect 32999 30617 33011 30651
rect 32953 30611 33011 30617
rect 33870 30580 33876 30592
rect 28951 30552 29960 30580
rect 33831 30552 33876 30580
rect 28951 30549 28963 30552
rect 28905 30543 28963 30549
rect 33870 30540 33876 30552
rect 33928 30540 33934 30592
rect 34256 30580 34284 30688
rect 34514 30608 34520 30660
rect 34572 30648 34578 30660
rect 34977 30651 35035 30657
rect 34977 30648 34989 30651
rect 34572 30620 34989 30648
rect 34572 30608 34578 30620
rect 34977 30617 34989 30620
rect 35023 30617 35035 30651
rect 34977 30611 35035 30617
rect 35986 30608 35992 30660
rect 36044 30608 36050 30660
rect 46106 30608 46112 30660
rect 46164 30648 46170 30660
rect 46845 30651 46903 30657
rect 46845 30648 46857 30651
rect 46164 30620 46857 30648
rect 46164 30608 46170 30620
rect 46845 30617 46857 30620
rect 46891 30617 46903 30651
rect 46845 30611 46903 30617
rect 46937 30651 46995 30657
rect 46937 30617 46949 30651
rect 46983 30648 46995 30651
rect 47302 30648 47308 30660
rect 46983 30620 47308 30648
rect 46983 30617 46995 30620
rect 46937 30611 46995 30617
rect 47302 30608 47308 30620
rect 47360 30648 47366 30660
rect 47946 30648 47952 30660
rect 47360 30620 47952 30648
rect 47360 30608 47366 30620
rect 47946 30608 47952 30620
rect 48004 30608 48010 30660
rect 36449 30583 36507 30589
rect 36449 30580 36461 30583
rect 34256 30552 36461 30580
rect 36449 30549 36461 30552
rect 36495 30549 36507 30583
rect 36449 30543 36507 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 4614 30336 4620 30388
rect 4672 30376 4678 30388
rect 20898 30376 20904 30388
rect 4672 30348 20904 30376
rect 4672 30336 4678 30348
rect 20898 30336 20904 30348
rect 20956 30336 20962 30388
rect 27249 30379 27307 30385
rect 27249 30376 27261 30379
rect 27172 30348 27261 30376
rect 23658 30308 23664 30320
rect 20732 30280 23664 30308
rect 14090 30200 14096 30252
rect 14148 30240 14154 30252
rect 15105 30243 15163 30249
rect 15105 30240 15117 30243
rect 14148 30212 15117 30240
rect 14148 30200 14154 30212
rect 15105 30209 15117 30212
rect 15151 30240 15163 30243
rect 17310 30240 17316 30252
rect 15151 30212 17316 30240
rect 15151 30209 15163 30212
rect 15105 30203 15163 30209
rect 17310 30200 17316 30212
rect 17368 30200 17374 30252
rect 19334 30200 19340 30252
rect 19392 30240 19398 30252
rect 19705 30243 19763 30249
rect 19705 30240 19717 30243
rect 19392 30212 19717 30240
rect 19392 30200 19398 30212
rect 19705 30209 19717 30212
rect 19751 30209 19763 30243
rect 19705 30203 19763 30209
rect 20533 30243 20591 30249
rect 20533 30209 20545 30243
rect 20579 30240 20591 30243
rect 20622 30240 20628 30252
rect 20579 30212 20628 30240
rect 20579 30209 20591 30212
rect 20533 30203 20591 30209
rect 20622 30200 20628 30212
rect 20680 30200 20686 30252
rect 20732 30249 20760 30280
rect 23658 30268 23664 30280
rect 23716 30308 23722 30320
rect 24121 30311 24179 30317
rect 23716 30280 24072 30308
rect 23716 30268 23722 30280
rect 20717 30243 20775 30249
rect 20717 30209 20729 30243
rect 20763 30209 20775 30243
rect 20717 30203 20775 30209
rect 20806 30200 20812 30252
rect 20864 30240 20870 30252
rect 21085 30243 21143 30249
rect 20864 30212 20909 30240
rect 20864 30200 20870 30212
rect 21085 30209 21097 30243
rect 21131 30240 21143 30243
rect 21174 30240 21180 30252
rect 21131 30212 21180 30240
rect 21131 30209 21143 30212
rect 21085 30203 21143 30209
rect 21174 30200 21180 30212
rect 21232 30200 21238 30252
rect 17402 30172 17408 30184
rect 17363 30144 17408 30172
rect 17402 30132 17408 30144
rect 17460 30132 17466 30184
rect 17586 30172 17592 30184
rect 17547 30144 17592 30172
rect 17586 30132 17592 30144
rect 17644 30132 17650 30184
rect 19245 30175 19303 30181
rect 19245 30141 19257 30175
rect 19291 30141 19303 30175
rect 19245 30135 19303 30141
rect 20901 30175 20959 30181
rect 20901 30141 20913 30175
rect 20947 30172 20959 30175
rect 20990 30172 20996 30184
rect 20947 30144 20996 30172
rect 20947 30141 20959 30144
rect 20901 30135 20959 30141
rect 19260 30104 19288 30135
rect 20990 30132 20996 30144
rect 21048 30172 21054 30184
rect 23198 30172 23204 30184
rect 21048 30144 23204 30172
rect 21048 30132 21054 30144
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 24044 30172 24072 30280
rect 24121 30277 24133 30311
rect 24167 30308 24179 30311
rect 24946 30308 24952 30320
rect 24167 30280 24952 30308
rect 24167 30277 24179 30280
rect 24121 30271 24179 30277
rect 24946 30268 24952 30280
rect 25004 30268 25010 30320
rect 25130 30308 25136 30320
rect 25056 30280 25136 30308
rect 25056 30249 25084 30280
rect 25130 30268 25136 30280
rect 25188 30268 25194 30320
rect 27172 30308 27200 30348
rect 27249 30345 27261 30348
rect 27295 30345 27307 30379
rect 27249 30339 27307 30345
rect 29549 30379 29607 30385
rect 29549 30345 29561 30379
rect 29595 30376 29607 30379
rect 29822 30376 29828 30388
rect 29595 30348 29828 30376
rect 29595 30345 29607 30348
rect 29549 30339 29607 30345
rect 29822 30336 29828 30348
rect 29880 30336 29886 30388
rect 29270 30308 29276 30320
rect 26068 30280 27200 30308
rect 29231 30280 29276 30308
rect 25041 30243 25099 30249
rect 25041 30209 25053 30243
rect 25087 30209 25099 30243
rect 25222 30240 25228 30252
rect 25183 30212 25228 30240
rect 25041 30203 25099 30209
rect 25222 30200 25228 30212
rect 25280 30200 25286 30252
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 25372 30212 25417 30240
rect 25372 30200 25378 30212
rect 26068 30172 26096 30280
rect 29270 30268 29276 30280
rect 29328 30268 29334 30320
rect 30466 30268 30472 30320
rect 30524 30308 30530 30320
rect 34149 30311 34207 30317
rect 30524 30280 33640 30308
rect 30524 30268 30530 30280
rect 27062 30240 27068 30252
rect 27023 30212 27068 30240
rect 27062 30200 27068 30212
rect 27120 30200 27126 30252
rect 28166 30240 28172 30252
rect 28127 30212 28172 30240
rect 28166 30200 28172 30212
rect 28224 30200 28230 30252
rect 28718 30200 28724 30252
rect 28776 30240 28782 30252
rect 29086 30249 29092 30254
rect 28912 30243 28970 30249
rect 28912 30240 28924 30243
rect 28776 30212 28924 30240
rect 28776 30200 28782 30212
rect 28912 30209 28924 30212
rect 28958 30209 28970 30243
rect 28912 30203 28970 30209
rect 29043 30243 29092 30249
rect 29043 30209 29055 30243
rect 29089 30209 29092 30243
rect 29043 30203 29092 30209
rect 29086 30202 29092 30203
rect 29144 30202 29150 30254
rect 29178 30200 29184 30252
rect 29236 30240 29242 30252
rect 29454 30249 29460 30252
rect 29411 30243 29460 30249
rect 29236 30212 29281 30240
rect 29236 30200 29242 30212
rect 29411 30209 29423 30243
rect 29457 30209 29460 30243
rect 29411 30203 29460 30209
rect 29454 30200 29460 30203
rect 29512 30200 29518 30252
rect 30837 30243 30895 30249
rect 30837 30209 30849 30243
rect 30883 30240 30895 30243
rect 30926 30240 30932 30252
rect 30883 30212 30932 30240
rect 30883 30209 30895 30212
rect 30837 30203 30895 30209
rect 30926 30200 30932 30212
rect 30984 30200 30990 30252
rect 31021 30243 31079 30249
rect 31021 30209 31033 30243
rect 31067 30240 31079 30243
rect 31386 30240 31392 30252
rect 31067 30212 31392 30240
rect 31067 30209 31079 30212
rect 31021 30203 31079 30209
rect 31386 30200 31392 30212
rect 31444 30200 31450 30252
rect 32030 30200 32036 30252
rect 32088 30240 32094 30252
rect 32125 30243 32183 30249
rect 32125 30240 32137 30243
rect 32088 30212 32137 30240
rect 32088 30200 32094 30212
rect 32125 30209 32137 30212
rect 32171 30240 32183 30243
rect 32766 30240 32772 30252
rect 32171 30212 32772 30240
rect 32171 30209 32183 30212
rect 32125 30203 32183 30209
rect 32766 30200 32772 30212
rect 32824 30200 32830 30252
rect 33410 30240 33416 30252
rect 33371 30212 33416 30240
rect 33410 30200 33416 30212
rect 33468 30200 33474 30252
rect 33502 30200 33508 30252
rect 33560 30240 33566 30252
rect 33612 30249 33640 30280
rect 34149 30277 34161 30311
rect 34195 30308 34207 30311
rect 34514 30308 34520 30320
rect 34195 30280 34520 30308
rect 34195 30277 34207 30280
rect 34149 30271 34207 30277
rect 34514 30268 34520 30280
rect 34572 30268 34578 30320
rect 34793 30311 34851 30317
rect 34793 30277 34805 30311
rect 34839 30308 34851 30311
rect 35986 30308 35992 30320
rect 34839 30280 35992 30308
rect 34839 30277 34851 30280
rect 34793 30271 34851 30277
rect 35986 30268 35992 30280
rect 36044 30268 36050 30320
rect 33597 30243 33655 30249
rect 33597 30240 33609 30243
rect 33560 30212 33609 30240
rect 33560 30200 33566 30212
rect 33597 30209 33609 30212
rect 33643 30209 33655 30243
rect 33597 30203 33655 30209
rect 33686 30200 33692 30252
rect 33744 30240 33750 30252
rect 33962 30240 33968 30252
rect 33744 30212 33789 30240
rect 33923 30212 33968 30240
rect 33744 30200 33750 30212
rect 33962 30200 33968 30212
rect 34020 30200 34026 30252
rect 34606 30200 34612 30252
rect 34664 30240 34670 30252
rect 34701 30243 34759 30249
rect 34701 30240 34713 30243
rect 34664 30212 34713 30240
rect 34664 30200 34670 30212
rect 34701 30209 34713 30212
rect 34747 30209 34759 30243
rect 34701 30203 34759 30209
rect 24044 30144 26096 30172
rect 27522 30132 27528 30184
rect 27580 30172 27586 30184
rect 28442 30172 28448 30184
rect 27580 30144 28448 30172
rect 27580 30132 27586 30144
rect 28442 30132 28448 30144
rect 28500 30132 28506 30184
rect 32398 30172 32404 30184
rect 32359 30144 32404 30172
rect 32398 30132 32404 30144
rect 32456 30132 32462 30184
rect 33781 30175 33839 30181
rect 33781 30141 33793 30175
rect 33827 30172 33839 30175
rect 34146 30172 34152 30184
rect 33827 30144 34152 30172
rect 33827 30141 33839 30144
rect 33781 30135 33839 30141
rect 34146 30132 34152 30144
rect 34204 30132 34210 30184
rect 46842 30172 46848 30184
rect 41386 30144 46848 30172
rect 41386 30104 41414 30144
rect 46842 30132 46848 30144
rect 46900 30132 46906 30184
rect 19260 30076 41414 30104
rect 14918 29996 14924 30048
rect 14976 30036 14982 30048
rect 15197 30039 15255 30045
rect 15197 30036 15209 30039
rect 14976 30008 15209 30036
rect 14976 29996 14982 30008
rect 15197 30005 15209 30008
rect 15243 30005 15255 30039
rect 19794 30036 19800 30048
rect 19755 30008 19800 30036
rect 15197 29999 15255 30005
rect 19794 29996 19800 30008
rect 19852 29996 19858 30048
rect 21266 30036 21272 30048
rect 21227 30008 21272 30036
rect 21266 29996 21272 30008
rect 21324 29996 21330 30048
rect 24210 30036 24216 30048
rect 24171 30008 24216 30036
rect 24210 29996 24216 30008
rect 24268 29996 24274 30048
rect 24486 29996 24492 30048
rect 24544 30036 24550 30048
rect 24857 30039 24915 30045
rect 24857 30036 24869 30039
rect 24544 30008 24869 30036
rect 24544 29996 24550 30008
rect 24857 30005 24869 30008
rect 24903 30005 24915 30039
rect 24857 29999 24915 30005
rect 26878 29996 26884 30048
rect 26936 30036 26942 30048
rect 27522 30036 27528 30048
rect 26936 30008 27528 30036
rect 26936 29996 26942 30008
rect 27522 29996 27528 30008
rect 27580 29996 27586 30048
rect 28350 30036 28356 30048
rect 28311 30008 28356 30036
rect 28350 29996 28356 30008
rect 28408 29996 28414 30048
rect 29178 29996 29184 30048
rect 29236 30036 29242 30048
rect 29362 30036 29368 30048
rect 29236 30008 29368 30036
rect 29236 29996 29242 30008
rect 29362 29996 29368 30008
rect 29420 29996 29426 30048
rect 30098 29996 30104 30048
rect 30156 30036 30162 30048
rect 30834 30036 30840 30048
rect 30156 30008 30840 30036
rect 30156 29996 30162 30008
rect 30834 29996 30840 30008
rect 30892 29996 30898 30048
rect 32030 29996 32036 30048
rect 32088 30036 32094 30048
rect 33042 30036 33048 30048
rect 32088 30008 33048 30036
rect 32088 29996 32094 30008
rect 33042 29996 33048 30008
rect 33100 29996 33106 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 27065 29835 27123 29841
rect 27065 29801 27077 29835
rect 27111 29832 27123 29835
rect 28074 29832 28080 29844
rect 27111 29804 28080 29832
rect 27111 29801 27123 29804
rect 27065 29795 27123 29801
rect 28074 29792 28080 29804
rect 28132 29792 28138 29844
rect 28626 29832 28632 29844
rect 28587 29804 28632 29832
rect 28626 29792 28632 29804
rect 28684 29792 28690 29844
rect 31573 29835 31631 29841
rect 31573 29801 31585 29835
rect 31619 29832 31631 29835
rect 32490 29832 32496 29844
rect 31619 29804 32496 29832
rect 31619 29801 31631 29804
rect 31573 29795 31631 29801
rect 32490 29792 32496 29804
rect 32548 29792 32554 29844
rect 32677 29835 32735 29841
rect 32677 29801 32689 29835
rect 32723 29832 32735 29835
rect 33410 29832 33416 29844
rect 32723 29804 33416 29832
rect 32723 29801 32735 29804
rect 32677 29795 32735 29801
rect 33410 29792 33416 29804
rect 33468 29792 33474 29844
rect 27249 29767 27307 29773
rect 27249 29733 27261 29767
rect 27295 29764 27307 29767
rect 27522 29764 27528 29776
rect 27295 29736 27528 29764
rect 27295 29733 27307 29736
rect 27249 29727 27307 29733
rect 27522 29724 27528 29736
rect 27580 29724 27586 29776
rect 30742 29764 30748 29776
rect 27632 29736 30748 29764
rect 14918 29696 14924 29708
rect 14879 29668 14924 29696
rect 14918 29656 14924 29668
rect 14976 29656 14982 29708
rect 16482 29696 16488 29708
rect 16443 29668 16488 29696
rect 16482 29656 16488 29668
rect 16540 29656 16546 29708
rect 19521 29699 19579 29705
rect 19521 29665 19533 29699
rect 19567 29696 19579 29699
rect 21266 29696 21272 29708
rect 19567 29668 21272 29696
rect 19567 29665 19579 29668
rect 19521 29659 19579 29665
rect 21266 29656 21272 29668
rect 21324 29656 21330 29708
rect 23750 29696 23756 29708
rect 23032 29668 23756 29696
rect 14090 29628 14096 29640
rect 14051 29600 14096 29628
rect 14090 29588 14096 29600
rect 14148 29588 14154 29640
rect 14734 29628 14740 29640
rect 14695 29600 14740 29628
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 19150 29588 19156 29640
rect 19208 29628 19214 29640
rect 23032 29637 23060 29668
rect 23750 29656 23756 29668
rect 23808 29656 23814 29708
rect 24762 29696 24768 29708
rect 24320 29668 24768 29696
rect 19245 29631 19303 29637
rect 19245 29628 19257 29631
rect 19208 29600 19257 29628
rect 19208 29588 19214 29600
rect 19245 29597 19257 29600
rect 19291 29597 19303 29631
rect 19245 29591 19303 29597
rect 23017 29631 23075 29637
rect 23017 29597 23029 29631
rect 23063 29597 23075 29631
rect 23198 29628 23204 29640
rect 23159 29600 23204 29628
rect 23017 29591 23075 29597
rect 23198 29588 23204 29600
rect 23256 29588 23262 29640
rect 23293 29631 23351 29637
rect 23293 29597 23305 29631
rect 23339 29597 23351 29631
rect 23293 29591 23351 29597
rect 19794 29520 19800 29572
rect 19852 29560 19858 29572
rect 23308 29560 23336 29591
rect 23382 29588 23388 29640
rect 23440 29628 23446 29640
rect 23569 29631 23627 29637
rect 23440 29600 23485 29628
rect 23440 29588 23446 29600
rect 23569 29597 23581 29631
rect 23615 29628 23627 29631
rect 23658 29628 23664 29640
rect 23615 29600 23664 29628
rect 23615 29597 23627 29600
rect 23569 29591 23627 29597
rect 23658 29588 23664 29600
rect 23716 29588 23722 29640
rect 24320 29560 24348 29668
rect 24762 29656 24768 29668
rect 24820 29656 24826 29708
rect 26050 29696 26056 29708
rect 24872 29668 26056 29696
rect 24486 29628 24492 29640
rect 24447 29600 24492 29628
rect 24486 29588 24492 29600
rect 24544 29588 24550 29640
rect 24637 29631 24695 29637
rect 24637 29597 24649 29631
rect 24683 29628 24695 29631
rect 24872 29628 24900 29668
rect 26050 29656 26056 29668
rect 26108 29656 26114 29708
rect 24683 29600 24900 29628
rect 24995 29631 25053 29637
rect 24683 29597 24695 29600
rect 24637 29591 24695 29597
rect 24995 29597 25007 29631
rect 25041 29628 25053 29631
rect 25222 29628 25228 29640
rect 25041 29600 25228 29628
rect 25041 29597 25053 29600
rect 24995 29591 25053 29597
rect 25222 29588 25228 29600
rect 25280 29588 25286 29640
rect 25590 29628 25596 29640
rect 25551 29600 25596 29628
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 27632 29628 27660 29736
rect 30742 29724 30748 29736
rect 30800 29724 30806 29776
rect 30926 29724 30932 29776
rect 30984 29764 30990 29776
rect 31757 29767 31815 29773
rect 31757 29764 31769 29767
rect 30984 29736 31769 29764
rect 30984 29724 30990 29736
rect 31757 29733 31769 29736
rect 31803 29733 31815 29767
rect 33870 29764 33876 29776
rect 31757 29727 31815 29733
rect 32416 29736 33876 29764
rect 27982 29656 27988 29708
rect 28040 29696 28046 29708
rect 30466 29696 30472 29708
rect 28040 29668 30472 29696
rect 28040 29656 28046 29668
rect 30466 29656 30472 29668
rect 30524 29656 30530 29708
rect 30834 29656 30840 29708
rect 30892 29696 30898 29708
rect 32309 29699 32367 29705
rect 32309 29696 32321 29699
rect 30892 29668 32321 29696
rect 30892 29656 30898 29668
rect 32309 29665 32321 29668
rect 32355 29665 32367 29699
rect 32309 29659 32367 29665
rect 25700 29600 27660 29628
rect 27803 29631 27861 29637
rect 24762 29560 24768 29572
rect 19852 29532 20010 29560
rect 23308 29532 24348 29560
rect 24723 29532 24768 29560
rect 19852 29520 19858 29532
rect 24762 29520 24768 29532
rect 24820 29520 24826 29572
rect 24857 29563 24915 29569
rect 24857 29529 24869 29563
rect 24903 29560 24915 29563
rect 25700 29560 25728 29600
rect 27803 29597 27815 29631
rect 27849 29626 27861 29631
rect 28074 29628 28080 29640
rect 27908 29626 28080 29628
rect 27849 29600 28080 29626
rect 27849 29598 27936 29600
rect 27849 29597 27861 29598
rect 27803 29591 27861 29597
rect 28074 29588 28080 29600
rect 28132 29588 28138 29640
rect 28166 29588 28172 29640
rect 28224 29628 28230 29640
rect 28445 29631 28503 29637
rect 28445 29628 28457 29631
rect 28224 29600 28457 29628
rect 28224 29588 28230 29600
rect 28445 29597 28457 29600
rect 28491 29597 28503 29631
rect 30558 29628 30564 29640
rect 30519 29600 30564 29628
rect 28445 29591 28503 29597
rect 30558 29588 30564 29600
rect 30616 29588 30622 29640
rect 31389 29631 31447 29637
rect 31389 29597 31401 29631
rect 31435 29628 31447 29631
rect 31478 29628 31484 29640
rect 31435 29600 31484 29628
rect 31435 29597 31447 29600
rect 31389 29591 31447 29597
rect 31478 29588 31484 29600
rect 31536 29588 31542 29640
rect 31573 29631 31631 29637
rect 31573 29597 31585 29631
rect 31619 29628 31631 29631
rect 32122 29628 32128 29640
rect 31619 29600 32128 29628
rect 31619 29597 31631 29600
rect 31573 29591 31631 29597
rect 32122 29588 32128 29600
rect 32180 29588 32186 29640
rect 32217 29631 32275 29637
rect 32217 29597 32229 29631
rect 32263 29628 32275 29631
rect 32416 29628 32444 29736
rect 33870 29724 33876 29736
rect 33928 29724 33934 29776
rect 32582 29696 32588 29708
rect 32543 29668 32588 29696
rect 32582 29656 32588 29668
rect 32640 29656 32646 29708
rect 33689 29699 33747 29705
rect 33689 29665 33701 29699
rect 33735 29696 33747 29699
rect 40218 29696 40224 29708
rect 33735 29668 40224 29696
rect 33735 29665 33747 29668
rect 33689 29659 33747 29665
rect 40218 29656 40224 29668
rect 40276 29656 40282 29708
rect 47210 29656 47216 29708
rect 47268 29696 47274 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 47268 29668 47593 29696
rect 47268 29656 47274 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 32263 29600 32444 29628
rect 32493 29631 32551 29637
rect 32263 29597 32275 29600
rect 32217 29591 32275 29597
rect 32493 29597 32505 29631
rect 32539 29628 32551 29631
rect 32539 29600 32628 29628
rect 32539 29597 32551 29600
rect 32493 29591 32551 29597
rect 24903 29532 25728 29560
rect 24903 29529 24915 29532
rect 24857 29523 24915 29529
rect 14185 29495 14243 29501
rect 14185 29461 14197 29495
rect 14231 29492 14243 29495
rect 14458 29492 14464 29504
rect 14231 29464 14464 29492
rect 14231 29461 14243 29464
rect 14185 29455 14243 29461
rect 14458 29452 14464 29464
rect 14516 29452 14522 29504
rect 20993 29495 21051 29501
rect 20993 29461 21005 29495
rect 21039 29492 21051 29495
rect 21174 29492 21180 29504
rect 21039 29464 21180 29492
rect 21039 29461 21051 29464
rect 20993 29455 21051 29461
rect 21174 29452 21180 29464
rect 21232 29452 21238 29504
rect 23566 29452 23572 29504
rect 23624 29492 23630 29504
rect 23753 29495 23811 29501
rect 23753 29492 23765 29495
rect 23624 29464 23765 29492
rect 23624 29452 23630 29464
rect 23753 29461 23765 29464
rect 23799 29461 23811 29495
rect 23753 29455 23811 29461
rect 23842 29452 23848 29504
rect 23900 29492 23906 29504
rect 24872 29492 24900 29523
rect 26694 29520 26700 29572
rect 26752 29560 26758 29572
rect 26881 29563 26939 29569
rect 26881 29560 26893 29563
rect 26752 29532 26893 29560
rect 26752 29520 26758 29532
rect 26881 29529 26893 29532
rect 26927 29529 26939 29563
rect 26881 29523 26939 29529
rect 27430 29520 27436 29572
rect 27488 29560 27494 29572
rect 29270 29560 29276 29572
rect 27488 29532 29276 29560
rect 27488 29520 27494 29532
rect 29270 29520 29276 29532
rect 29328 29520 29334 29572
rect 30745 29563 30803 29569
rect 30745 29529 30757 29563
rect 30791 29560 30803 29563
rect 32030 29560 32036 29572
rect 30791 29532 32036 29560
rect 30791 29529 30803 29532
rect 30745 29523 30803 29529
rect 32030 29520 32036 29532
rect 32088 29520 32094 29572
rect 32600 29560 32628 29600
rect 32950 29588 32956 29640
rect 33008 29628 33014 29640
rect 33321 29631 33379 29637
rect 33321 29628 33333 29631
rect 33008 29600 33333 29628
rect 33008 29588 33014 29600
rect 33321 29597 33333 29600
rect 33367 29597 33379 29631
rect 33502 29628 33508 29640
rect 33463 29600 33508 29628
rect 33321 29591 33379 29597
rect 33502 29588 33508 29600
rect 33560 29588 33566 29640
rect 33594 29588 33600 29640
rect 33652 29628 33658 29640
rect 33870 29628 33876 29640
rect 33652 29600 33697 29628
rect 33831 29600 33876 29628
rect 33652 29588 33658 29600
rect 33870 29588 33876 29600
rect 33928 29588 33934 29640
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 32508 29532 32628 29560
rect 32508 29504 32536 29532
rect 23900 29464 24900 29492
rect 23900 29452 23906 29464
rect 24946 29452 24952 29504
rect 25004 29492 25010 29504
rect 25133 29495 25191 29501
rect 25133 29492 25145 29495
rect 25004 29464 25145 29492
rect 25004 29452 25010 29464
rect 25133 29461 25145 29464
rect 25179 29461 25191 29495
rect 25682 29492 25688 29504
rect 25643 29464 25688 29492
rect 25133 29455 25191 29461
rect 25682 29452 25688 29464
rect 25740 29452 25746 29504
rect 26234 29452 26240 29504
rect 26292 29492 26298 29504
rect 26970 29492 26976 29504
rect 26292 29464 26976 29492
rect 26292 29452 26298 29464
rect 26970 29452 26976 29464
rect 27028 29492 27034 29504
rect 27081 29495 27139 29501
rect 27081 29492 27093 29495
rect 27028 29464 27093 29492
rect 27028 29452 27034 29464
rect 27081 29461 27093 29464
rect 27127 29461 27139 29495
rect 27081 29455 27139 29461
rect 27246 29452 27252 29504
rect 27304 29492 27310 29504
rect 27893 29495 27951 29501
rect 27893 29492 27905 29495
rect 27304 29464 27905 29492
rect 27304 29452 27310 29464
rect 27893 29461 27905 29464
rect 27939 29461 27951 29495
rect 27893 29455 27951 29461
rect 31478 29452 31484 29504
rect 31536 29492 31542 29504
rect 32398 29492 32404 29504
rect 31536 29464 32404 29492
rect 31536 29452 31542 29464
rect 32398 29452 32404 29464
rect 32456 29452 32462 29504
rect 32490 29452 32496 29504
rect 32548 29452 32554 29504
rect 34057 29495 34115 29501
rect 34057 29461 34069 29495
rect 34103 29492 34115 29495
rect 34238 29492 34244 29504
rect 34103 29464 34244 29492
rect 34103 29461 34115 29464
rect 34057 29455 34115 29461
rect 34238 29452 34244 29464
rect 34296 29452 34302 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 10965 29291 11023 29297
rect 10965 29257 10977 29291
rect 11011 29257 11023 29291
rect 20346 29288 20352 29300
rect 10965 29251 11023 29257
rect 20088 29260 20352 29288
rect 10980 29220 11008 29251
rect 11793 29223 11851 29229
rect 11793 29220 11805 29223
rect 10980 29192 11805 29220
rect 11793 29189 11805 29192
rect 11839 29189 11851 29223
rect 11793 29183 11851 29189
rect 12434 29180 12440 29232
rect 12492 29180 12498 29232
rect 14458 29220 14464 29232
rect 14419 29192 14464 29220
rect 14458 29180 14464 29192
rect 14516 29180 14522 29232
rect 10597 29155 10655 29161
rect 10597 29121 10609 29155
rect 10643 29152 10655 29155
rect 11054 29152 11060 29164
rect 10643 29124 11060 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 11054 29112 11060 29124
rect 11112 29112 11118 29164
rect 18506 29112 18512 29164
rect 18564 29152 18570 29164
rect 19153 29155 19211 29161
rect 19153 29152 19165 29155
rect 18564 29124 19165 29152
rect 18564 29112 18570 29124
rect 19153 29121 19165 29124
rect 19199 29152 19211 29155
rect 19334 29152 19340 29164
rect 19199 29124 19340 29152
rect 19199 29121 19211 29124
rect 19153 29115 19211 29121
rect 19334 29112 19340 29124
rect 19392 29112 19398 29164
rect 20088 29161 20116 29260
rect 20346 29248 20352 29260
rect 20404 29248 20410 29300
rect 20990 29248 20996 29300
rect 21048 29288 21054 29300
rect 21913 29291 21971 29297
rect 21913 29288 21925 29291
rect 21048 29260 21925 29288
rect 21048 29248 21054 29260
rect 21913 29257 21925 29260
rect 21959 29257 21971 29291
rect 21913 29251 21971 29257
rect 24854 29248 24860 29300
rect 24912 29288 24918 29300
rect 25041 29291 25099 29297
rect 25041 29288 25053 29291
rect 24912 29260 25053 29288
rect 24912 29248 24918 29260
rect 25041 29257 25053 29260
rect 25087 29257 25099 29291
rect 27706 29288 27712 29300
rect 27667 29260 27712 29288
rect 25041 29251 25099 29257
rect 27706 29248 27712 29260
rect 27764 29248 27770 29300
rect 28074 29248 28080 29300
rect 28132 29288 28138 29300
rect 28353 29291 28411 29297
rect 28353 29288 28365 29291
rect 28132 29260 28365 29288
rect 28132 29248 28138 29260
rect 28353 29257 28365 29260
rect 28399 29257 28411 29291
rect 28353 29251 28411 29257
rect 30285 29291 30343 29297
rect 30285 29257 30297 29291
rect 30331 29288 30343 29291
rect 30742 29288 30748 29300
rect 30331 29260 30748 29288
rect 30331 29257 30343 29260
rect 30285 29251 30343 29257
rect 30742 29248 30748 29260
rect 30800 29248 30806 29300
rect 31570 29288 31576 29300
rect 31531 29260 31576 29288
rect 31570 29248 31576 29260
rect 31628 29248 31634 29300
rect 31754 29248 31760 29300
rect 31812 29288 31818 29300
rect 32490 29288 32496 29300
rect 31812 29260 32496 29288
rect 31812 29248 31818 29260
rect 32490 29248 32496 29260
rect 32548 29248 32554 29300
rect 32950 29288 32956 29300
rect 32911 29260 32956 29288
rect 32950 29248 32956 29260
rect 33008 29248 33014 29300
rect 33594 29248 33600 29300
rect 33652 29288 33658 29300
rect 33778 29288 33784 29300
rect 33652 29260 33784 29288
rect 33652 29248 33658 29260
rect 33778 29248 33784 29260
rect 33836 29288 33842 29300
rect 35713 29291 35771 29297
rect 35713 29288 35725 29291
rect 33836 29260 35725 29288
rect 33836 29248 33842 29260
rect 35713 29257 35725 29260
rect 35759 29257 35771 29291
rect 35713 29251 35771 29257
rect 20165 29223 20223 29229
rect 20165 29189 20177 29223
rect 20211 29220 20223 29223
rect 23566 29220 23572 29232
rect 20211 29192 21864 29220
rect 23527 29192 23572 29220
rect 20211 29189 20223 29192
rect 20165 29183 20223 29189
rect 20073 29155 20131 29161
rect 20073 29121 20085 29155
rect 20119 29121 20131 29155
rect 20073 29115 20131 29121
rect 20257 29155 20315 29161
rect 20257 29121 20269 29155
rect 20303 29121 20315 29155
rect 20898 29152 20904 29164
rect 20859 29124 20904 29152
rect 20257 29115 20315 29121
rect 10686 29084 10692 29096
rect 10647 29056 10692 29084
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 11514 29084 11520 29096
rect 11475 29056 11520 29084
rect 11514 29044 11520 29056
rect 11572 29044 11578 29096
rect 14277 29087 14335 29093
rect 11624 29056 14228 29084
rect 8294 28976 8300 29028
rect 8352 29016 8358 29028
rect 11624 29016 11652 29056
rect 8352 28988 11652 29016
rect 13265 29019 13323 29025
rect 8352 28976 8358 28988
rect 13265 28985 13277 29019
rect 13311 28985 13323 29019
rect 14200 29016 14228 29056
rect 14277 29053 14289 29087
rect 14323 29084 14335 29087
rect 14458 29084 14464 29096
rect 14323 29056 14464 29084
rect 14323 29053 14335 29056
rect 14277 29047 14335 29053
rect 14458 29044 14464 29056
rect 14516 29044 14522 29096
rect 14737 29087 14795 29093
rect 14737 29053 14749 29087
rect 14783 29053 14795 29087
rect 14737 29047 14795 29053
rect 14752 29016 14780 29047
rect 14826 29044 14832 29096
rect 14884 29084 14890 29096
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 14884 29056 16681 29084
rect 14884 29044 14890 29056
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 16850 29084 16856 29096
rect 16811 29056 16856 29084
rect 16669 29047 16727 29053
rect 16850 29044 16856 29056
rect 16908 29044 16914 29096
rect 17129 29087 17187 29093
rect 17129 29053 17141 29087
rect 17175 29053 17187 29087
rect 17129 29047 17187 29053
rect 19245 29087 19303 29093
rect 19245 29053 19257 29087
rect 19291 29084 19303 29087
rect 19978 29084 19984 29096
rect 19291 29056 19984 29084
rect 19291 29053 19303 29056
rect 19245 29047 19303 29053
rect 14200 28988 14780 29016
rect 13265 28979 13323 28985
rect 11054 28908 11060 28960
rect 11112 28948 11118 28960
rect 12158 28948 12164 28960
rect 11112 28920 12164 28948
rect 11112 28908 11118 28920
rect 12158 28908 12164 28920
rect 12216 28948 12222 28960
rect 13280 28948 13308 28979
rect 16758 28976 16764 29028
rect 16816 29016 16822 29028
rect 17144 29016 17172 29047
rect 19978 29044 19984 29056
rect 20036 29044 20042 29096
rect 20272 29084 20300 29115
rect 20898 29112 20904 29124
rect 20956 29112 20962 29164
rect 21082 29152 21088 29164
rect 21043 29124 21088 29152
rect 21082 29112 21088 29124
rect 21140 29152 21146 29164
rect 21726 29152 21732 29164
rect 21140 29124 21732 29152
rect 21140 29112 21146 29124
rect 21726 29112 21732 29124
rect 21784 29112 21790 29164
rect 21836 29161 21864 29192
rect 23566 29180 23572 29192
rect 23624 29180 23630 29232
rect 25682 29220 25688 29232
rect 24794 29192 25688 29220
rect 25682 29180 25688 29192
rect 25740 29180 25746 29232
rect 27430 29180 27436 29232
rect 27488 29220 27494 29232
rect 31205 29223 31263 29229
rect 27488 29192 28304 29220
rect 27488 29180 27502 29192
rect 21821 29155 21879 29161
rect 21821 29121 21833 29155
rect 21867 29121 21879 29155
rect 22005 29155 22063 29161
rect 22005 29152 22017 29155
rect 21821 29115 21879 29121
rect 21928 29124 22017 29152
rect 20806 29084 20812 29096
rect 20272 29056 20812 29084
rect 20806 29044 20812 29056
rect 20864 29044 20870 29096
rect 21174 29084 21180 29096
rect 21135 29056 21180 29084
rect 21174 29044 21180 29056
rect 21232 29044 21238 29096
rect 21744 29084 21772 29112
rect 21928 29084 21956 29124
rect 22005 29121 22017 29124
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 25590 29112 25596 29164
rect 25648 29152 25654 29164
rect 25869 29155 25927 29161
rect 25869 29152 25881 29155
rect 25648 29124 25881 29152
rect 25648 29112 25654 29124
rect 25869 29121 25881 29124
rect 25915 29121 25927 29155
rect 25869 29115 25927 29121
rect 27474 29142 27502 29180
rect 27798 29152 27804 29164
rect 27474 29127 27568 29142
rect 27474 29121 27583 29127
rect 27759 29124 27804 29152
rect 27474 29114 27537 29121
rect 21744 29056 21956 29084
rect 23293 29087 23351 29093
rect 23293 29053 23305 29087
rect 23339 29084 23351 29087
rect 23339 29056 23373 29084
rect 23339 29053 23351 29056
rect 23293 29047 23351 29053
rect 16816 28988 17172 29016
rect 16816 28976 16822 28988
rect 19150 28976 19156 29028
rect 19208 29016 19214 29028
rect 23308 29016 23336 29047
rect 23658 29044 23664 29096
rect 23716 29084 23722 29096
rect 27525 29087 27537 29114
rect 27571 29087 27583 29121
rect 27798 29112 27804 29124
rect 27856 29112 27862 29164
rect 28276 29161 28304 29192
rect 31205 29189 31217 29223
rect 31251 29220 31263 29223
rect 34238 29220 34244 29232
rect 31251 29192 31616 29220
rect 34199 29192 34244 29220
rect 31251 29189 31263 29192
rect 31205 29183 31263 29189
rect 28261 29155 28319 29161
rect 28261 29121 28273 29155
rect 28307 29121 28319 29155
rect 28261 29115 28319 29121
rect 28350 29112 28356 29164
rect 28408 29152 28414 29164
rect 29457 29155 29515 29161
rect 29457 29152 29469 29155
rect 28408 29124 29469 29152
rect 28408 29112 28414 29124
rect 29457 29121 29469 29124
rect 29503 29152 29515 29155
rect 30006 29152 30012 29164
rect 29503 29124 30012 29152
rect 29503 29121 29515 29124
rect 29457 29115 29515 29121
rect 30006 29112 30012 29124
rect 30064 29112 30070 29164
rect 30101 29155 30159 29161
rect 30101 29121 30113 29155
rect 30147 29152 30159 29155
rect 30742 29152 30748 29164
rect 30147 29124 30748 29152
rect 30147 29121 30159 29124
rect 30101 29115 30159 29121
rect 30742 29112 30748 29124
rect 30800 29112 30806 29164
rect 31386 29152 31392 29164
rect 31347 29124 31392 29152
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 31588 29150 31616 29192
rect 34238 29180 34244 29192
rect 34296 29180 34302 29232
rect 34790 29180 34796 29232
rect 34848 29180 34854 29232
rect 32122 29152 32128 29164
rect 31772 29150 32128 29152
rect 31588 29124 32128 29150
rect 31588 29122 31800 29124
rect 32122 29112 32128 29124
rect 32180 29112 32186 29164
rect 32398 29152 32404 29164
rect 32359 29124 32404 29152
rect 32398 29112 32404 29124
rect 32456 29112 32462 29164
rect 33042 29112 33048 29164
rect 33100 29152 33106 29164
rect 33965 29155 34023 29161
rect 33965 29152 33977 29155
rect 33100 29124 33977 29152
rect 33100 29112 33106 29124
rect 33965 29121 33977 29124
rect 34011 29121 34023 29155
rect 33965 29115 34023 29121
rect 23716 29056 24624 29084
rect 27525 29081 27583 29087
rect 29730 29084 29736 29096
rect 23716 29044 23722 29056
rect 24596 29016 24624 29056
rect 27908 29056 29736 29084
rect 27341 29019 27399 29025
rect 19208 28988 23428 29016
rect 24596 28988 27292 29016
rect 19208 28976 19214 28988
rect 14826 28948 14832 28960
rect 12216 28920 14832 28948
rect 12216 28908 12222 28920
rect 14826 28908 14832 28920
rect 14884 28908 14890 28960
rect 20714 28948 20720 28960
rect 20675 28920 20720 28948
rect 20714 28908 20720 28920
rect 20772 28908 20778 28960
rect 23400 28948 23428 28988
rect 24210 28948 24216 28960
rect 23400 28920 24216 28948
rect 24210 28908 24216 28920
rect 24268 28948 24274 28960
rect 24670 28948 24676 28960
rect 24268 28920 24676 28948
rect 24268 28908 24274 28920
rect 24670 28908 24676 28920
rect 24728 28908 24734 28960
rect 25958 28948 25964 28960
rect 25919 28920 25964 28948
rect 25958 28908 25964 28920
rect 26016 28908 26022 28960
rect 27264 28948 27292 28988
rect 27341 28985 27353 29019
rect 27387 29016 27399 29019
rect 27614 29016 27620 29028
rect 27387 28988 27620 29016
rect 27387 28985 27399 28988
rect 27341 28979 27399 28985
rect 27614 28976 27620 28988
rect 27672 28976 27678 29028
rect 27908 29016 27936 29056
rect 29730 29044 29736 29056
rect 29788 29044 29794 29096
rect 32677 29087 32735 29093
rect 32677 29084 32689 29087
rect 31772 29056 32689 29084
rect 27724 28988 27936 29016
rect 31772 28994 31800 29056
rect 32677 29053 32689 29056
rect 32723 29053 32735 29087
rect 32677 29047 32735 29053
rect 27724 28948 27752 28988
rect 31680 28966 31800 28994
rect 29546 28948 29552 28960
rect 27264 28920 27752 28948
rect 29507 28920 29552 28948
rect 29546 28908 29552 28920
rect 29604 28908 29610 28960
rect 29638 28908 29644 28960
rect 29696 28948 29702 28960
rect 31680 28948 31708 28966
rect 29696 28920 31708 28948
rect 32769 28951 32827 28957
rect 29696 28908 29702 28920
rect 32769 28917 32781 28951
rect 32815 28948 32827 28951
rect 33502 28948 33508 28960
rect 32815 28920 33508 28948
rect 32815 28917 32827 28920
rect 32769 28911 32827 28917
rect 33502 28908 33508 28920
rect 33560 28908 33566 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 10686 28744 10692 28756
rect 10647 28716 10692 28744
rect 10686 28704 10692 28716
rect 10744 28704 10750 28756
rect 12434 28704 12440 28756
rect 12492 28744 12498 28756
rect 12492 28716 12537 28744
rect 12492 28704 12498 28716
rect 14458 28704 14464 28756
rect 14516 28744 14522 28756
rect 15841 28747 15899 28753
rect 15841 28744 15853 28747
rect 14516 28716 15853 28744
rect 14516 28704 14522 28716
rect 15841 28713 15853 28716
rect 15887 28713 15899 28747
rect 15841 28707 15899 28713
rect 16393 28747 16451 28753
rect 16393 28713 16405 28747
rect 16439 28744 16451 28747
rect 16850 28744 16856 28756
rect 16439 28716 16856 28744
rect 16439 28713 16451 28716
rect 16393 28707 16451 28713
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 17405 28747 17463 28753
rect 17405 28713 17417 28747
rect 17451 28744 17463 28747
rect 17586 28744 17592 28756
rect 17451 28716 17592 28744
rect 17451 28713 17463 28716
rect 17405 28707 17463 28713
rect 17586 28704 17592 28716
rect 17644 28704 17650 28756
rect 20714 28704 20720 28756
rect 20772 28744 20778 28756
rect 21545 28747 21603 28753
rect 21545 28744 21557 28747
rect 20772 28716 21557 28744
rect 20772 28704 20778 28716
rect 21545 28713 21557 28716
rect 21591 28713 21603 28747
rect 21545 28707 21603 28713
rect 21726 28704 21732 28756
rect 21784 28744 21790 28756
rect 22833 28747 22891 28753
rect 22833 28744 22845 28747
rect 21784 28716 22845 28744
rect 21784 28704 21790 28716
rect 22833 28713 22845 28716
rect 22879 28713 22891 28747
rect 22833 28707 22891 28713
rect 23106 28704 23112 28756
rect 23164 28744 23170 28756
rect 23164 28716 26004 28744
rect 23164 28704 23170 28716
rect 10045 28679 10103 28685
rect 10045 28645 10057 28679
rect 10091 28676 10103 28679
rect 11514 28676 11520 28688
rect 10091 28648 11520 28676
rect 10091 28645 10103 28648
rect 10045 28639 10103 28645
rect 11514 28636 11520 28648
rect 11572 28636 11578 28688
rect 20806 28636 20812 28688
rect 20864 28676 20870 28688
rect 20993 28679 21051 28685
rect 20993 28676 21005 28679
rect 20864 28648 21005 28676
rect 20864 28636 20870 28648
rect 20993 28645 21005 28648
rect 21039 28676 21051 28679
rect 21266 28676 21272 28688
rect 21039 28648 21272 28676
rect 21039 28645 21051 28648
rect 20993 28639 21051 28645
rect 21266 28636 21272 28648
rect 21324 28676 21330 28688
rect 25976 28676 26004 28716
rect 26050 28704 26056 28756
rect 26108 28744 26114 28756
rect 26421 28747 26479 28753
rect 26421 28744 26433 28747
rect 26108 28716 26433 28744
rect 26108 28704 26114 28716
rect 26421 28713 26433 28716
rect 26467 28713 26479 28747
rect 26421 28707 26479 28713
rect 26970 28704 26976 28756
rect 27028 28744 27034 28756
rect 27065 28747 27123 28753
rect 27065 28744 27077 28747
rect 27028 28716 27077 28744
rect 27028 28704 27034 28716
rect 27065 28713 27077 28716
rect 27111 28713 27123 28747
rect 27065 28707 27123 28713
rect 27614 28704 27620 28756
rect 27672 28744 27678 28756
rect 28902 28744 28908 28756
rect 27672 28716 28908 28744
rect 27672 28704 27678 28716
rect 28902 28704 28908 28716
rect 28960 28744 28966 28756
rect 30101 28747 30159 28753
rect 30101 28744 30113 28747
rect 28960 28716 30113 28744
rect 28960 28704 28966 28716
rect 30101 28713 30113 28716
rect 30147 28713 30159 28747
rect 30101 28707 30159 28713
rect 31938 28704 31944 28756
rect 31996 28744 32002 28756
rect 32125 28747 32183 28753
rect 32125 28744 32137 28747
rect 31996 28716 32137 28744
rect 31996 28704 32002 28716
rect 32125 28713 32137 28716
rect 32171 28713 32183 28747
rect 32125 28707 32183 28713
rect 32398 28704 32404 28756
rect 32456 28744 32462 28756
rect 32769 28747 32827 28753
rect 32769 28744 32781 28747
rect 32456 28716 32781 28744
rect 32456 28704 32462 28716
rect 32769 28713 32781 28716
rect 32815 28713 32827 28747
rect 34790 28744 34796 28756
rect 34751 28716 34796 28744
rect 32769 28707 32827 28713
rect 34790 28704 34796 28716
rect 34848 28704 34854 28756
rect 27801 28679 27859 28685
rect 27801 28676 27813 28679
rect 21324 28648 22692 28676
rect 25976 28648 27813 28676
rect 21324 28636 21330 28648
rect 11790 28608 11796 28620
rect 10796 28580 11796 28608
rect 9950 28540 9956 28552
rect 9911 28512 9956 28540
rect 9950 28500 9956 28512
rect 10008 28500 10014 28552
rect 10796 28549 10824 28580
rect 11790 28568 11796 28580
rect 11848 28568 11854 28620
rect 19150 28568 19156 28620
rect 19208 28608 19214 28620
rect 19245 28611 19303 28617
rect 19245 28608 19257 28611
rect 19208 28580 19257 28608
rect 19208 28568 19214 28580
rect 19245 28577 19257 28580
rect 19291 28577 19303 28611
rect 19245 28571 19303 28577
rect 19521 28611 19579 28617
rect 19521 28577 19533 28611
rect 19567 28608 19579 28611
rect 21358 28608 21364 28620
rect 19567 28580 21364 28608
rect 19567 28577 19579 28580
rect 19521 28571 19579 28577
rect 21358 28568 21364 28580
rect 21416 28568 21422 28620
rect 10597 28543 10655 28549
rect 10597 28509 10609 28543
rect 10643 28509 10655 28543
rect 10597 28503 10655 28509
rect 10781 28543 10839 28549
rect 10781 28509 10793 28543
rect 10827 28509 10839 28543
rect 11238 28540 11244 28552
rect 11199 28512 11244 28540
rect 10781 28503 10839 28509
rect 10612 28472 10640 28503
rect 11238 28500 11244 28512
rect 11296 28500 11302 28552
rect 11422 28540 11428 28552
rect 11383 28512 11428 28540
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 12342 28540 12348 28552
rect 12303 28512 12348 28540
rect 12342 28500 12348 28512
rect 12400 28500 12406 28552
rect 14090 28540 14096 28552
rect 14051 28512 14096 28540
rect 14090 28500 14096 28512
rect 14148 28500 14154 28552
rect 16301 28543 16359 28549
rect 16301 28509 16313 28543
rect 16347 28540 16359 28543
rect 16574 28540 16580 28552
rect 16347 28512 16580 28540
rect 16347 28509 16359 28512
rect 16301 28503 16359 28509
rect 16574 28500 16580 28512
rect 16632 28500 16638 28552
rect 17310 28540 17316 28552
rect 17223 28512 17316 28540
rect 17310 28500 17316 28512
rect 17368 28540 17374 28552
rect 17862 28540 17868 28552
rect 17368 28512 17868 28540
rect 17368 28500 17374 28512
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 18506 28540 18512 28552
rect 18467 28512 18512 28540
rect 18506 28500 18512 28512
rect 18564 28500 18570 28552
rect 21453 28543 21511 28549
rect 21453 28509 21465 28543
rect 21499 28540 21511 28543
rect 21726 28540 21732 28552
rect 21499 28512 21732 28540
rect 21499 28509 21511 28512
rect 21453 28503 21511 28509
rect 21726 28500 21732 28512
rect 21784 28500 21790 28552
rect 22664 28549 22692 28648
rect 27801 28645 27813 28648
rect 27847 28645 27859 28679
rect 27801 28639 27859 28645
rect 24946 28608 24952 28620
rect 24907 28580 24952 28608
rect 24946 28568 24952 28580
rect 25004 28568 25010 28620
rect 27816 28608 27844 28639
rect 28626 28636 28632 28688
rect 28684 28676 28690 28688
rect 29638 28676 29644 28688
rect 28684 28648 29644 28676
rect 28684 28636 28690 28648
rect 29638 28636 29644 28648
rect 29696 28636 29702 28688
rect 30653 28611 30711 28617
rect 27816 28580 29868 28608
rect 21821 28543 21879 28549
rect 21821 28509 21833 28543
rect 21867 28540 21879 28543
rect 22649 28543 22707 28549
rect 21867 28512 22600 28540
rect 21867 28509 21879 28512
rect 21821 28503 21879 28509
rect 11974 28472 11980 28484
rect 10612 28444 11980 28472
rect 11974 28432 11980 28444
rect 12032 28432 12038 28484
rect 13170 28432 13176 28484
rect 13228 28472 13234 28484
rect 14369 28475 14427 28481
rect 14369 28472 14381 28475
rect 13228 28444 14381 28472
rect 13228 28432 13234 28444
rect 14369 28441 14381 28444
rect 14415 28441 14427 28475
rect 14369 28435 14427 28441
rect 15378 28432 15384 28484
rect 15436 28432 15442 28484
rect 19978 28432 19984 28484
rect 20036 28432 20042 28484
rect 22094 28472 22100 28484
rect 21744 28444 22100 28472
rect 11330 28404 11336 28416
rect 11291 28376 11336 28404
rect 11330 28364 11336 28376
rect 11388 28364 11394 28416
rect 11790 28364 11796 28416
rect 11848 28404 11854 28416
rect 14734 28404 14740 28416
rect 11848 28376 14740 28404
rect 11848 28364 11854 28376
rect 14734 28364 14740 28376
rect 14792 28364 14798 28416
rect 18601 28407 18659 28413
rect 18601 28373 18613 28407
rect 18647 28404 18659 28407
rect 19334 28404 19340 28416
rect 18647 28376 19340 28404
rect 18647 28373 18659 28376
rect 18601 28367 18659 28373
rect 19334 28364 19340 28376
rect 19392 28364 19398 28416
rect 20346 28364 20352 28416
rect 20404 28404 20410 28416
rect 21744 28404 21772 28444
rect 22094 28432 22100 28444
rect 22152 28472 22158 28484
rect 22465 28475 22523 28481
rect 22465 28472 22477 28475
rect 22152 28444 22477 28472
rect 22152 28432 22158 28444
rect 22465 28441 22477 28444
rect 22511 28441 22523 28475
rect 22572 28472 22600 28512
rect 22649 28509 22661 28543
rect 22695 28509 22707 28543
rect 22649 28503 22707 28509
rect 23014 28500 23020 28552
rect 23072 28540 23078 28552
rect 23293 28543 23351 28549
rect 23293 28540 23305 28543
rect 23072 28512 23305 28540
rect 23072 28500 23078 28512
rect 23293 28509 23305 28512
rect 23339 28509 23351 28543
rect 24670 28540 24676 28552
rect 24631 28512 24676 28540
rect 23293 28503 23351 28509
rect 24670 28500 24676 28512
rect 24728 28500 24734 28552
rect 27062 28500 27068 28552
rect 27120 28540 27126 28552
rect 27522 28540 27528 28552
rect 27120 28512 27528 28540
rect 27120 28500 27126 28512
rect 27522 28500 27528 28512
rect 27580 28540 27586 28552
rect 29840 28549 29868 28580
rect 30653 28577 30665 28611
rect 30699 28608 30711 28611
rect 31386 28608 31392 28620
rect 30699 28580 31392 28608
rect 30699 28577 30711 28580
rect 30653 28571 30711 28577
rect 27617 28543 27675 28549
rect 27617 28540 27629 28543
rect 27580 28512 27629 28540
rect 27580 28500 27586 28512
rect 27617 28509 27629 28512
rect 27663 28540 27675 28543
rect 28445 28543 28503 28549
rect 28445 28540 28457 28543
rect 27663 28512 28457 28540
rect 27663 28509 27675 28512
rect 27617 28503 27675 28509
rect 28445 28509 28457 28512
rect 28491 28509 28503 28543
rect 28445 28503 28503 28509
rect 29825 28543 29883 28549
rect 29825 28509 29837 28543
rect 29871 28509 29883 28543
rect 29825 28503 29883 28509
rect 29977 28543 30035 28549
rect 29977 28509 29989 28543
rect 30023 28540 30035 28543
rect 30098 28540 30104 28552
rect 30023 28512 30104 28540
rect 30023 28509 30035 28512
rect 29977 28503 30035 28509
rect 23934 28472 23940 28484
rect 22572 28444 23940 28472
rect 22465 28435 22523 28441
rect 23934 28432 23940 28444
rect 23992 28432 23998 28484
rect 25958 28432 25964 28484
rect 26016 28432 26022 28484
rect 26970 28472 26976 28484
rect 26931 28444 26976 28472
rect 26970 28432 26976 28444
rect 27028 28432 27034 28484
rect 29840 28472 29868 28503
rect 30098 28500 30104 28512
rect 30156 28500 30162 28552
rect 30193 28543 30251 28549
rect 30193 28509 30205 28543
rect 30239 28540 30251 28543
rect 30374 28540 30380 28552
rect 30239 28512 30380 28540
rect 30239 28509 30251 28512
rect 30193 28503 30251 28509
rect 30374 28500 30380 28512
rect 30432 28540 30438 28552
rect 30668 28540 30696 28571
rect 31386 28568 31392 28580
rect 31444 28568 31450 28620
rect 32122 28568 32128 28620
rect 32180 28608 32186 28620
rect 32217 28611 32275 28617
rect 32217 28608 32229 28611
rect 32180 28580 32229 28608
rect 32180 28568 32186 28580
rect 32217 28577 32229 28580
rect 32263 28608 32275 28611
rect 32950 28608 32956 28620
rect 32263 28580 32956 28608
rect 32263 28577 32275 28580
rect 32217 28571 32275 28577
rect 32950 28568 32956 28580
rect 33008 28568 33014 28620
rect 30432 28512 30696 28540
rect 30837 28543 30895 28549
rect 30432 28500 30438 28512
rect 30837 28509 30849 28543
rect 30883 28540 30895 28543
rect 30926 28540 30932 28552
rect 30883 28512 30932 28540
rect 30883 28509 30895 28512
rect 30837 28503 30895 28509
rect 30926 28500 30932 28512
rect 30984 28500 30990 28552
rect 31662 28540 31668 28552
rect 31036 28512 31668 28540
rect 30650 28472 30656 28484
rect 29840 28444 30656 28472
rect 30650 28432 30656 28444
rect 30708 28472 30714 28484
rect 31036 28472 31064 28512
rect 31662 28500 31668 28512
rect 31720 28500 31726 28552
rect 31938 28540 31944 28552
rect 31899 28512 31944 28540
rect 31938 28500 31944 28512
rect 31996 28500 32002 28552
rect 32674 28540 32680 28552
rect 32635 28512 32680 28540
rect 32674 28500 32680 28512
rect 32732 28500 32738 28552
rect 34606 28500 34612 28552
rect 34664 28540 34670 28552
rect 34701 28543 34759 28549
rect 34701 28540 34713 28543
rect 34664 28512 34713 28540
rect 34664 28500 34670 28512
rect 34701 28509 34713 28512
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 46934 28500 46940 28552
rect 46992 28540 46998 28552
rect 47673 28543 47731 28549
rect 47673 28540 47685 28543
rect 46992 28512 47685 28540
rect 46992 28500 46998 28512
rect 47673 28509 47685 28512
rect 47719 28509 47731 28543
rect 47673 28503 47731 28509
rect 30708 28444 31064 28472
rect 30708 28432 30714 28444
rect 31570 28432 31576 28484
rect 31628 28472 31634 28484
rect 32953 28475 33011 28481
rect 32953 28472 32965 28475
rect 31628 28444 32965 28472
rect 31628 28432 31634 28444
rect 32953 28441 32965 28444
rect 32999 28441 33011 28475
rect 32953 28435 33011 28441
rect 20404 28376 21772 28404
rect 20404 28364 20410 28376
rect 21818 28364 21824 28416
rect 21876 28404 21882 28416
rect 22005 28407 22063 28413
rect 22005 28404 22017 28407
rect 21876 28376 22017 28404
rect 21876 28364 21882 28376
rect 22005 28373 22017 28376
rect 22051 28373 22063 28407
rect 22005 28367 22063 28373
rect 23382 28364 23388 28416
rect 23440 28404 23446 28416
rect 23477 28407 23535 28413
rect 23477 28404 23489 28407
rect 23440 28376 23489 28404
rect 23440 28364 23446 28376
rect 23477 28373 23489 28376
rect 23523 28373 23535 28407
rect 23952 28404 23980 28432
rect 28537 28407 28595 28413
rect 28537 28404 28549 28407
rect 23952 28376 28549 28404
rect 23477 28367 23535 28373
rect 28537 28373 28549 28376
rect 28583 28404 28595 28407
rect 28626 28404 28632 28416
rect 28583 28376 28632 28404
rect 28583 28373 28595 28376
rect 28537 28367 28595 28373
rect 28626 28364 28632 28376
rect 28684 28364 28690 28416
rect 29641 28407 29699 28413
rect 29641 28373 29653 28407
rect 29687 28404 29699 28407
rect 29822 28404 29828 28416
rect 29687 28376 29828 28404
rect 29687 28373 29699 28376
rect 29641 28367 29699 28373
rect 29822 28364 29828 28376
rect 29880 28364 29886 28416
rect 31018 28404 31024 28416
rect 30979 28376 31024 28404
rect 31018 28364 31024 28376
rect 31076 28364 31082 28416
rect 31757 28407 31815 28413
rect 31757 28373 31769 28407
rect 31803 28404 31815 28407
rect 32582 28404 32588 28416
rect 31803 28376 32588 28404
rect 31803 28373 31815 28376
rect 31757 28367 31815 28373
rect 32582 28364 32588 28376
rect 32640 28364 32646 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 3602 28160 3608 28212
rect 3660 28200 3666 28212
rect 11790 28200 11796 28212
rect 3660 28172 11376 28200
rect 11751 28172 11796 28200
rect 3660 28160 3666 28172
rect 3326 28024 3332 28076
rect 3384 28064 3390 28076
rect 3602 28064 3608 28076
rect 3384 28036 3608 28064
rect 3384 28024 3390 28036
rect 3602 28024 3608 28036
rect 3660 28024 3666 28076
rect 9950 28024 9956 28076
rect 10008 28064 10014 28076
rect 10321 28067 10379 28073
rect 10321 28064 10333 28067
rect 10008 28036 10333 28064
rect 10008 28024 10014 28036
rect 10321 28033 10333 28036
rect 10367 28033 10379 28067
rect 10321 28027 10379 28033
rect 10502 27860 10508 27872
rect 10463 27832 10508 27860
rect 10502 27820 10508 27832
rect 10560 27820 10566 27872
rect 11348 27860 11376 28172
rect 11790 28160 11796 28172
rect 11848 28160 11854 28212
rect 13170 28200 13176 28212
rect 13131 28172 13176 28200
rect 13170 28160 13176 28172
rect 13228 28160 13234 28212
rect 14458 28200 14464 28212
rect 14108 28172 14464 28200
rect 11701 28135 11759 28141
rect 11701 28101 11713 28135
rect 11747 28132 11759 28135
rect 12158 28132 12164 28144
rect 11747 28104 12164 28132
rect 11747 28101 11759 28104
rect 11701 28095 11759 28101
rect 12158 28092 12164 28104
rect 12216 28092 12222 28144
rect 13814 28132 13820 28144
rect 12544 28104 13820 28132
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 11974 28064 11980 28076
rect 11931 28036 11980 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 11974 28024 11980 28036
rect 12032 28024 12038 28076
rect 12342 28024 12348 28076
rect 12400 28064 12406 28076
rect 12544 28073 12572 28104
rect 13814 28092 13820 28104
rect 13872 28092 13878 28144
rect 14108 28141 14136 28172
rect 14458 28160 14464 28172
rect 14516 28160 14522 28212
rect 15197 28203 15255 28209
rect 15197 28169 15209 28203
rect 15243 28200 15255 28203
rect 15378 28200 15384 28212
rect 15243 28172 15384 28200
rect 15243 28169 15255 28172
rect 15197 28163 15255 28169
rect 15378 28160 15384 28172
rect 15436 28160 15442 28212
rect 16574 28200 16580 28212
rect 15948 28172 16580 28200
rect 14093 28135 14151 28141
rect 14093 28101 14105 28135
rect 14139 28101 14151 28135
rect 14093 28095 14151 28101
rect 14369 28135 14427 28141
rect 14369 28101 14381 28135
rect 14415 28132 14427 28135
rect 14826 28132 14832 28144
rect 14415 28104 14832 28132
rect 14415 28101 14427 28104
rect 14369 28095 14427 28101
rect 12529 28067 12587 28073
rect 12529 28064 12541 28067
rect 12400 28036 12541 28064
rect 12400 28024 12406 28036
rect 12529 28033 12541 28036
rect 12575 28033 12587 28067
rect 12529 28027 12587 28033
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28064 13415 28067
rect 13998 28064 14004 28076
rect 13403 28036 14004 28064
rect 13403 28033 13415 28036
rect 13357 28027 13415 28033
rect 13998 28024 14004 28036
rect 14056 28024 14062 28076
rect 11422 27956 11428 28008
rect 11480 27996 11486 28008
rect 12069 27999 12127 28005
rect 12069 27996 12081 27999
rect 11480 27968 12081 27996
rect 11480 27956 11486 27968
rect 12069 27965 12081 27968
rect 12115 27996 12127 27999
rect 13541 27999 13599 28005
rect 13541 27996 13553 27999
rect 12115 27968 13553 27996
rect 12115 27965 12127 27968
rect 12069 27959 12127 27965
rect 13541 27965 13553 27968
rect 13587 27965 13599 27999
rect 13541 27959 13599 27965
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27996 13691 27999
rect 14108 27996 14136 28095
rect 14826 28092 14832 28104
rect 14884 28092 14890 28144
rect 14274 28064 14280 28076
rect 14235 28036 14280 28064
rect 14274 28024 14280 28036
rect 14332 28024 14338 28076
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28064 14519 28067
rect 14734 28064 14740 28076
rect 14507 28036 14740 28064
rect 14507 28033 14519 28036
rect 14461 28027 14519 28033
rect 14734 28024 14740 28036
rect 14792 28024 14798 28076
rect 15102 28064 15108 28076
rect 15063 28036 15108 28064
rect 15102 28024 15108 28036
rect 15160 28024 15166 28076
rect 15948 28073 15976 28172
rect 16574 28160 16580 28172
rect 16632 28200 16638 28212
rect 17586 28200 17592 28212
rect 16632 28172 17592 28200
rect 16632 28160 16638 28172
rect 17586 28160 17592 28172
rect 17644 28160 17650 28212
rect 22557 28203 22615 28209
rect 22557 28200 22569 28203
rect 19260 28172 22569 28200
rect 16025 28135 16083 28141
rect 16025 28101 16037 28135
rect 16071 28132 16083 28135
rect 16853 28135 16911 28141
rect 16853 28132 16865 28135
rect 16071 28104 16865 28132
rect 16071 28101 16083 28104
rect 16025 28095 16083 28101
rect 16853 28101 16865 28104
rect 16899 28101 16911 28135
rect 19150 28132 19156 28144
rect 16853 28095 16911 28101
rect 18984 28104 19156 28132
rect 18984 28073 19012 28104
rect 19150 28092 19156 28104
rect 19208 28092 19214 28144
rect 19260 28141 19288 28172
rect 22557 28169 22569 28172
rect 22603 28169 22615 28203
rect 27522 28200 27528 28212
rect 27483 28172 27528 28200
rect 22557 28163 22615 28169
rect 27522 28160 27528 28172
rect 27580 28160 27586 28212
rect 32030 28200 32036 28212
rect 28552 28172 32036 28200
rect 19245 28135 19303 28141
rect 19245 28101 19257 28135
rect 19291 28101 19303 28135
rect 19245 28095 19303 28101
rect 19334 28092 19340 28144
rect 19392 28132 19398 28144
rect 19392 28104 19734 28132
rect 19392 28092 19398 28104
rect 21542 28092 21548 28144
rect 21600 28132 21606 28144
rect 21600 28104 22048 28132
rect 21600 28092 21606 28104
rect 22020 28076 22048 28104
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28033 15991 28067
rect 15933 28027 15991 28033
rect 18969 28067 19027 28073
rect 18969 28033 18981 28067
rect 19015 28033 19027 28067
rect 21818 28064 21824 28076
rect 21779 28036 21824 28064
rect 18969 28027 19027 28033
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 22002 28064 22008 28076
rect 21915 28036 22008 28064
rect 22002 28024 22008 28036
rect 22060 28024 22066 28076
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28064 22431 28067
rect 22830 28064 22836 28076
rect 22419 28036 22836 28064
rect 22419 28033 22431 28036
rect 22373 28027 22431 28033
rect 22830 28024 22836 28036
rect 22888 28064 22894 28076
rect 23382 28064 23388 28076
rect 22888 28036 23388 28064
rect 22888 28024 22894 28036
rect 23382 28024 23388 28036
rect 23440 28024 23446 28076
rect 25498 28024 25504 28076
rect 25556 28064 25562 28076
rect 26970 28064 26976 28076
rect 25556 28036 26976 28064
rect 25556 28024 25562 28036
rect 26970 28024 26976 28036
rect 27028 28024 27034 28076
rect 27062 28024 27068 28076
rect 27120 28064 27126 28076
rect 27341 28067 27399 28073
rect 27341 28064 27353 28067
rect 27120 28036 27353 28064
rect 27120 28024 27126 28036
rect 27341 28033 27353 28036
rect 27387 28064 27399 28067
rect 28258 28064 28264 28076
rect 27387 28036 28264 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 28258 28024 28264 28036
rect 28316 28024 28322 28076
rect 13679 27968 14136 27996
rect 13679 27965 13691 27968
rect 13633 27959 13691 27965
rect 16574 27956 16580 28008
rect 16632 27996 16638 28008
rect 16669 27999 16727 28005
rect 16669 27996 16681 27999
rect 16632 27968 16681 27996
rect 16632 27956 16638 27968
rect 16669 27965 16681 27968
rect 16715 27965 16727 27999
rect 16669 27959 16727 27965
rect 17129 27999 17187 28005
rect 17129 27965 17141 27999
rect 17175 27965 17187 27999
rect 20898 27996 20904 28008
rect 17129 27959 17187 27965
rect 20732 27968 20904 27996
rect 11514 27928 11520 27940
rect 11475 27900 11520 27928
rect 11514 27888 11520 27900
rect 11572 27888 11578 27940
rect 17144 27928 17172 27959
rect 11624 27900 14044 27928
rect 11624 27860 11652 27900
rect 12618 27860 12624 27872
rect 11348 27832 11652 27860
rect 12579 27832 12624 27860
rect 12618 27820 12624 27832
rect 12676 27820 12682 27872
rect 14016 27860 14044 27900
rect 14200 27900 17172 27928
rect 14200 27860 14228 27900
rect 20732 27872 20760 27968
rect 20898 27956 20904 27968
rect 20956 27996 20962 28008
rect 22097 27999 22155 28005
rect 22097 27996 22109 27999
rect 20956 27968 22109 27996
rect 20956 27956 20962 27968
rect 22097 27965 22109 27968
rect 22143 27965 22155 27999
rect 22097 27959 22155 27965
rect 22186 27956 22192 28008
rect 22244 27996 22250 28008
rect 22244 27968 22289 27996
rect 22244 27956 22250 27968
rect 28074 27956 28080 28008
rect 28132 27996 28138 28008
rect 28552 28005 28580 28172
rect 32030 28160 32036 28172
rect 32088 28160 32094 28212
rect 32950 28160 32956 28212
rect 33008 28200 33014 28212
rect 34057 28203 34115 28209
rect 34057 28200 34069 28203
rect 33008 28172 34069 28200
rect 33008 28160 33014 28172
rect 34057 28169 34069 28172
rect 34103 28169 34115 28203
rect 34057 28163 34115 28169
rect 29546 28092 29552 28144
rect 29604 28092 29610 28144
rect 30926 28092 30932 28144
rect 30984 28132 30990 28144
rect 31481 28135 31539 28141
rect 31481 28132 31493 28135
rect 30984 28104 31493 28132
rect 30984 28092 30990 28104
rect 31481 28101 31493 28104
rect 31527 28101 31539 28135
rect 31481 28095 31539 28101
rect 30834 28024 30840 28076
rect 30892 28064 30898 28076
rect 31297 28067 31355 28073
rect 31297 28064 31309 28067
rect 30892 28036 31309 28064
rect 30892 28024 30898 28036
rect 31297 28033 31309 28036
rect 31343 28033 31355 28067
rect 31297 28027 31355 28033
rect 31570 28024 31576 28076
rect 31628 28064 31634 28076
rect 32048 28064 32076 28160
rect 32582 28132 32588 28144
rect 32543 28104 32588 28132
rect 32582 28092 32588 28104
rect 32640 28092 32646 28144
rect 33594 28092 33600 28144
rect 33652 28092 33658 28144
rect 32306 28064 32312 28076
rect 31628 28036 31673 28064
rect 32048 28036 32312 28064
rect 31628 28024 31634 28036
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 45830 28024 45836 28076
rect 45888 28064 45894 28076
rect 47581 28067 47639 28073
rect 47581 28064 47593 28067
rect 45888 28036 47593 28064
rect 45888 28024 45894 28036
rect 47581 28033 47593 28036
rect 47627 28033 47639 28067
rect 47581 28027 47639 28033
rect 28537 27999 28595 28005
rect 28537 27996 28549 27999
rect 28132 27968 28549 27996
rect 28132 27956 28138 27968
rect 28537 27965 28549 27968
rect 28583 27965 28595 27999
rect 28537 27959 28595 27965
rect 28813 27999 28871 28005
rect 28813 27965 28825 27999
rect 28859 27996 28871 27999
rect 29546 27996 29552 28008
rect 28859 27968 29552 27996
rect 28859 27965 28871 27968
rect 28813 27959 28871 27965
rect 29546 27956 29552 27968
rect 29604 27956 29610 28008
rect 30285 27999 30343 28005
rect 30285 27965 30297 27999
rect 30331 27996 30343 27999
rect 30374 27996 30380 28008
rect 30331 27968 30380 27996
rect 30331 27965 30343 27968
rect 30285 27959 30343 27965
rect 30374 27956 30380 27968
rect 30432 27956 30438 28008
rect 14016 27832 14228 27860
rect 14645 27863 14703 27869
rect 14645 27829 14657 27863
rect 14691 27860 14703 27863
rect 14826 27860 14832 27872
rect 14691 27832 14832 27860
rect 14691 27829 14703 27832
rect 14645 27823 14703 27829
rect 14826 27820 14832 27832
rect 14884 27820 14890 27872
rect 20714 27860 20720 27872
rect 20675 27832 20720 27860
rect 20714 27820 20720 27832
rect 20772 27820 20778 27872
rect 27341 27863 27399 27869
rect 27341 27829 27353 27863
rect 27387 27860 27399 27863
rect 27430 27860 27436 27872
rect 27387 27832 27436 27860
rect 27387 27829 27399 27832
rect 27341 27823 27399 27829
rect 27430 27820 27436 27832
rect 27488 27820 27494 27872
rect 31297 27863 31355 27869
rect 31297 27829 31309 27863
rect 31343 27860 31355 27863
rect 32122 27860 32128 27872
rect 31343 27832 32128 27860
rect 31343 27829 31355 27832
rect 31297 27823 31355 27829
rect 32122 27820 32128 27832
rect 32180 27820 32186 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 10860 27659 10918 27665
rect 10860 27625 10872 27659
rect 10906 27656 10918 27659
rect 11330 27656 11336 27668
rect 10906 27628 11336 27656
rect 10906 27625 10918 27628
rect 10860 27619 10918 27625
rect 11330 27616 11336 27628
rect 11388 27616 11394 27668
rect 11514 27616 11520 27668
rect 11572 27656 11578 27668
rect 11882 27656 11888 27668
rect 11572 27628 11888 27656
rect 11572 27616 11578 27628
rect 11882 27616 11888 27628
rect 11940 27656 11946 27668
rect 12345 27659 12403 27665
rect 12345 27656 12357 27659
rect 11940 27628 12357 27656
rect 11940 27616 11946 27628
rect 12345 27625 12357 27628
rect 12391 27656 12403 27659
rect 14274 27656 14280 27668
rect 12391 27628 14280 27656
rect 12391 27625 12403 27628
rect 12345 27619 12403 27625
rect 14274 27616 14280 27628
rect 14332 27616 14338 27668
rect 31573 27659 31631 27665
rect 31573 27625 31585 27659
rect 31619 27656 31631 27659
rect 31938 27656 31944 27668
rect 31619 27628 31944 27656
rect 31619 27625 31631 27628
rect 31573 27619 31631 27625
rect 31938 27616 31944 27628
rect 31996 27616 32002 27668
rect 42518 27616 42524 27668
rect 42576 27656 42582 27668
rect 46198 27656 46204 27668
rect 42576 27628 46204 27656
rect 42576 27616 42582 27628
rect 46198 27616 46204 27628
rect 46256 27616 46262 27668
rect 7466 27548 7472 27600
rect 7524 27588 7530 27600
rect 13449 27591 13507 27597
rect 7524 27560 10732 27588
rect 7524 27548 7530 27560
rect 10502 27480 10508 27532
rect 10560 27520 10566 27532
rect 10597 27523 10655 27529
rect 10597 27520 10609 27523
rect 10560 27492 10609 27520
rect 10560 27480 10566 27492
rect 10597 27489 10609 27492
rect 10643 27489 10655 27523
rect 10704 27520 10732 27560
rect 13449 27557 13461 27591
rect 13495 27588 13507 27591
rect 14090 27588 14096 27600
rect 13495 27560 14096 27588
rect 13495 27557 13507 27560
rect 13449 27551 13507 27557
rect 14090 27548 14096 27560
rect 14148 27548 14154 27600
rect 21358 27548 21364 27600
rect 21416 27588 21422 27600
rect 21453 27591 21511 27597
rect 21453 27588 21465 27591
rect 21416 27560 21465 27588
rect 21416 27548 21422 27560
rect 21453 27557 21465 27560
rect 21499 27557 21511 27591
rect 21453 27551 21511 27557
rect 23014 27548 23020 27600
rect 23072 27588 23078 27600
rect 26510 27588 26516 27600
rect 23072 27560 26516 27588
rect 23072 27548 23078 27560
rect 26510 27548 26516 27560
rect 26568 27548 26574 27600
rect 29546 27588 29552 27600
rect 29507 27560 29552 27588
rect 29546 27548 29552 27560
rect 29604 27548 29610 27600
rect 31018 27588 31024 27600
rect 29748 27560 31024 27588
rect 23201 27523 23259 27529
rect 23201 27520 23213 27523
rect 10704 27492 23213 27520
rect 10597 27483 10655 27489
rect 23201 27489 23213 27492
rect 23247 27489 23259 27523
rect 23201 27483 23259 27489
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 13906 27452 13912 27464
rect 13403 27424 13912 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 13906 27412 13912 27424
rect 13964 27412 13970 27464
rect 14090 27412 14096 27464
rect 14148 27452 14154 27464
rect 14185 27455 14243 27461
rect 14185 27452 14197 27455
rect 14148 27424 14197 27452
rect 14148 27412 14154 27424
rect 14185 27421 14197 27424
rect 14231 27421 14243 27455
rect 14185 27415 14243 27421
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27452 14427 27455
rect 14826 27452 14832 27464
rect 14415 27424 14832 27452
rect 14415 27421 14427 27424
rect 14369 27415 14427 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 20806 27452 20812 27464
rect 20767 27424 20812 27452
rect 20806 27412 20812 27424
rect 20864 27412 20870 27464
rect 20990 27461 20996 27464
rect 20957 27455 20996 27461
rect 20957 27421 20969 27455
rect 20957 27415 20996 27421
rect 20990 27412 20996 27415
rect 21048 27412 21054 27464
rect 21315 27455 21373 27461
rect 21315 27421 21327 27455
rect 21361 27452 21373 27455
rect 21910 27452 21916 27464
rect 21361 27424 21916 27452
rect 21361 27421 21373 27424
rect 21315 27415 21373 27421
rect 21910 27412 21916 27424
rect 21968 27412 21974 27464
rect 22830 27452 22836 27464
rect 22791 27424 22836 27452
rect 22830 27412 22836 27424
rect 22888 27412 22894 27464
rect 23017 27455 23075 27461
rect 23017 27421 23029 27455
rect 23063 27421 23075 27455
rect 23017 27415 23075 27421
rect 23109 27455 23167 27461
rect 23109 27421 23121 27455
rect 23155 27421 23167 27455
rect 23382 27452 23388 27464
rect 23295 27424 23388 27452
rect 23109 27415 23167 27421
rect 12618 27384 12624 27396
rect 12098 27356 12624 27384
rect 12618 27344 12624 27356
rect 12676 27344 12682 27396
rect 13998 27344 14004 27396
rect 14056 27384 14062 27396
rect 14277 27387 14335 27393
rect 14277 27384 14289 27387
rect 14056 27356 14289 27384
rect 14056 27344 14062 27356
rect 14277 27353 14289 27356
rect 14323 27353 14335 27387
rect 21082 27384 21088 27396
rect 21043 27356 21088 27384
rect 14277 27347 14335 27353
rect 21082 27344 21088 27356
rect 21140 27344 21146 27396
rect 21177 27387 21235 27393
rect 21177 27353 21189 27387
rect 21223 27384 21235 27387
rect 21223 27356 21312 27384
rect 21223 27353 21235 27356
rect 21177 27347 21235 27353
rect 21284 27328 21312 27356
rect 22002 27344 22008 27396
rect 22060 27384 22066 27396
rect 23032 27384 23060 27415
rect 22060 27356 23060 27384
rect 23124 27384 23152 27415
rect 23382 27412 23388 27424
rect 23440 27452 23446 27464
rect 26329 27455 26387 27461
rect 23440 27424 24440 27452
rect 23440 27412 23446 27424
rect 23658 27384 23664 27396
rect 23124 27356 23664 27384
rect 22060 27344 22066 27356
rect 23658 27344 23664 27356
rect 23716 27344 23722 27396
rect 21266 27276 21272 27328
rect 21324 27276 21330 27328
rect 23566 27316 23572 27328
rect 23527 27288 23572 27316
rect 23566 27276 23572 27288
rect 23624 27276 23630 27328
rect 24412 27316 24440 27424
rect 26329 27421 26341 27455
rect 26375 27452 26387 27455
rect 27246 27452 27252 27464
rect 26375 27424 27252 27452
rect 26375 27421 26387 27424
rect 26329 27415 26387 27421
rect 27246 27412 27252 27424
rect 27304 27412 27310 27464
rect 29748 27461 29776 27560
rect 31018 27548 31024 27560
rect 31076 27548 31082 27600
rect 33594 27588 33600 27600
rect 33555 27560 33600 27588
rect 33594 27548 33600 27560
rect 33652 27548 33658 27600
rect 46934 27588 46940 27600
rect 46308 27560 46940 27588
rect 30009 27523 30067 27529
rect 30009 27489 30021 27523
rect 30055 27489 30067 27523
rect 45646 27520 45652 27532
rect 30009 27483 30067 27489
rect 31772 27492 45652 27520
rect 29733 27455 29791 27461
rect 29733 27421 29745 27455
rect 29779 27421 29791 27455
rect 29733 27415 29791 27421
rect 29822 27412 29828 27464
rect 29880 27452 29886 27464
rect 29880 27424 29925 27452
rect 29880 27412 29886 27424
rect 29362 27344 29368 27396
rect 29420 27384 29426 27396
rect 30024 27384 30052 27483
rect 31772 27461 31800 27492
rect 45646 27480 45652 27492
rect 45704 27480 45710 27532
rect 46308 27529 46336 27560
rect 46934 27548 46940 27560
rect 46992 27548 46998 27600
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46293 27483 46351 27489
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 47670 27520 47676 27532
rect 46523 27492 47676 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 47670 27480 47676 27492
rect 47728 27480 47734 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 30101 27455 30159 27461
rect 30101 27421 30113 27455
rect 30147 27421 30159 27455
rect 30101 27415 30159 27421
rect 31757 27455 31815 27461
rect 31757 27421 31769 27455
rect 31803 27421 31815 27455
rect 31757 27415 31815 27421
rect 31849 27455 31907 27461
rect 31849 27421 31861 27455
rect 31895 27452 31907 27455
rect 31938 27452 31944 27464
rect 31895 27424 31944 27452
rect 31895 27421 31907 27424
rect 31849 27415 31907 27421
rect 29420 27356 30052 27384
rect 29420 27344 29426 27356
rect 30116 27316 30144 27415
rect 31938 27412 31944 27424
rect 31996 27412 32002 27464
rect 32033 27455 32091 27461
rect 32033 27421 32045 27455
rect 32079 27421 32091 27455
rect 32033 27415 32091 27421
rect 31202 27344 31208 27396
rect 31260 27384 31266 27396
rect 31662 27384 31668 27396
rect 31260 27356 31668 27384
rect 31260 27344 31266 27356
rect 31662 27344 31668 27356
rect 31720 27384 31726 27396
rect 32048 27384 32076 27415
rect 32122 27412 32128 27464
rect 32180 27452 32186 27464
rect 33505 27455 33563 27461
rect 32180 27424 32225 27452
rect 32180 27412 32186 27424
rect 33505 27421 33517 27455
rect 33551 27452 33563 27455
rect 34606 27452 34612 27464
rect 33551 27424 34612 27452
rect 33551 27421 33563 27424
rect 33505 27415 33563 27421
rect 34606 27412 34612 27424
rect 34664 27412 34670 27464
rect 31720 27356 32076 27384
rect 31720 27344 31726 27356
rect 24412 27288 30144 27316
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 11238 27072 11244 27124
rect 11296 27112 11302 27124
rect 11793 27115 11851 27121
rect 11793 27112 11805 27115
rect 11296 27084 11805 27112
rect 11296 27072 11302 27084
rect 11793 27081 11805 27084
rect 11839 27081 11851 27115
rect 11793 27075 11851 27081
rect 26878 27072 26884 27124
rect 26936 27112 26942 27124
rect 27522 27112 27528 27124
rect 26936 27084 27528 27112
rect 26936 27072 26942 27084
rect 27522 27072 27528 27084
rect 27580 27112 27586 27124
rect 28353 27115 28411 27121
rect 28353 27112 28365 27115
rect 27580 27084 28365 27112
rect 27580 27072 27586 27084
rect 28353 27081 28365 27084
rect 28399 27081 28411 27115
rect 28353 27075 28411 27081
rect 11609 27047 11667 27053
rect 11609 27013 11621 27047
rect 11655 27044 11667 27047
rect 11698 27044 11704 27056
rect 11655 27016 11704 27044
rect 11655 27013 11667 27016
rect 11609 27007 11667 27013
rect 11698 27004 11704 27016
rect 11756 27004 11762 27056
rect 21266 27044 21272 27056
rect 20640 27016 21272 27044
rect 11514 26976 11520 26988
rect 11475 26948 11520 26976
rect 11514 26936 11520 26948
rect 11572 26936 11578 26988
rect 11882 26976 11888 26988
rect 11843 26948 11888 26976
rect 11882 26936 11888 26948
rect 11940 26936 11946 26988
rect 13814 26936 13820 26988
rect 13872 26976 13878 26988
rect 14093 26979 14151 26985
rect 14093 26976 14105 26979
rect 13872 26948 14105 26976
rect 13872 26936 13878 26948
rect 14093 26945 14105 26948
rect 14139 26976 14151 26979
rect 15102 26976 15108 26988
rect 14139 26948 15108 26976
rect 14139 26945 14151 26948
rect 14093 26939 14151 26945
rect 15102 26936 15108 26948
rect 15160 26976 15166 26988
rect 15286 26976 15292 26988
rect 15160 26948 15292 26976
rect 15160 26936 15166 26948
rect 15286 26936 15292 26948
rect 15344 26936 15350 26988
rect 20640 26985 20668 27016
rect 21266 27004 21272 27016
rect 21324 27004 21330 27056
rect 21910 27004 21916 27056
rect 21968 27044 21974 27056
rect 23109 27047 23167 27053
rect 23109 27044 23121 27047
rect 21968 27016 23121 27044
rect 21968 27004 21974 27016
rect 23109 27013 23121 27016
rect 23155 27044 23167 27047
rect 23382 27044 23388 27056
rect 23155 27016 23388 27044
rect 23155 27013 23167 27016
rect 23109 27007 23167 27013
rect 23382 27004 23388 27016
rect 23440 27004 23446 27056
rect 30650 27004 30656 27056
rect 30708 27044 30714 27056
rect 30929 27047 30987 27053
rect 30929 27044 30941 27047
rect 30708 27016 30941 27044
rect 30708 27004 30714 27016
rect 30929 27013 30941 27016
rect 30975 27013 30987 27047
rect 30929 27007 30987 27013
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26945 20683 26979
rect 20625 26939 20683 26945
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 21821 26979 21879 26985
rect 20772 26948 20817 26976
rect 20772 26936 20778 26948
rect 21821 26945 21833 26979
rect 21867 26976 21879 26979
rect 22462 26976 22468 26988
rect 21867 26948 22468 26976
rect 21867 26945 21879 26948
rect 21821 26939 21879 26945
rect 22462 26936 22468 26948
rect 22520 26936 22526 26988
rect 23293 26979 23351 26985
rect 23293 26945 23305 26979
rect 23339 26945 23351 26979
rect 23293 26939 23351 26945
rect 23937 26979 23995 26985
rect 23937 26945 23949 26979
rect 23983 26945 23995 26979
rect 24118 26976 24124 26988
rect 24079 26948 24124 26976
rect 23937 26939 23995 26945
rect 11701 26911 11759 26917
rect 11701 26877 11713 26911
rect 11747 26908 11759 26911
rect 12158 26908 12164 26920
rect 11747 26880 12164 26908
rect 11747 26877 11759 26880
rect 11701 26871 11759 26877
rect 12158 26868 12164 26880
rect 12216 26868 12222 26920
rect 22094 26868 22100 26920
rect 22152 26908 22158 26920
rect 23308 26908 23336 26939
rect 23658 26908 23664 26920
rect 22152 26880 22197 26908
rect 23308 26880 23664 26908
rect 22152 26868 22158 26880
rect 23658 26868 23664 26880
rect 23716 26868 23722 26920
rect 21174 26840 21180 26852
rect 20824 26812 21180 26840
rect 14182 26772 14188 26784
rect 14143 26744 14188 26772
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 20824 26781 20852 26812
rect 21174 26800 21180 26812
rect 21232 26800 21238 26852
rect 21358 26800 21364 26852
rect 21416 26840 21422 26852
rect 23477 26843 23535 26849
rect 23477 26840 23489 26843
rect 21416 26812 23489 26840
rect 21416 26800 21422 26812
rect 23477 26809 23489 26812
rect 23523 26840 23535 26843
rect 23952 26840 23980 26939
rect 24118 26936 24124 26948
rect 24176 26936 24182 26988
rect 25682 26976 25688 26988
rect 25643 26948 25688 26976
rect 25682 26936 25688 26948
rect 25740 26936 25746 26988
rect 28166 26976 28172 26988
rect 28127 26948 28172 26976
rect 28166 26936 28172 26948
rect 28224 26976 28230 26988
rect 28902 26976 28908 26988
rect 28224 26948 28908 26976
rect 28224 26936 28230 26948
rect 28902 26936 28908 26948
rect 28960 26936 28966 26988
rect 31110 26976 31116 26988
rect 31071 26948 31116 26976
rect 31110 26936 31116 26948
rect 31168 26936 31174 26988
rect 31205 26979 31263 26985
rect 31205 26945 31217 26979
rect 31251 26976 31263 26979
rect 32214 26976 32220 26988
rect 31251 26948 32220 26976
rect 31251 26945 31263 26948
rect 31205 26939 31263 26945
rect 32214 26936 32220 26948
rect 32272 26936 32278 26988
rect 25774 26908 25780 26920
rect 25735 26880 25780 26908
rect 25774 26868 25780 26880
rect 25832 26868 25838 26920
rect 24394 26840 24400 26852
rect 23523 26812 24400 26840
rect 23523 26809 23535 26812
rect 23477 26803 23535 26809
rect 24394 26800 24400 26812
rect 24452 26800 24458 26852
rect 25590 26800 25596 26852
rect 25648 26840 25654 26852
rect 26053 26843 26111 26849
rect 26053 26840 26065 26843
rect 25648 26812 26065 26840
rect 25648 26800 25654 26812
rect 26053 26809 26065 26812
rect 26099 26809 26111 26843
rect 26053 26803 26111 26809
rect 20809 26775 20867 26781
rect 20809 26741 20821 26775
rect 20855 26741 20867 26775
rect 20809 26735 20867 26741
rect 20993 26775 21051 26781
rect 20993 26741 21005 26775
rect 21039 26772 21051 26775
rect 21542 26772 21548 26784
rect 21039 26744 21548 26772
rect 21039 26741 21051 26744
rect 20993 26735 21051 26741
rect 21542 26732 21548 26744
rect 21600 26732 21606 26784
rect 23842 26732 23848 26784
rect 23900 26772 23906 26784
rect 23937 26775 23995 26781
rect 23937 26772 23949 26775
rect 23900 26744 23949 26772
rect 23900 26732 23906 26744
rect 23937 26741 23949 26744
rect 23983 26741 23995 26775
rect 23937 26735 23995 26741
rect 25869 26775 25927 26781
rect 25869 26741 25881 26775
rect 25915 26772 25927 26775
rect 26234 26772 26240 26784
rect 25915 26744 26240 26772
rect 25915 26741 25927 26744
rect 25869 26735 25927 26741
rect 26234 26732 26240 26744
rect 26292 26772 26298 26784
rect 27062 26772 27068 26784
rect 26292 26744 27068 26772
rect 26292 26732 26298 26744
rect 27062 26732 27068 26744
rect 27120 26732 27126 26784
rect 30929 26775 30987 26781
rect 30929 26741 30941 26775
rect 30975 26772 30987 26775
rect 31202 26772 31208 26784
rect 30975 26744 31208 26772
rect 30975 26741 30987 26744
rect 30929 26735 30987 26741
rect 31202 26732 31208 26744
rect 31260 26732 31266 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 2038 26528 2044 26580
rect 2096 26568 2102 26580
rect 2096 26540 28672 26568
rect 2096 26528 2102 26540
rect 11514 26460 11520 26512
rect 11572 26500 11578 26512
rect 12250 26500 12256 26512
rect 11572 26472 12256 26500
rect 11572 26460 11578 26472
rect 12250 26460 12256 26472
rect 12308 26460 12314 26512
rect 14090 26460 14096 26512
rect 14148 26500 14154 26512
rect 15473 26503 15531 26509
rect 15473 26500 15485 26503
rect 14148 26472 15485 26500
rect 14148 26460 14154 26472
rect 15473 26469 15485 26472
rect 15519 26469 15531 26503
rect 15473 26463 15531 26469
rect 16577 26503 16635 26509
rect 16577 26469 16589 26503
rect 16623 26469 16635 26503
rect 16577 26463 16635 26469
rect 13998 26392 14004 26444
rect 14056 26432 14062 26444
rect 14185 26435 14243 26441
rect 14185 26432 14197 26435
rect 14056 26404 14197 26432
rect 14056 26392 14062 26404
rect 14185 26401 14197 26404
rect 14231 26401 14243 26435
rect 16592 26432 16620 26463
rect 20346 26460 20352 26512
rect 20404 26500 20410 26512
rect 21174 26500 21180 26512
rect 20404 26472 21180 26500
rect 20404 26460 20410 26472
rect 21174 26460 21180 26472
rect 21232 26460 21238 26512
rect 21542 26460 21548 26512
rect 21600 26500 21606 26512
rect 21600 26472 21645 26500
rect 21600 26460 21606 26472
rect 21726 26460 21732 26512
rect 21784 26500 21790 26512
rect 23293 26503 23351 26509
rect 23293 26500 23305 26503
rect 21784 26472 23305 26500
rect 21784 26460 21790 26472
rect 23293 26469 23305 26472
rect 23339 26500 23351 26503
rect 24118 26500 24124 26512
rect 23339 26472 24124 26500
rect 23339 26469 23351 26472
rect 23293 26463 23351 26469
rect 24118 26460 24124 26472
rect 24176 26500 24182 26512
rect 26510 26500 26516 26512
rect 24176 26472 24624 26500
rect 24176 26460 24182 26472
rect 16592 26404 18092 26432
rect 14185 26395 14243 26401
rect 9950 26324 9956 26376
rect 10008 26364 10014 26376
rect 10045 26367 10103 26373
rect 10045 26364 10057 26367
rect 10008 26336 10057 26364
rect 10008 26324 10014 26336
rect 10045 26333 10057 26336
rect 10091 26333 10103 26367
rect 10045 26327 10103 26333
rect 11974 26324 11980 26376
rect 12032 26364 12038 26376
rect 12069 26367 12127 26373
rect 12069 26364 12081 26367
rect 12032 26336 12081 26364
rect 12032 26324 12038 26336
rect 12069 26333 12081 26336
rect 12115 26364 12127 26367
rect 14090 26364 14096 26376
rect 12115 26336 14096 26364
rect 12115 26333 12127 26336
rect 12069 26327 12127 26333
rect 14090 26324 14096 26336
rect 14148 26324 14154 26376
rect 14274 26364 14280 26376
rect 14235 26336 14280 26364
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 15010 26324 15016 26376
rect 15068 26364 15074 26376
rect 15105 26367 15163 26373
rect 15105 26364 15117 26367
rect 15068 26336 15117 26364
rect 15068 26324 15074 26336
rect 15105 26333 15117 26336
rect 15151 26333 15163 26367
rect 15105 26327 15163 26333
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26333 15347 26367
rect 16574 26364 16580 26376
rect 16535 26336 16580 26364
rect 15289 26327 15347 26333
rect 14734 26256 14740 26308
rect 14792 26296 14798 26308
rect 15304 26296 15332 26327
rect 16574 26324 16580 26336
rect 16632 26324 16638 26376
rect 16850 26364 16856 26376
rect 16811 26336 16856 26364
rect 16850 26324 16856 26336
rect 16908 26324 16914 26376
rect 16942 26324 16948 26376
rect 17000 26364 17006 26376
rect 18064 26373 18092 26404
rect 20898 26392 20904 26444
rect 20956 26432 20962 26444
rect 21358 26432 21364 26444
rect 20956 26404 21364 26432
rect 20956 26392 20962 26404
rect 21358 26392 21364 26404
rect 21416 26441 21422 26444
rect 21416 26435 21474 26441
rect 21416 26401 21428 26435
rect 21462 26401 21474 26435
rect 21416 26395 21474 26401
rect 21637 26435 21695 26441
rect 21637 26401 21649 26435
rect 21683 26432 21695 26435
rect 22554 26432 22560 26444
rect 21683 26404 22560 26432
rect 21683 26401 21695 26404
rect 21637 26395 21695 26401
rect 21416 26392 21422 26395
rect 22554 26392 22560 26404
rect 22612 26392 22618 26444
rect 23382 26432 23388 26444
rect 23343 26404 23388 26432
rect 23382 26392 23388 26404
rect 23440 26392 23446 26444
rect 17313 26367 17371 26373
rect 17313 26364 17325 26367
rect 17000 26336 17325 26364
rect 17000 26324 17006 26336
rect 17313 26333 17325 26336
rect 17359 26333 17371 26367
rect 17313 26327 17371 26333
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26333 18107 26367
rect 18049 26327 18107 26333
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26364 18291 26367
rect 19978 26364 19984 26376
rect 18279 26336 19984 26364
rect 18279 26333 18291 26336
rect 18233 26327 18291 26333
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 20441 26367 20499 26373
rect 20441 26333 20453 26367
rect 20487 26364 20499 26367
rect 21542 26364 21548 26376
rect 20487 26336 21548 26364
rect 20487 26333 20499 26336
rect 20441 26327 20499 26333
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26333 23167 26367
rect 24394 26364 24400 26376
rect 24355 26336 24400 26364
rect 23109 26327 23167 26333
rect 14792 26268 15332 26296
rect 16592 26296 16620 26324
rect 18874 26296 18880 26308
rect 16592 26268 18880 26296
rect 14792 26256 14798 26268
rect 18874 26256 18880 26268
rect 18932 26256 18938 26308
rect 20346 26256 20352 26308
rect 20404 26296 20410 26308
rect 20625 26299 20683 26305
rect 20625 26296 20637 26299
rect 20404 26268 20637 26296
rect 20404 26256 20410 26268
rect 20625 26265 20637 26268
rect 20671 26265 20683 26299
rect 20625 26259 20683 26265
rect 20809 26299 20867 26305
rect 20809 26265 20821 26299
rect 20855 26296 20867 26299
rect 20990 26296 20996 26308
rect 20855 26268 20996 26296
rect 20855 26265 20867 26268
rect 20809 26259 20867 26265
rect 20990 26256 20996 26268
rect 21048 26296 21054 26308
rect 21266 26296 21272 26308
rect 21048 26268 21128 26296
rect 21227 26268 21272 26296
rect 21048 26256 21054 26268
rect 10226 26228 10232 26240
rect 10187 26200 10232 26228
rect 10226 26188 10232 26200
rect 10284 26188 10290 26240
rect 13814 26188 13820 26240
rect 13872 26228 13878 26240
rect 14645 26231 14703 26237
rect 14645 26228 14657 26231
rect 13872 26200 14657 26228
rect 13872 26188 13878 26200
rect 14645 26197 14657 26200
rect 14691 26197 14703 26231
rect 14645 26191 14703 26197
rect 16666 26188 16672 26240
rect 16724 26228 16730 26240
rect 16761 26231 16819 26237
rect 16761 26228 16773 26231
rect 16724 26200 16773 26228
rect 16724 26188 16730 26200
rect 16761 26197 16773 26200
rect 16807 26197 16819 26231
rect 16761 26191 16819 26197
rect 17126 26188 17132 26240
rect 17184 26228 17190 26240
rect 17497 26231 17555 26237
rect 17497 26228 17509 26231
rect 17184 26200 17509 26228
rect 17184 26188 17190 26200
rect 17497 26197 17509 26200
rect 17543 26197 17555 26231
rect 18138 26228 18144 26240
rect 18099 26200 18144 26228
rect 17497 26191 17555 26197
rect 18138 26188 18144 26200
rect 18196 26188 18202 26240
rect 21100 26228 21128 26268
rect 21266 26256 21272 26268
rect 21324 26256 21330 26308
rect 21726 26296 21732 26308
rect 21376 26268 21732 26296
rect 21376 26228 21404 26268
rect 21726 26256 21732 26268
rect 21784 26256 21790 26308
rect 21818 26256 21824 26308
rect 21876 26296 21882 26308
rect 22005 26299 22063 26305
rect 22005 26296 22017 26299
rect 21876 26268 22017 26296
rect 21876 26256 21882 26268
rect 22005 26265 22017 26268
rect 22051 26265 22063 26299
rect 23124 26296 23152 26327
rect 24394 26324 24400 26336
rect 24452 26324 24458 26376
rect 24596 26373 24624 26472
rect 26436 26472 26516 26500
rect 24765 26435 24823 26441
rect 24765 26401 24777 26435
rect 24811 26432 24823 26435
rect 25682 26432 25688 26444
rect 24811 26404 25688 26432
rect 24811 26401 24823 26404
rect 24765 26395 24823 26401
rect 25682 26392 25688 26404
rect 25740 26432 25746 26444
rect 25740 26404 26280 26432
rect 25740 26392 25746 26404
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26333 24639 26367
rect 26142 26364 26148 26376
rect 26103 26336 26148 26364
rect 24581 26327 24639 26333
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 26252 26373 26280 26404
rect 26237 26367 26295 26373
rect 26237 26333 26249 26367
rect 26283 26333 26295 26367
rect 26237 26327 26295 26333
rect 26329 26367 26387 26373
rect 26329 26333 26341 26367
rect 26375 26364 26387 26367
rect 26436 26364 26464 26472
rect 26510 26460 26516 26472
rect 26568 26460 26574 26512
rect 27522 26392 27528 26444
rect 27580 26432 27586 26444
rect 27580 26404 28580 26432
rect 27580 26392 27586 26404
rect 26375 26336 26464 26364
rect 26375 26333 26387 26336
rect 26329 26327 26387 26333
rect 26510 26324 26516 26376
rect 26568 26364 26574 26376
rect 27062 26364 27068 26376
rect 26568 26336 26613 26364
rect 27023 26336 27068 26364
rect 26568 26324 26574 26336
rect 27062 26324 27068 26336
rect 27120 26324 27126 26376
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26364 27215 26367
rect 27246 26364 27252 26376
rect 27203 26336 27252 26364
rect 27203 26333 27215 26336
rect 27157 26327 27215 26333
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 28552 26373 28580 26404
rect 28644 26373 28672 26540
rect 28902 26528 28908 26580
rect 28960 26568 28966 26580
rect 30929 26571 30987 26577
rect 30929 26568 30941 26571
rect 28960 26540 30941 26568
rect 28960 26528 28966 26540
rect 30929 26537 30941 26540
rect 30975 26537 30987 26571
rect 32674 26568 32680 26580
rect 30929 26531 30987 26537
rect 31680 26540 32680 26568
rect 29549 26503 29607 26509
rect 29549 26469 29561 26503
rect 29595 26469 29607 26503
rect 29549 26463 29607 26469
rect 29564 26432 29592 26463
rect 28828 26404 29592 26432
rect 30193 26435 30251 26441
rect 28353 26367 28411 26373
rect 28353 26333 28365 26367
rect 28399 26333 28411 26367
rect 28353 26327 28411 26333
rect 28537 26367 28595 26373
rect 28537 26333 28549 26367
rect 28583 26333 28595 26367
rect 28537 26327 28595 26333
rect 28629 26367 28687 26373
rect 28629 26333 28641 26367
rect 28675 26333 28687 26367
rect 28629 26327 28687 26333
rect 23658 26296 23664 26308
rect 23124 26268 23664 26296
rect 22005 26259 22063 26265
rect 23658 26256 23664 26268
rect 23716 26256 23722 26308
rect 25869 26299 25927 26305
rect 25869 26265 25881 26299
rect 25915 26296 25927 26299
rect 26970 26296 26976 26308
rect 25915 26268 26976 26296
rect 25915 26265 25927 26268
rect 25869 26259 25927 26265
rect 26970 26256 26976 26268
rect 27028 26256 27034 26308
rect 28169 26299 28227 26305
rect 28169 26265 28181 26299
rect 28215 26296 28227 26299
rect 28258 26296 28264 26308
rect 28215 26268 28264 26296
rect 28215 26265 28227 26268
rect 28169 26259 28227 26265
rect 28258 26256 28264 26268
rect 28316 26256 28322 26308
rect 28368 26296 28396 26327
rect 28828 26296 28856 26404
rect 30193 26401 30205 26435
rect 30239 26432 30251 26435
rect 30374 26432 30380 26444
rect 30239 26404 30380 26432
rect 30239 26401 30251 26404
rect 30193 26395 30251 26401
rect 30374 26392 30380 26404
rect 30432 26392 30438 26444
rect 29178 26324 29184 26376
rect 29236 26364 29242 26376
rect 29917 26367 29975 26373
rect 29917 26364 29929 26367
rect 29236 26336 29929 26364
rect 29236 26324 29242 26336
rect 29917 26333 29929 26336
rect 29963 26333 29975 26367
rect 29917 26327 29975 26333
rect 28368 26268 28856 26296
rect 29546 26256 29552 26308
rect 29604 26296 29610 26308
rect 30009 26299 30067 26305
rect 30009 26296 30021 26299
rect 29604 26268 30021 26296
rect 29604 26256 29610 26268
rect 30009 26265 30021 26268
rect 30055 26265 30067 26299
rect 30834 26296 30840 26308
rect 30795 26268 30840 26296
rect 30009 26259 30067 26265
rect 30834 26256 30840 26268
rect 30892 26256 30898 26308
rect 30944 26296 30972 26531
rect 31680 26373 31708 26540
rect 32674 26528 32680 26540
rect 32732 26528 32738 26580
rect 32766 26528 32772 26580
rect 32824 26568 32830 26580
rect 33137 26571 33195 26577
rect 33137 26568 33149 26571
rect 32824 26540 33149 26568
rect 32824 26528 32830 26540
rect 33137 26537 33149 26540
rect 33183 26537 33195 26571
rect 33137 26531 33195 26537
rect 33502 26528 33508 26580
rect 33560 26568 33566 26580
rect 33597 26571 33655 26577
rect 33597 26568 33609 26571
rect 33560 26540 33609 26568
rect 33560 26528 33566 26540
rect 33597 26537 33609 26540
rect 33643 26537 33655 26571
rect 33597 26531 33655 26537
rect 32217 26503 32275 26509
rect 32217 26469 32229 26503
rect 32263 26500 32275 26503
rect 33962 26500 33968 26512
rect 32263 26472 33968 26500
rect 32263 26469 32275 26472
rect 32217 26463 32275 26469
rect 33962 26460 33968 26472
rect 34020 26460 34026 26512
rect 32582 26392 32588 26444
rect 32640 26432 32646 26444
rect 32769 26435 32827 26441
rect 32769 26432 32781 26435
rect 32640 26404 32781 26432
rect 32640 26392 32646 26404
rect 32769 26401 32781 26404
rect 32815 26401 32827 26435
rect 32769 26395 32827 26401
rect 33686 26392 33692 26444
rect 33744 26432 33750 26444
rect 34057 26435 34115 26441
rect 34057 26432 34069 26435
rect 33744 26404 34069 26432
rect 33744 26392 33750 26404
rect 34057 26401 34069 26404
rect 34103 26401 34115 26435
rect 34057 26395 34115 26401
rect 31665 26367 31723 26373
rect 31665 26333 31677 26367
rect 31711 26333 31723 26367
rect 31665 26327 31723 26333
rect 31754 26324 31760 26376
rect 31812 26364 31818 26376
rect 31849 26367 31907 26373
rect 31849 26364 31861 26367
rect 31812 26336 31861 26364
rect 31812 26324 31818 26336
rect 31849 26333 31861 26336
rect 31895 26333 31907 26367
rect 32030 26364 32036 26376
rect 31991 26336 32036 26364
rect 31849 26327 31907 26333
rect 32030 26324 32036 26336
rect 32088 26324 32094 26376
rect 32953 26367 33011 26373
rect 32953 26333 32965 26367
rect 32999 26364 33011 26367
rect 33778 26364 33784 26376
rect 32999 26336 33784 26364
rect 32999 26333 33011 26336
rect 32953 26327 33011 26333
rect 33778 26324 33784 26336
rect 33836 26324 33842 26376
rect 33965 26367 34023 26373
rect 33965 26333 33977 26367
rect 34011 26333 34023 26367
rect 33965 26327 34023 26333
rect 31938 26296 31944 26308
rect 30944 26268 31944 26296
rect 31938 26256 31944 26268
rect 31996 26256 32002 26308
rect 32122 26256 32128 26308
rect 32180 26296 32186 26308
rect 32677 26299 32735 26305
rect 32677 26296 32689 26299
rect 32180 26268 32689 26296
rect 32180 26256 32186 26268
rect 32677 26265 32689 26268
rect 32723 26265 32735 26299
rect 32677 26259 32735 26265
rect 33042 26256 33048 26308
rect 33100 26296 33106 26308
rect 33980 26296 34008 26327
rect 46382 26324 46388 26376
rect 46440 26364 46446 26376
rect 47673 26367 47731 26373
rect 47673 26364 47685 26367
rect 46440 26336 47685 26364
rect 46440 26324 46446 26336
rect 47673 26333 47685 26336
rect 47719 26333 47731 26367
rect 47673 26327 47731 26333
rect 33100 26268 34008 26296
rect 33100 26256 33106 26268
rect 21100 26200 21404 26228
rect 22925 26231 22983 26237
rect 22925 26197 22937 26231
rect 22971 26228 22983 26231
rect 23014 26228 23020 26240
rect 22971 26200 23020 26228
rect 22971 26197 22983 26200
rect 22925 26191 22983 26197
rect 23014 26188 23020 26200
rect 23072 26188 23078 26240
rect 26234 26188 26240 26240
rect 26292 26228 26298 26240
rect 27341 26231 27399 26237
rect 27341 26228 27353 26231
rect 26292 26200 27353 26228
rect 26292 26188 26298 26200
rect 27341 26197 27353 26200
rect 27387 26197 27399 26231
rect 27341 26191 27399 26197
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 12250 25984 12256 26036
rect 12308 26024 12314 26036
rect 18874 26024 18880 26036
rect 12308 25996 15148 26024
rect 18835 25996 18880 26024
rect 12308 25984 12314 25996
rect 10321 25891 10379 25897
rect 10321 25857 10333 25891
rect 10367 25888 10379 25891
rect 11790 25888 11796 25900
rect 10367 25860 11796 25888
rect 10367 25857 10379 25860
rect 10321 25851 10379 25857
rect 11790 25848 11796 25860
rect 11848 25848 11854 25900
rect 10413 25823 10471 25829
rect 10413 25789 10425 25823
rect 10459 25820 10471 25823
rect 10962 25820 10968 25832
rect 10459 25792 10968 25820
rect 10459 25789 10471 25792
rect 10413 25783 10471 25789
rect 10962 25780 10968 25792
rect 11020 25820 11026 25832
rect 12268 25820 12296 25984
rect 13541 25959 13599 25965
rect 13541 25925 13553 25959
rect 13587 25956 13599 25959
rect 13814 25956 13820 25968
rect 13587 25928 13820 25956
rect 13587 25925 13599 25928
rect 13541 25919 13599 25925
rect 13814 25916 13820 25928
rect 13872 25916 13878 25968
rect 14182 25916 14188 25968
rect 14240 25916 14246 25968
rect 12713 25891 12771 25897
rect 12713 25857 12725 25891
rect 12759 25857 12771 25891
rect 15120 25888 15148 25996
rect 18874 25984 18880 25996
rect 18932 25984 18938 26036
rect 19889 26027 19947 26033
rect 19889 25993 19901 26027
rect 19935 26024 19947 26027
rect 20806 26024 20812 26036
rect 19935 25996 20812 26024
rect 19935 25993 19947 25996
rect 19889 25987 19947 25993
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 27341 26027 27399 26033
rect 27341 26024 27353 26027
rect 22066 25996 27353 26024
rect 16025 25959 16083 25965
rect 16025 25925 16037 25959
rect 16071 25956 16083 25959
rect 16574 25956 16580 25968
rect 16071 25928 16580 25956
rect 16071 25925 16083 25928
rect 16025 25919 16083 25925
rect 16574 25916 16580 25928
rect 16632 25916 16638 25968
rect 19978 25916 19984 25968
rect 20036 25956 20042 25968
rect 20441 25959 20499 25965
rect 20441 25956 20453 25959
rect 20036 25928 20453 25956
rect 20036 25916 20042 25928
rect 20441 25925 20453 25928
rect 20487 25956 20499 25959
rect 20622 25956 20628 25968
rect 20487 25928 20628 25956
rect 20487 25925 20499 25928
rect 20441 25919 20499 25925
rect 20622 25916 20628 25928
rect 20680 25916 20686 25968
rect 16117 25891 16175 25897
rect 16117 25888 16129 25891
rect 15120 25860 16129 25888
rect 12713 25851 12771 25857
rect 16117 25857 16129 25860
rect 16163 25888 16175 25891
rect 16850 25888 16856 25900
rect 16163 25860 16856 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 11020 25792 12296 25820
rect 11020 25780 11026 25792
rect 12728 25752 12756 25851
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 17126 25888 17132 25900
rect 17087 25860 17132 25888
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 19334 25888 19340 25900
rect 18538 25860 19340 25888
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 19705 25891 19763 25897
rect 19705 25857 19717 25891
rect 19751 25888 19763 25891
rect 20346 25888 20352 25900
rect 19751 25860 20352 25888
rect 19751 25857 19763 25860
rect 19705 25851 19763 25857
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 20714 25888 20720 25900
rect 20675 25860 20720 25888
rect 20714 25848 20720 25860
rect 20772 25848 20778 25900
rect 20898 25888 20904 25900
rect 20859 25860 20904 25888
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 21174 25888 21180 25900
rect 21135 25860 21180 25888
rect 21174 25848 21180 25860
rect 21232 25848 21238 25900
rect 12805 25823 12863 25829
rect 12805 25789 12817 25823
rect 12851 25820 12863 25823
rect 13265 25823 13323 25829
rect 13265 25820 13277 25823
rect 12851 25792 13277 25820
rect 12851 25789 12863 25792
rect 12805 25783 12863 25789
rect 13265 25789 13277 25792
rect 13311 25789 13323 25823
rect 13906 25820 13912 25832
rect 13265 25783 13323 25789
rect 13372 25792 13912 25820
rect 13372 25752 13400 25792
rect 13906 25780 13912 25792
rect 13964 25820 13970 25832
rect 14918 25820 14924 25832
rect 13964 25792 14924 25820
rect 13964 25780 13970 25792
rect 14918 25780 14924 25792
rect 14976 25780 14982 25832
rect 15654 25820 15660 25832
rect 15615 25792 15660 25820
rect 15654 25780 15660 25792
rect 15712 25780 15718 25832
rect 17405 25823 17463 25829
rect 17405 25789 17417 25823
rect 17451 25820 17463 25823
rect 18138 25820 18144 25832
rect 17451 25792 18144 25820
rect 17451 25789 17463 25792
rect 17405 25783 17463 25789
rect 18138 25780 18144 25792
rect 18196 25780 18202 25832
rect 19518 25820 19524 25832
rect 19479 25792 19524 25820
rect 19518 25780 19524 25792
rect 19576 25780 19582 25832
rect 20993 25823 21051 25829
rect 20993 25789 21005 25823
rect 21039 25820 21051 25823
rect 21542 25820 21548 25832
rect 21039 25792 21548 25820
rect 21039 25789 21051 25792
rect 20993 25783 21051 25789
rect 21542 25780 21548 25792
rect 21600 25780 21606 25832
rect 12728 25724 13400 25752
rect 20809 25755 20867 25761
rect 20809 25721 20821 25755
rect 20855 25752 20867 25755
rect 21266 25752 21272 25764
rect 20855 25724 21272 25752
rect 20855 25721 20867 25724
rect 20809 25715 20867 25721
rect 21266 25712 21272 25724
rect 21324 25752 21330 25764
rect 22066 25752 22094 25996
rect 27341 25993 27353 25996
rect 27387 25993 27399 26027
rect 29825 26027 29883 26033
rect 29825 26024 29837 26027
rect 27341 25987 27399 25993
rect 28368 25996 29837 26024
rect 24486 25956 24492 25968
rect 24242 25928 24492 25956
rect 24486 25916 24492 25928
rect 24544 25916 24550 25968
rect 28368 25965 28396 25996
rect 29825 25993 29837 25996
rect 29871 26024 29883 26027
rect 30834 26024 30840 26036
rect 29871 25996 30840 26024
rect 29871 25993 29883 25996
rect 29825 25987 29883 25993
rect 30834 25984 30840 25996
rect 30892 25984 30898 26036
rect 31110 25984 31116 26036
rect 31168 26024 31174 26036
rect 31573 26027 31631 26033
rect 31573 26024 31585 26027
rect 31168 25996 31585 26024
rect 31168 25984 31174 25996
rect 31573 25993 31585 25996
rect 31619 26024 31631 26027
rect 32214 26024 32220 26036
rect 31619 25996 31754 26024
rect 32175 25996 32220 26024
rect 31619 25993 31631 25996
rect 31573 25987 31631 25993
rect 26053 25959 26111 25965
rect 26053 25925 26065 25959
rect 26099 25956 26111 25959
rect 28353 25959 28411 25965
rect 26099 25928 27292 25956
rect 26099 25925 26111 25928
rect 26053 25919 26111 25925
rect 25774 25888 25780 25900
rect 25735 25860 25780 25888
rect 25774 25848 25780 25860
rect 25832 25888 25838 25900
rect 26510 25888 26516 25900
rect 25832 25860 26516 25888
rect 25832 25848 25838 25860
rect 26510 25848 26516 25860
rect 26568 25888 26574 25900
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 26568 25860 26985 25888
rect 26568 25848 26574 25860
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 27154 25888 27160 25900
rect 27115 25860 27160 25888
rect 26973 25851 27031 25857
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 27264 25888 27292 25928
rect 28353 25925 28365 25959
rect 28399 25925 28411 25959
rect 28353 25919 28411 25925
rect 29546 25916 29552 25968
rect 29604 25956 29610 25968
rect 31726 25956 31754 25996
rect 32214 25984 32220 25996
rect 32272 25984 32278 26036
rect 33321 26027 33379 26033
rect 33321 25993 33333 26027
rect 33367 25993 33379 26027
rect 33321 25987 33379 25993
rect 33042 25956 33048 25968
rect 29604 25928 30420 25956
rect 31726 25928 33048 25956
rect 29604 25916 29610 25928
rect 27706 25888 27712 25900
rect 27264 25860 27712 25888
rect 27706 25848 27712 25860
rect 27764 25888 27770 25900
rect 28537 25891 28595 25897
rect 28537 25888 28549 25891
rect 27764 25860 28549 25888
rect 27764 25848 27770 25860
rect 28537 25857 28549 25860
rect 28583 25857 28595 25891
rect 28537 25851 28595 25857
rect 28626 25848 28632 25900
rect 28684 25888 28690 25900
rect 29733 25891 29791 25897
rect 28684 25860 28729 25888
rect 28684 25848 28690 25860
rect 29733 25857 29745 25891
rect 29779 25888 29791 25891
rect 29914 25888 29920 25900
rect 29779 25860 29920 25888
rect 29779 25857 29791 25860
rect 29733 25851 29791 25857
rect 22741 25823 22799 25829
rect 22741 25789 22753 25823
rect 22787 25820 22799 25823
rect 23017 25823 23075 25829
rect 22787 25792 22876 25820
rect 22787 25789 22799 25792
rect 22741 25783 22799 25789
rect 21324 25724 22094 25752
rect 21324 25712 21330 25724
rect 10502 25644 10508 25696
rect 10560 25684 10566 25696
rect 10689 25687 10747 25693
rect 10689 25684 10701 25687
rect 10560 25656 10701 25684
rect 10560 25644 10566 25656
rect 10689 25653 10701 25656
rect 10735 25653 10747 25687
rect 10689 25647 10747 25653
rect 14090 25644 14096 25696
rect 14148 25684 14154 25696
rect 14274 25684 14280 25696
rect 14148 25656 14280 25684
rect 14148 25644 14154 25656
rect 14274 25644 14280 25656
rect 14332 25684 14338 25696
rect 15013 25687 15071 25693
rect 15013 25684 15025 25687
rect 14332 25656 15025 25684
rect 14332 25644 14338 25656
rect 15013 25653 15025 25656
rect 15059 25684 15071 25687
rect 15102 25684 15108 25696
rect 15059 25656 15108 25684
rect 15059 25653 15071 25656
rect 15013 25647 15071 25653
rect 15102 25644 15108 25656
rect 15160 25644 15166 25696
rect 15841 25687 15899 25693
rect 15841 25653 15853 25687
rect 15887 25684 15899 25687
rect 16942 25684 16948 25696
rect 15887 25656 16948 25684
rect 15887 25653 15899 25656
rect 15841 25647 15899 25653
rect 16942 25644 16948 25656
rect 17000 25644 17006 25696
rect 22848 25684 22876 25792
rect 23017 25789 23029 25823
rect 23063 25820 23075 25823
rect 23566 25820 23572 25832
rect 23063 25792 23572 25820
rect 23063 25789 23075 25792
rect 23017 25783 23075 25789
rect 23566 25780 23572 25792
rect 23624 25780 23630 25832
rect 23658 25780 23664 25832
rect 23716 25820 23722 25832
rect 24489 25823 24547 25829
rect 24489 25820 24501 25823
rect 23716 25792 24501 25820
rect 23716 25780 23722 25792
rect 24489 25789 24501 25792
rect 24535 25789 24547 25823
rect 24489 25783 24547 25789
rect 26145 25823 26203 25829
rect 26145 25789 26157 25823
rect 26191 25789 26203 25823
rect 26145 25783 26203 25789
rect 24026 25712 24032 25764
rect 24084 25752 24090 25764
rect 26160 25752 26188 25783
rect 26234 25780 26240 25832
rect 26292 25829 26298 25832
rect 26292 25823 26320 25829
rect 26308 25789 26320 25823
rect 26292 25783 26320 25789
rect 26292 25780 26298 25783
rect 27430 25780 27436 25832
rect 27488 25820 27494 25832
rect 29748 25820 29776 25851
rect 29914 25848 29920 25860
rect 29972 25848 29978 25900
rect 30392 25897 30420 25928
rect 33042 25916 33048 25928
rect 33100 25916 33106 25968
rect 33336 25956 33364 25987
rect 33336 25928 34284 25956
rect 30377 25891 30435 25897
rect 30377 25857 30389 25891
rect 30423 25857 30435 25891
rect 30377 25851 30435 25857
rect 30466 25848 30472 25900
rect 30524 25888 30530 25900
rect 31205 25891 31263 25897
rect 31205 25888 31217 25891
rect 30524 25860 31217 25888
rect 30524 25848 30530 25860
rect 31205 25857 31217 25860
rect 31251 25857 31263 25891
rect 31386 25888 31392 25900
rect 31347 25860 31392 25888
rect 31205 25851 31263 25857
rect 27488 25792 29776 25820
rect 31220 25820 31248 25851
rect 31386 25848 31392 25860
rect 31444 25848 31450 25900
rect 32122 25888 32128 25900
rect 31726 25860 32128 25888
rect 31726 25820 31754 25860
rect 32122 25848 32128 25860
rect 32180 25848 32186 25900
rect 32309 25891 32367 25897
rect 32309 25857 32321 25891
rect 32355 25888 32367 25891
rect 32582 25888 32588 25900
rect 32355 25860 32588 25888
rect 32355 25857 32367 25860
rect 32309 25851 32367 25857
rect 32582 25848 32588 25860
rect 32640 25848 32646 25900
rect 32674 25848 32680 25900
rect 32732 25888 32738 25900
rect 32953 25891 33011 25897
rect 32953 25888 32965 25891
rect 32732 25860 32965 25888
rect 32732 25848 32738 25860
rect 32953 25857 32965 25860
rect 32999 25888 33011 25891
rect 33686 25888 33692 25900
rect 32999 25860 33692 25888
rect 32999 25857 33011 25860
rect 32953 25851 33011 25857
rect 33686 25848 33692 25860
rect 33744 25848 33750 25900
rect 33962 25888 33968 25900
rect 33923 25860 33968 25888
rect 33962 25848 33968 25860
rect 34020 25848 34026 25900
rect 34256 25897 34284 25928
rect 34149 25891 34207 25897
rect 34149 25857 34161 25891
rect 34195 25857 34207 25891
rect 34149 25851 34207 25857
rect 34241 25891 34299 25897
rect 34241 25857 34253 25891
rect 34287 25857 34299 25891
rect 34241 25851 34299 25857
rect 33042 25820 33048 25832
rect 31220 25792 31754 25820
rect 33003 25792 33048 25820
rect 27488 25780 27494 25792
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 28166 25752 28172 25764
rect 24084 25724 26188 25752
rect 26344 25724 28172 25752
rect 24084 25712 24090 25724
rect 23474 25684 23480 25696
rect 22848 25656 23480 25684
rect 23474 25644 23480 25656
rect 23532 25644 23538 25696
rect 24854 25644 24860 25696
rect 24912 25684 24918 25696
rect 26344 25684 26372 25724
rect 28166 25712 28172 25724
rect 28224 25712 28230 25764
rect 30561 25755 30619 25761
rect 30561 25721 30573 25755
rect 30607 25752 30619 25755
rect 31662 25752 31668 25764
rect 30607 25724 31668 25752
rect 30607 25721 30619 25724
rect 30561 25715 30619 25721
rect 31662 25712 31668 25724
rect 31720 25712 31726 25764
rect 32214 25712 32220 25764
rect 32272 25752 32278 25764
rect 32490 25752 32496 25764
rect 32272 25724 32496 25752
rect 32272 25712 32278 25724
rect 32490 25712 32496 25724
rect 32548 25752 32554 25764
rect 34164 25752 34192 25851
rect 32548 25724 34192 25752
rect 32548 25712 32554 25724
rect 24912 25656 26372 25684
rect 26421 25687 26479 25693
rect 24912 25644 24918 25656
rect 26421 25653 26433 25687
rect 26467 25684 26479 25687
rect 26878 25684 26884 25696
rect 26467 25656 26884 25684
rect 26467 25653 26479 25656
rect 26421 25647 26479 25653
rect 26878 25644 26884 25656
rect 26936 25644 26942 25696
rect 28353 25687 28411 25693
rect 28353 25653 28365 25687
rect 28399 25684 28411 25687
rect 29546 25684 29552 25696
rect 28399 25656 29552 25684
rect 28399 25653 28411 25656
rect 28353 25647 28411 25653
rect 29546 25644 29552 25656
rect 29604 25644 29610 25696
rect 33318 25644 33324 25696
rect 33376 25684 33382 25696
rect 33781 25687 33839 25693
rect 33781 25684 33793 25687
rect 33376 25656 33793 25684
rect 33376 25644 33382 25656
rect 33781 25653 33793 25656
rect 33827 25653 33839 25687
rect 33781 25647 33839 25653
rect 46290 25644 46296 25696
rect 46348 25684 46354 25696
rect 47765 25687 47823 25693
rect 47765 25684 47777 25687
rect 46348 25656 47777 25684
rect 46348 25644 46354 25656
rect 47765 25653 47777 25656
rect 47811 25653 47823 25687
rect 47765 25647 47823 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 15562 25480 15568 25492
rect 15396 25452 15568 25480
rect 15396 25421 15424 25452
rect 15562 25440 15568 25452
rect 15620 25480 15626 25492
rect 17402 25480 17408 25492
rect 15620 25452 17408 25480
rect 15620 25440 15626 25452
rect 17402 25440 17408 25452
rect 17460 25480 17466 25492
rect 18417 25483 18475 25489
rect 18417 25480 18429 25483
rect 17460 25452 18429 25480
rect 17460 25440 17466 25452
rect 18417 25449 18429 25452
rect 18463 25449 18475 25483
rect 19334 25480 19340 25492
rect 19295 25452 19340 25480
rect 18417 25443 18475 25449
rect 19334 25440 19340 25452
rect 19392 25440 19398 25492
rect 23014 25480 23020 25492
rect 22975 25452 23020 25480
rect 23014 25440 23020 25452
rect 23072 25440 23078 25492
rect 24486 25480 24492 25492
rect 24447 25452 24492 25480
rect 24486 25440 24492 25452
rect 24544 25440 24550 25492
rect 24964 25452 31754 25480
rect 15381 25415 15439 25421
rect 15381 25381 15393 25415
rect 15427 25381 15439 25415
rect 15381 25375 15439 25381
rect 21542 25372 21548 25424
rect 21600 25412 21606 25424
rect 21910 25412 21916 25424
rect 21600 25384 21916 25412
rect 21600 25372 21606 25384
rect 21910 25372 21916 25384
rect 21968 25372 21974 25424
rect 22830 25372 22836 25424
rect 22888 25412 22894 25424
rect 23385 25415 23443 25421
rect 23385 25412 23397 25415
rect 22888 25384 23397 25412
rect 22888 25372 22894 25384
rect 23385 25381 23397 25384
rect 23431 25381 23443 25415
rect 23385 25375 23443 25381
rect 10226 25344 10232 25356
rect 10187 25316 10232 25344
rect 10226 25304 10232 25316
rect 10284 25304 10290 25356
rect 10502 25344 10508 25356
rect 10463 25316 10508 25344
rect 10502 25304 10508 25316
rect 10560 25304 10566 25356
rect 11790 25304 11796 25356
rect 11848 25344 11854 25356
rect 12253 25347 12311 25353
rect 12253 25344 12265 25347
rect 11848 25316 12265 25344
rect 11848 25304 11854 25316
rect 12253 25313 12265 25316
rect 12299 25313 12311 25347
rect 12253 25307 12311 25313
rect 15470 25304 15476 25356
rect 15528 25344 15534 25356
rect 16942 25344 16948 25356
rect 15528 25316 15884 25344
rect 16903 25316 16948 25344
rect 15528 25304 15534 25316
rect 11606 25236 11612 25288
rect 11664 25236 11670 25288
rect 14734 25276 14740 25288
rect 14695 25248 14740 25276
rect 14734 25236 14740 25248
rect 14792 25236 14798 25288
rect 14826 25236 14832 25288
rect 14884 25276 14890 25288
rect 15749 25279 15807 25285
rect 15749 25276 15761 25279
rect 14884 25248 15761 25276
rect 14884 25236 14890 25248
rect 15749 25245 15761 25248
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 14090 25168 14096 25220
rect 14148 25208 14154 25220
rect 14369 25211 14427 25217
rect 14369 25208 14381 25211
rect 14148 25180 14381 25208
rect 14148 25168 14154 25180
rect 14369 25177 14381 25180
rect 14415 25177 14427 25211
rect 14369 25171 14427 25177
rect 14553 25211 14611 25217
rect 14553 25177 14565 25211
rect 14599 25208 14611 25211
rect 15010 25208 15016 25220
rect 14599 25180 15016 25208
rect 14599 25177 14611 25180
rect 14553 25171 14611 25177
rect 15010 25168 15016 25180
rect 15068 25168 15074 25220
rect 15102 25168 15108 25220
rect 15160 25208 15166 25220
rect 15657 25211 15715 25217
rect 15657 25208 15669 25211
rect 15160 25180 15332 25208
rect 15160 25168 15166 25180
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 2038 25140 2044 25152
rect 1995 25112 2044 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 14645 25143 14703 25149
rect 14645 25109 14657 25143
rect 14691 25140 14703 25143
rect 14826 25140 14832 25152
rect 14691 25112 14832 25140
rect 14691 25109 14703 25112
rect 14645 25103 14703 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 14921 25143 14979 25149
rect 14921 25109 14933 25143
rect 14967 25140 14979 25143
rect 15194 25140 15200 25152
rect 14967 25112 15200 25140
rect 14967 25109 14979 25112
rect 14921 25103 14979 25109
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 15304 25140 15332 25180
rect 15488 25180 15669 25208
rect 15488 25140 15516 25180
rect 15657 25177 15669 25180
rect 15703 25177 15715 25211
rect 15856 25208 15884 25316
rect 16942 25304 16948 25316
rect 17000 25304 17006 25356
rect 19518 25304 19524 25356
rect 19576 25344 19582 25356
rect 20257 25347 20315 25353
rect 20257 25344 20269 25347
rect 19576 25316 20269 25344
rect 19576 25304 19582 25316
rect 20257 25313 20269 25316
rect 20303 25344 20315 25347
rect 24854 25344 24860 25356
rect 20303 25316 24860 25344
rect 20303 25313 20315 25316
rect 20257 25307 20315 25313
rect 24854 25304 24860 25316
rect 24912 25304 24918 25356
rect 16666 25276 16672 25288
rect 16627 25248 16672 25276
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 19242 25276 19248 25288
rect 18288 25248 19248 25276
rect 18288 25236 18294 25248
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 20441 25279 20499 25285
rect 20441 25245 20453 25279
rect 20487 25245 20499 25279
rect 20441 25239 20499 25245
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25276 20683 25279
rect 21177 25279 21235 25285
rect 21177 25276 21189 25279
rect 20671 25248 21189 25276
rect 20671 25245 20683 25248
rect 20625 25239 20683 25245
rect 21177 25245 21189 25248
rect 21223 25245 21235 25279
rect 21177 25239 21235 25245
rect 18322 25208 18328 25220
rect 15856 25180 17172 25208
rect 18170 25180 18328 25208
rect 15657 25171 15715 25177
rect 15304 25112 15516 25140
rect 15565 25143 15623 25149
rect 15565 25109 15577 25143
rect 15611 25140 15623 25143
rect 15838 25140 15844 25152
rect 15611 25112 15844 25140
rect 15611 25109 15623 25112
rect 15565 25103 15623 25109
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 15933 25143 15991 25149
rect 15933 25109 15945 25143
rect 15979 25140 15991 25143
rect 16574 25140 16580 25152
rect 15979 25112 16580 25140
rect 15979 25109 15991 25112
rect 15933 25103 15991 25109
rect 16574 25100 16580 25112
rect 16632 25140 16638 25152
rect 17034 25140 17040 25152
rect 16632 25112 17040 25140
rect 16632 25100 16638 25112
rect 17034 25100 17040 25112
rect 17092 25100 17098 25152
rect 17144 25140 17172 25180
rect 18322 25168 18328 25180
rect 18380 25168 18386 25220
rect 20456 25140 20484 25239
rect 21266 25236 21272 25288
rect 21324 25276 21330 25288
rect 21542 25276 21548 25288
rect 21324 25248 21369 25276
rect 21503 25248 21548 25276
rect 21324 25236 21330 25248
rect 21542 25236 21548 25248
rect 21600 25236 21606 25288
rect 21683 25279 21741 25285
rect 21683 25245 21695 25279
rect 21729 25276 21741 25279
rect 22002 25276 22008 25288
rect 21729 25248 22008 25276
rect 21729 25245 21741 25248
rect 21683 25239 21741 25245
rect 22002 25236 22008 25248
rect 22060 25236 22066 25288
rect 23017 25279 23075 25285
rect 23017 25245 23029 25279
rect 23063 25276 23075 25279
rect 23106 25276 23112 25288
rect 23063 25248 23112 25276
rect 23063 25245 23075 25248
rect 23017 25239 23075 25245
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25276 23259 25279
rect 23842 25276 23848 25288
rect 23247 25248 23848 25276
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 23842 25236 23848 25248
rect 23900 25236 23906 25288
rect 24394 25276 24400 25288
rect 24355 25248 24400 25276
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 21082 25168 21088 25220
rect 21140 25208 21146 25220
rect 21453 25211 21511 25217
rect 21453 25208 21465 25211
rect 21140 25180 21465 25208
rect 21140 25168 21146 25180
rect 21453 25177 21465 25180
rect 21499 25177 21511 25211
rect 24964 25208 24992 25452
rect 26234 25412 26240 25424
rect 25424 25384 26240 25412
rect 25424 25285 25452 25384
rect 26234 25372 26240 25384
rect 26292 25372 26298 25424
rect 29270 25372 29276 25424
rect 29328 25412 29334 25424
rect 29733 25415 29791 25421
rect 29733 25412 29745 25415
rect 29328 25384 29745 25412
rect 29328 25372 29334 25384
rect 29733 25381 29745 25384
rect 29779 25381 29791 25415
rect 31726 25412 31754 25452
rect 33686 25440 33692 25492
rect 33744 25480 33750 25492
rect 34149 25483 34207 25489
rect 34149 25480 34161 25483
rect 33744 25452 34161 25480
rect 33744 25440 33750 25452
rect 34149 25449 34161 25452
rect 34195 25449 34207 25483
rect 34149 25443 34207 25449
rect 32214 25412 32220 25424
rect 31726 25384 32220 25412
rect 29733 25375 29791 25381
rect 32214 25372 32220 25384
rect 32272 25372 32278 25424
rect 25866 25304 25872 25356
rect 25924 25344 25930 25356
rect 28626 25344 28632 25356
rect 25924 25316 28632 25344
rect 25924 25304 25930 25316
rect 28626 25304 28632 25316
rect 28684 25304 28690 25356
rect 31386 25344 31392 25356
rect 30760 25316 31392 25344
rect 25409 25279 25467 25285
rect 25409 25245 25421 25279
rect 25455 25245 25467 25279
rect 25590 25276 25596 25288
rect 25551 25248 25596 25276
rect 25409 25239 25467 25245
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 25774 25276 25780 25288
rect 25735 25248 25780 25276
rect 25774 25236 25780 25248
rect 25832 25236 25838 25288
rect 26602 25276 26608 25288
rect 26563 25248 26608 25276
rect 26602 25236 26608 25248
rect 26660 25236 26666 25288
rect 26697 25279 26755 25285
rect 26697 25245 26709 25279
rect 26743 25245 26755 25279
rect 26878 25276 26884 25288
rect 26839 25248 26884 25276
rect 26697 25239 26755 25245
rect 21453 25171 21511 25177
rect 21652 25180 24992 25208
rect 25685 25211 25743 25217
rect 17144 25112 20484 25140
rect 21468 25140 21496 25171
rect 21652 25140 21680 25180
rect 25685 25177 25697 25211
rect 25731 25208 25743 25211
rect 26712 25208 26740 25239
rect 26878 25236 26884 25248
rect 26936 25236 26942 25288
rect 26970 25236 26976 25288
rect 27028 25276 27034 25288
rect 29546 25276 29552 25288
rect 27028 25248 27073 25276
rect 29507 25248 29552 25276
rect 27028 25236 27034 25248
rect 29546 25236 29552 25248
rect 29604 25236 29610 25288
rect 30760 25285 30788 25316
rect 31386 25304 31392 25316
rect 31444 25344 31450 25356
rect 31444 25316 31754 25344
rect 31444 25304 31450 25316
rect 30745 25279 30803 25285
rect 30745 25245 30757 25279
rect 30791 25245 30803 25279
rect 31110 25276 31116 25288
rect 31071 25248 31116 25276
rect 30745 25239 30803 25245
rect 31110 25236 31116 25248
rect 31168 25236 31174 25288
rect 27522 25208 27528 25220
rect 25731 25180 27528 25208
rect 25731 25177 25743 25180
rect 25685 25171 25743 25177
rect 27522 25168 27528 25180
rect 27580 25168 27586 25220
rect 29564 25208 29592 25236
rect 30929 25211 30987 25217
rect 30929 25208 30941 25211
rect 29564 25180 30941 25208
rect 30929 25177 30941 25180
rect 30975 25177 30987 25211
rect 30929 25171 30987 25177
rect 31021 25211 31079 25217
rect 31021 25177 31033 25211
rect 31067 25177 31079 25211
rect 31726 25208 31754 25316
rect 32306 25304 32312 25356
rect 32364 25344 32370 25356
rect 32401 25347 32459 25353
rect 32401 25344 32413 25347
rect 32364 25316 32413 25344
rect 32364 25304 32370 25316
rect 32401 25313 32413 25316
rect 32447 25313 32459 25347
rect 32401 25307 32459 25313
rect 32677 25347 32735 25353
rect 32677 25313 32689 25347
rect 32723 25344 32735 25347
rect 33318 25344 33324 25356
rect 32723 25316 33324 25344
rect 32723 25313 32735 25316
rect 32677 25307 32735 25313
rect 33318 25304 33324 25316
rect 33376 25304 33382 25356
rect 46290 25344 46296 25356
rect 46251 25316 46296 25344
rect 46290 25304 46296 25316
rect 46348 25304 46354 25356
rect 32582 25208 32588 25220
rect 31726 25180 32588 25208
rect 31021 25171 31079 25177
rect 21468 25112 21680 25140
rect 21821 25143 21879 25149
rect 21821 25109 21833 25143
rect 21867 25140 21879 25143
rect 22094 25140 22100 25152
rect 21867 25112 22100 25140
rect 21867 25109 21879 25112
rect 21821 25103 21879 25109
rect 22094 25100 22100 25112
rect 22152 25100 22158 25152
rect 25406 25100 25412 25152
rect 25464 25140 25470 25152
rect 25961 25143 26019 25149
rect 25961 25140 25973 25143
rect 25464 25112 25973 25140
rect 25464 25100 25470 25112
rect 25961 25109 25973 25112
rect 26007 25109 26019 25143
rect 25961 25103 26019 25109
rect 26234 25100 26240 25152
rect 26292 25140 26298 25152
rect 26421 25143 26479 25149
rect 26421 25140 26433 25143
rect 26292 25112 26433 25140
rect 26292 25100 26298 25112
rect 26421 25109 26433 25112
rect 26467 25109 26479 25143
rect 26421 25103 26479 25109
rect 30834 25100 30840 25152
rect 30892 25140 30898 25152
rect 31036 25140 31064 25171
rect 32582 25168 32588 25180
rect 32640 25168 32646 25220
rect 33134 25168 33140 25220
rect 33192 25168 33198 25220
rect 35158 25208 35164 25220
rect 35119 25180 35164 25208
rect 35158 25168 35164 25180
rect 35216 25168 35222 25220
rect 46477 25211 46535 25217
rect 46477 25177 46489 25211
rect 46523 25208 46535 25211
rect 47670 25208 47676 25220
rect 46523 25180 47676 25208
rect 46523 25177 46535 25180
rect 46477 25171 46535 25177
rect 47670 25168 47676 25180
rect 47728 25168 47734 25220
rect 48130 25208 48136 25220
rect 48091 25180 48136 25208
rect 48130 25168 48136 25180
rect 48188 25168 48194 25220
rect 31294 25140 31300 25152
rect 30892 25112 31064 25140
rect 31255 25112 31300 25140
rect 30892 25100 30898 25112
rect 31294 25100 31300 25112
rect 31352 25100 31358 25152
rect 34790 25100 34796 25152
rect 34848 25140 34854 25152
rect 35253 25143 35311 25149
rect 35253 25140 35265 25143
rect 34848 25112 35265 25140
rect 34848 25100 34854 25112
rect 35253 25109 35265 25112
rect 35299 25109 35311 25143
rect 35253 25103 35311 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 14734 24896 14740 24948
rect 14792 24936 14798 24948
rect 14921 24939 14979 24945
rect 14921 24936 14933 24939
rect 14792 24908 14933 24936
rect 14792 24896 14798 24908
rect 14921 24905 14933 24908
rect 14967 24905 14979 24939
rect 14921 24899 14979 24905
rect 15473 24939 15531 24945
rect 15473 24905 15485 24939
rect 15519 24936 15531 24939
rect 15654 24936 15660 24948
rect 15519 24908 15660 24936
rect 15519 24905 15531 24908
rect 15473 24899 15531 24905
rect 15654 24896 15660 24908
rect 15712 24896 15718 24948
rect 17034 24936 17040 24948
rect 16995 24908 17040 24936
rect 17034 24896 17040 24908
rect 17092 24896 17098 24948
rect 21266 24936 21272 24948
rect 21227 24908 21272 24936
rect 21266 24896 21272 24908
rect 21324 24896 21330 24948
rect 23474 24936 23480 24948
rect 22066 24908 23480 24936
rect 16853 24871 16911 24877
rect 16853 24868 16865 24871
rect 14568 24840 16865 24868
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10962 24800 10968 24812
rect 10923 24772 10968 24800
rect 10781 24763 10839 24769
rect 10796 24732 10824 24763
rect 10962 24760 10968 24772
rect 11020 24760 11026 24812
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 11330 24732 11336 24744
rect 10796 24704 11336 24732
rect 11330 24692 11336 24704
rect 11388 24692 11394 24744
rect 11532 24732 11560 24763
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11664 24772 11709 24800
rect 11664 24760 11670 24772
rect 14568 24744 14596 24840
rect 16853 24837 16865 24840
rect 16899 24837 16911 24871
rect 16853 24831 16911 24837
rect 16942 24828 16948 24880
rect 17000 24868 17006 24880
rect 22066 24868 22094 24908
rect 23474 24896 23480 24908
rect 23532 24936 23538 24948
rect 24670 24936 24676 24948
rect 23532 24908 24676 24936
rect 23532 24896 23538 24908
rect 24670 24896 24676 24908
rect 24728 24896 24734 24948
rect 25038 24896 25044 24948
rect 25096 24936 25102 24948
rect 25774 24936 25780 24948
rect 25096 24908 25780 24936
rect 25096 24896 25102 24908
rect 25774 24896 25780 24908
rect 25832 24896 25838 24948
rect 26421 24939 26479 24945
rect 26421 24905 26433 24939
rect 26467 24936 26479 24939
rect 26510 24936 26516 24948
rect 26467 24908 26516 24936
rect 26467 24905 26479 24908
rect 26421 24899 26479 24905
rect 26510 24896 26516 24908
rect 26568 24896 26574 24948
rect 17000 24840 17045 24868
rect 21836 24840 22094 24868
rect 31021 24871 31079 24877
rect 17000 24828 17006 24840
rect 14734 24800 14740 24812
rect 14695 24772 14740 24800
rect 14734 24760 14740 24772
rect 14792 24760 14798 24812
rect 15562 24760 15568 24812
rect 15620 24800 15626 24812
rect 15657 24803 15715 24809
rect 15657 24800 15669 24803
rect 15620 24772 15669 24800
rect 15620 24760 15626 24772
rect 15657 24769 15669 24772
rect 15703 24769 15715 24803
rect 15838 24800 15844 24812
rect 15799 24772 15844 24800
rect 15657 24763 15715 24769
rect 15838 24760 15844 24772
rect 15896 24760 15902 24812
rect 15933 24803 15991 24809
rect 15933 24769 15945 24803
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24800 16727 24803
rect 16758 24800 16764 24812
rect 16715 24772 16764 24800
rect 16715 24769 16727 24772
rect 16669 24763 16727 24769
rect 12342 24732 12348 24744
rect 11532 24704 12348 24732
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 14550 24732 14556 24744
rect 14511 24704 14556 24732
rect 14550 24692 14556 24704
rect 14608 24692 14614 24744
rect 15194 24692 15200 24744
rect 15252 24732 15258 24744
rect 15948 24732 15976 24763
rect 16758 24760 16764 24772
rect 16816 24760 16822 24812
rect 18230 24800 18236 24812
rect 18191 24772 18236 24800
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 20901 24803 20959 24809
rect 18380 24772 18425 24800
rect 18380 24760 18386 24772
rect 20901 24769 20913 24803
rect 20947 24800 20959 24803
rect 21542 24800 21548 24812
rect 20947 24772 21548 24800
rect 20947 24769 20959 24772
rect 20901 24763 20959 24769
rect 21542 24760 21548 24772
rect 21600 24760 21606 24812
rect 21836 24809 21864 24840
rect 31021 24837 31033 24871
rect 31067 24868 31079 24871
rect 31294 24868 31300 24880
rect 31067 24840 31300 24868
rect 31067 24837 31079 24840
rect 31021 24831 31079 24837
rect 31294 24828 31300 24840
rect 31352 24828 31358 24880
rect 34790 24828 34796 24880
rect 34848 24868 34854 24880
rect 34848 24840 35848 24868
rect 34848 24828 34854 24840
rect 21821 24803 21879 24809
rect 21821 24769 21833 24803
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 23198 24760 23204 24812
rect 23256 24760 23262 24812
rect 26970 24800 26976 24812
rect 15252 24704 15976 24732
rect 17221 24735 17279 24741
rect 15252 24692 15258 24704
rect 17221 24701 17233 24735
rect 17267 24732 17279 24735
rect 20714 24732 20720 24744
rect 17267 24704 20720 24732
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 20714 24692 20720 24704
rect 20772 24692 20778 24744
rect 20990 24732 20996 24744
rect 20951 24704 20996 24732
rect 20990 24692 20996 24704
rect 21048 24692 21054 24744
rect 22094 24692 22100 24744
rect 22152 24732 22158 24744
rect 24670 24732 24676 24744
rect 22152 24704 22197 24732
rect 24631 24704 24676 24732
rect 22152 24692 22158 24704
rect 24670 24692 24676 24704
rect 24728 24692 24734 24744
rect 24949 24735 25007 24741
rect 24949 24701 24961 24735
rect 24995 24732 25007 24735
rect 26068 24732 26096 24786
rect 26931 24772 26976 24800
rect 26970 24760 26976 24772
rect 27028 24760 27034 24812
rect 28074 24800 28080 24812
rect 28035 24772 28080 24800
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 29638 24800 29644 24812
rect 29486 24772 29644 24800
rect 29638 24760 29644 24772
rect 29696 24760 29702 24812
rect 30561 24803 30619 24809
rect 30561 24769 30573 24803
rect 30607 24769 30619 24803
rect 31202 24800 31208 24812
rect 31163 24772 31208 24800
rect 30561 24763 30619 24769
rect 27065 24735 27123 24741
rect 27065 24732 27077 24735
rect 24995 24704 26004 24732
rect 26068 24704 27077 24732
rect 24995 24701 25007 24704
rect 24949 24695 25007 24701
rect 25976 24664 26004 24704
rect 27065 24701 27077 24704
rect 27111 24701 27123 24735
rect 28350 24732 28356 24744
rect 28311 24704 28356 24732
rect 27065 24695 27123 24701
rect 28350 24692 28356 24704
rect 28408 24692 28414 24744
rect 29825 24735 29883 24741
rect 29825 24701 29837 24735
rect 29871 24732 29883 24735
rect 30374 24732 30380 24744
rect 29871 24704 30380 24732
rect 29871 24701 29883 24704
rect 29825 24695 29883 24701
rect 30374 24692 30380 24704
rect 30432 24692 30438 24744
rect 30576 24732 30604 24763
rect 31202 24760 31208 24772
rect 31260 24760 31266 24812
rect 32214 24800 32220 24812
rect 32175 24772 32220 24800
rect 32214 24760 32220 24772
rect 32272 24760 32278 24812
rect 32398 24800 32404 24812
rect 32359 24772 32404 24800
rect 32398 24760 32404 24772
rect 32456 24760 32462 24812
rect 32490 24760 32496 24812
rect 32548 24800 32554 24812
rect 32861 24803 32919 24809
rect 32861 24800 32873 24803
rect 32548 24772 32873 24800
rect 32548 24760 32554 24772
rect 32861 24769 32873 24772
rect 32907 24769 32919 24803
rect 32861 24763 32919 24769
rect 32953 24803 33011 24809
rect 32953 24769 32965 24803
rect 32999 24800 33011 24803
rect 33134 24800 33140 24812
rect 32999 24772 33140 24800
rect 32999 24769 33011 24772
rect 32953 24763 33011 24769
rect 33134 24760 33140 24772
rect 33192 24760 33198 24812
rect 35158 24800 35164 24812
rect 35119 24772 35164 24800
rect 35158 24760 35164 24772
rect 35216 24760 35222 24812
rect 35820 24800 35848 24840
rect 39945 24803 40003 24809
rect 39945 24800 39957 24803
rect 35820 24772 39957 24800
rect 39945 24769 39957 24772
rect 39991 24800 40003 24803
rect 45002 24800 45008 24812
rect 39991 24772 45008 24800
rect 39991 24769 40003 24772
rect 39945 24763 40003 24769
rect 45002 24760 45008 24772
rect 45060 24760 45066 24812
rect 47578 24800 47584 24812
rect 47539 24772 47584 24800
rect 47578 24760 47584 24772
rect 47636 24760 47642 24812
rect 47670 24760 47676 24812
rect 47728 24800 47734 24812
rect 47728 24772 47773 24800
rect 47728 24760 47734 24772
rect 31389 24735 31447 24741
rect 31389 24732 31401 24735
rect 30576 24704 31401 24732
rect 31389 24701 31401 24704
rect 31435 24701 31447 24735
rect 31389 24695 31447 24701
rect 32122 24692 32128 24744
rect 32180 24732 32186 24744
rect 35437 24735 35495 24741
rect 35437 24732 35449 24735
rect 32180 24704 35449 24732
rect 32180 24692 32186 24704
rect 35437 24701 35449 24704
rect 35483 24732 35495 24735
rect 44358 24732 44364 24744
rect 35483 24704 44364 24732
rect 35483 24701 35495 24704
rect 35437 24695 35495 24701
rect 44358 24692 44364 24704
rect 44416 24692 44422 24744
rect 45094 24692 45100 24744
rect 45152 24732 45158 24744
rect 45189 24735 45247 24741
rect 45189 24732 45201 24735
rect 45152 24704 45201 24732
rect 45152 24692 45158 24704
rect 45189 24701 45201 24704
rect 45235 24701 45247 24735
rect 45370 24732 45376 24744
rect 45331 24704 45376 24732
rect 45189 24695 45247 24701
rect 45370 24692 45376 24704
rect 45428 24692 45434 24744
rect 46750 24732 46756 24744
rect 46711 24704 46756 24732
rect 46750 24692 46756 24704
rect 46808 24692 46814 24744
rect 26234 24664 26240 24676
rect 25976 24636 26240 24664
rect 26234 24624 26240 24636
rect 26292 24624 26298 24676
rect 46842 24664 46848 24676
rect 29564 24636 46848 24664
rect 10594 24556 10600 24608
rect 10652 24596 10658 24608
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 10652 24568 10793 24596
rect 10652 24556 10658 24568
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 10781 24559 10839 24565
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 23569 24599 23627 24605
rect 23569 24596 23581 24599
rect 21968 24568 23581 24596
rect 21968 24556 21974 24568
rect 23569 24565 23581 24568
rect 23615 24565 23627 24599
rect 23569 24559 23627 24565
rect 27338 24556 27344 24608
rect 27396 24596 27402 24608
rect 29564 24596 29592 24636
rect 46842 24624 46848 24636
rect 46900 24624 46906 24676
rect 30374 24596 30380 24608
rect 27396 24568 29592 24596
rect 30335 24568 30380 24596
rect 27396 24556 27402 24568
rect 30374 24556 30380 24568
rect 30432 24556 30438 24608
rect 30650 24556 30656 24608
rect 30708 24596 30714 24608
rect 32122 24596 32128 24608
rect 30708 24568 32128 24596
rect 30708 24556 30714 24568
rect 32122 24556 32128 24568
rect 32180 24556 32186 24608
rect 32214 24556 32220 24608
rect 32272 24596 32278 24608
rect 34790 24596 34796 24608
rect 32272 24568 34796 24596
rect 32272 24556 32278 24568
rect 34790 24556 34796 24568
rect 34848 24556 34854 24608
rect 40034 24596 40040 24608
rect 39995 24568 40040 24596
rect 40034 24556 40040 24568
rect 40092 24556 40098 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 16577 24395 16635 24401
rect 16577 24361 16589 24395
rect 16623 24392 16635 24395
rect 16666 24392 16672 24404
rect 16623 24364 16672 24392
rect 16623 24361 16635 24364
rect 16577 24355 16635 24361
rect 16666 24352 16672 24364
rect 16724 24352 16730 24404
rect 19334 24352 19340 24404
rect 19392 24392 19398 24404
rect 23106 24392 23112 24404
rect 19392 24364 23112 24392
rect 19392 24352 19398 24364
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 23198 24352 23204 24404
rect 23256 24392 23262 24404
rect 23293 24395 23351 24401
rect 23293 24392 23305 24395
rect 23256 24364 23305 24392
rect 23256 24352 23262 24364
rect 23293 24361 23305 24364
rect 23339 24361 23351 24395
rect 23293 24355 23351 24361
rect 26050 24352 26056 24404
rect 26108 24392 26114 24404
rect 26881 24395 26939 24401
rect 26108 24364 26464 24392
rect 26108 24352 26114 24364
rect 19429 24327 19487 24333
rect 19429 24324 19441 24327
rect 17696 24296 19441 24324
rect 10594 24256 10600 24268
rect 10555 24228 10600 24256
rect 10594 24216 10600 24228
rect 10652 24216 10658 24268
rect 10318 24188 10324 24200
rect 10279 24160 10324 24188
rect 10318 24148 10324 24160
rect 10376 24148 10382 24200
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12400 24160 12541 24188
rect 12400 24148 12406 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 14918 24148 14924 24200
rect 14976 24188 14982 24200
rect 16485 24191 16543 24197
rect 16485 24188 16497 24191
rect 14976 24160 16497 24188
rect 14976 24148 14982 24160
rect 16485 24157 16497 24160
rect 16531 24188 16543 24191
rect 16850 24188 16856 24200
rect 16531 24160 16856 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 17696 24197 17724 24296
rect 19429 24293 19441 24296
rect 19475 24324 19487 24327
rect 20530 24324 20536 24336
rect 19475 24296 20536 24324
rect 19475 24293 19487 24296
rect 19429 24287 19487 24293
rect 20530 24284 20536 24296
rect 20588 24284 20594 24336
rect 26436 24324 26464 24364
rect 26881 24361 26893 24395
rect 26927 24392 26939 24395
rect 27154 24392 27160 24404
rect 26927 24364 27160 24392
rect 26927 24361 26939 24364
rect 26881 24355 26939 24361
rect 27154 24352 27160 24364
rect 27212 24352 27218 24404
rect 29638 24392 29644 24404
rect 29599 24364 29644 24392
rect 29638 24352 29644 24364
rect 29696 24352 29702 24404
rect 30374 24352 30380 24404
rect 30432 24392 30438 24404
rect 31002 24395 31060 24401
rect 31002 24392 31014 24395
rect 30432 24364 31014 24392
rect 30432 24352 30438 24364
rect 31002 24361 31014 24364
rect 31048 24361 31060 24395
rect 31002 24355 31060 24361
rect 32493 24395 32551 24401
rect 32493 24361 32505 24395
rect 32539 24392 32551 24395
rect 32582 24392 32588 24404
rect 32539 24364 32588 24392
rect 32539 24361 32551 24364
rect 32493 24355 32551 24361
rect 32582 24352 32588 24364
rect 32640 24352 32646 24404
rect 45097 24395 45155 24401
rect 45097 24361 45109 24395
rect 45143 24392 45155 24395
rect 45370 24392 45376 24404
rect 45143 24364 45376 24392
rect 45143 24361 45155 24364
rect 45097 24355 45155 24361
rect 45370 24352 45376 24364
rect 45428 24352 45434 24404
rect 30650 24324 30656 24336
rect 26436 24296 30656 24324
rect 30650 24284 30656 24296
rect 30708 24284 30714 24336
rect 45646 24324 45652 24336
rect 36924 24296 45652 24324
rect 17770 24216 17776 24268
rect 17828 24256 17834 24268
rect 17828 24228 20024 24256
rect 17828 24216 17834 24228
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 19058 24148 19064 24200
rect 19116 24188 19122 24200
rect 19996 24197 20024 24228
rect 24670 24216 24676 24268
rect 24728 24256 24734 24268
rect 25133 24259 25191 24265
rect 25133 24256 25145 24259
rect 24728 24228 25145 24256
rect 24728 24216 24734 24228
rect 25133 24225 25145 24228
rect 25179 24225 25191 24259
rect 25406 24256 25412 24268
rect 25367 24228 25412 24256
rect 25133 24219 25191 24225
rect 25406 24216 25412 24228
rect 25464 24216 25470 24268
rect 30745 24259 30803 24265
rect 30745 24225 30757 24259
rect 30791 24256 30803 24259
rect 32306 24256 32312 24268
rect 30791 24228 32312 24256
rect 30791 24225 30803 24228
rect 30745 24219 30803 24225
rect 32306 24216 32312 24228
rect 32364 24216 32370 24268
rect 34149 24259 34207 24265
rect 34149 24225 34161 24259
rect 34195 24256 34207 24259
rect 35342 24256 35348 24268
rect 34195 24228 35348 24256
rect 34195 24225 34207 24228
rect 34149 24219 34207 24225
rect 35342 24216 35348 24228
rect 35400 24216 35406 24268
rect 36924 24265 36952 24296
rect 45646 24284 45652 24296
rect 45704 24284 45710 24336
rect 36909 24259 36967 24265
rect 36909 24225 36921 24259
rect 36955 24225 36967 24259
rect 40034 24256 40040 24268
rect 39995 24228 40040 24256
rect 36909 24219 36967 24225
rect 40034 24216 40040 24228
rect 40092 24216 40098 24268
rect 40310 24256 40316 24268
rect 40271 24228 40316 24256
rect 40310 24216 40316 24228
rect 40368 24216 40374 24268
rect 44358 24216 44364 24268
rect 44416 24256 44422 24268
rect 44416 24228 45692 24256
rect 44416 24216 44422 24228
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 19116 24160 19257 24188
rect 19116 24148 19122 24160
rect 19245 24157 19257 24160
rect 19291 24157 19303 24191
rect 19245 24151 19303 24157
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24188 20039 24191
rect 22830 24188 22836 24200
rect 20027 24160 22836 24188
rect 20027 24157 20039 24160
rect 19981 24151 20039 24157
rect 12621 24123 12679 24129
rect 12621 24120 12633 24123
rect 11822 24092 12633 24120
rect 12621 24089 12633 24092
rect 12667 24089 12679 24123
rect 19260 24120 19288 24151
rect 22830 24148 22836 24160
rect 22888 24148 22894 24200
rect 23201 24191 23259 24197
rect 23201 24157 23213 24191
rect 23247 24188 23259 24191
rect 24394 24188 24400 24200
rect 23247 24160 24400 24188
rect 23247 24157 23259 24160
rect 23201 24151 23259 24157
rect 24394 24148 24400 24160
rect 24452 24148 24458 24200
rect 28626 24148 28632 24200
rect 28684 24188 28690 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 28684 24160 29561 24188
rect 28684 24148 28690 24160
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 29549 24151 29607 24157
rect 32122 24148 32128 24200
rect 32180 24148 32186 24200
rect 34606 24148 34612 24200
rect 34664 24188 34670 24200
rect 35069 24191 35127 24197
rect 35069 24188 35081 24191
rect 34664 24160 35081 24188
rect 34664 24148 34670 24160
rect 35069 24157 35081 24160
rect 35115 24157 35127 24191
rect 35069 24151 35127 24157
rect 39853 24191 39911 24197
rect 39853 24157 39865 24191
rect 39899 24157 39911 24191
rect 45002 24188 45008 24200
rect 44963 24160 45008 24188
rect 39853 24151 39911 24157
rect 19260 24092 22094 24120
rect 12621 24083 12679 24089
rect 11882 24012 11888 24064
rect 11940 24052 11946 24064
rect 12069 24055 12127 24061
rect 12069 24052 12081 24055
rect 11940 24024 12081 24052
rect 11940 24012 11946 24024
rect 12069 24021 12081 24024
rect 12115 24021 12127 24055
rect 12069 24015 12127 24021
rect 14366 24012 14372 24064
rect 14424 24052 14430 24064
rect 17678 24052 17684 24064
rect 14424 24024 17684 24052
rect 14424 24012 14430 24024
rect 17678 24012 17684 24024
rect 17736 24012 17742 24064
rect 17862 24052 17868 24064
rect 17823 24024 17868 24052
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 20070 24052 20076 24064
rect 20031 24024 20076 24052
rect 20070 24012 20076 24024
rect 20128 24012 20134 24064
rect 22066 24052 22094 24092
rect 25958 24080 25964 24132
rect 26016 24080 26022 24132
rect 33965 24123 34023 24129
rect 33965 24120 33977 24123
rect 26712 24092 27016 24120
rect 26712 24052 26740 24092
rect 22066 24024 26740 24052
rect 26988 24052 27016 24092
rect 32416 24092 33977 24120
rect 32416 24052 32444 24092
rect 33965 24089 33977 24092
rect 34011 24120 34023 24123
rect 34011 24092 34468 24120
rect 34011 24089 34023 24092
rect 33965 24083 34023 24089
rect 26988 24024 32444 24052
rect 34440 24052 34468 24092
rect 34514 24080 34520 24132
rect 34572 24120 34578 24132
rect 35253 24123 35311 24129
rect 35253 24120 35265 24123
rect 34572 24092 35265 24120
rect 34572 24080 34578 24092
rect 35253 24089 35265 24092
rect 35299 24089 35311 24123
rect 39868 24120 39896 24151
rect 45002 24148 45008 24160
rect 45060 24148 45066 24200
rect 45664 24197 45692 24228
rect 46474 24216 46480 24268
rect 46532 24256 46538 24268
rect 46937 24259 46995 24265
rect 46937 24256 46949 24259
rect 46532 24228 46949 24256
rect 46532 24216 46538 24228
rect 46937 24225 46949 24228
rect 46983 24225 46995 24259
rect 46937 24219 46995 24225
rect 45649 24191 45707 24197
rect 45649 24157 45661 24191
rect 45695 24188 45707 24191
rect 45830 24188 45836 24200
rect 45695 24160 45836 24188
rect 45695 24157 45707 24160
rect 45649 24151 45707 24157
rect 45830 24148 45836 24160
rect 45888 24148 45894 24200
rect 46290 24188 46296 24200
rect 46251 24160 46296 24188
rect 46290 24148 46296 24160
rect 46348 24148 46354 24200
rect 40034 24120 40040 24132
rect 39868 24092 40040 24120
rect 35253 24083 35311 24089
rect 40034 24080 40040 24092
rect 40092 24120 40098 24132
rect 41046 24120 41052 24132
rect 40092 24092 41052 24120
rect 40092 24080 40098 24092
rect 41046 24080 41052 24092
rect 41104 24080 41110 24132
rect 45741 24123 45799 24129
rect 41800 24092 45554 24120
rect 41800 24052 41828 24092
rect 34440 24024 41828 24052
rect 45526 24052 45554 24092
rect 45741 24089 45753 24123
rect 45787 24120 45799 24123
rect 46477 24123 46535 24129
rect 46477 24120 46489 24123
rect 45787 24092 46489 24120
rect 45787 24089 45799 24092
rect 45741 24083 45799 24089
rect 46477 24089 46489 24092
rect 46523 24089 46535 24123
rect 46477 24083 46535 24089
rect 47762 24052 47768 24064
rect 45526 24024 47768 24052
rect 47762 24012 47768 24024
rect 47820 24012 47826 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 17586 23848 17592 23860
rect 3568 23820 16896 23848
rect 17547 23820 17592 23848
rect 3568 23808 3574 23820
rect 3878 23740 3884 23792
rect 3936 23780 3942 23792
rect 3936 23752 10272 23780
rect 3936 23740 3942 23752
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 9950 23672 9956 23724
rect 10008 23712 10014 23724
rect 10137 23715 10195 23721
rect 10137 23712 10149 23715
rect 10008 23684 10149 23712
rect 10008 23672 10014 23684
rect 10137 23681 10149 23684
rect 10183 23681 10195 23715
rect 10244 23712 10272 23752
rect 10318 23740 10324 23792
rect 10376 23780 10382 23792
rect 10413 23783 10471 23789
rect 10413 23780 10425 23783
rect 10376 23752 10425 23780
rect 10376 23740 10382 23752
rect 10413 23749 10425 23752
rect 10459 23749 10471 23783
rect 14185 23783 14243 23789
rect 10413 23743 10471 23749
rect 10520 23752 13216 23780
rect 10520 23712 10548 23752
rect 10244 23684 10548 23712
rect 10137 23675 10195 23681
rect 11790 23644 11796 23656
rect 11751 23616 11796 23644
rect 11790 23604 11796 23616
rect 11848 23604 11854 23656
rect 11974 23644 11980 23656
rect 11935 23616 11980 23644
rect 11974 23604 11980 23616
rect 12032 23604 12038 23656
rect 13188 23653 13216 23752
rect 14185 23749 14197 23783
rect 14231 23780 14243 23783
rect 14366 23780 14372 23792
rect 14231 23752 14372 23780
rect 14231 23749 14243 23752
rect 14185 23743 14243 23749
rect 14366 23740 14372 23752
rect 14424 23740 14430 23792
rect 16868 23780 16896 23820
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 17678 23808 17684 23860
rect 17736 23848 17742 23860
rect 19334 23848 19340 23860
rect 17736 23820 19340 23848
rect 17736 23808 17742 23820
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 23474 23808 23480 23860
rect 23532 23848 23538 23860
rect 23753 23851 23811 23857
rect 23753 23848 23765 23851
rect 23532 23820 23765 23848
rect 23532 23808 23538 23820
rect 23753 23817 23765 23820
rect 23799 23848 23811 23851
rect 24394 23848 24400 23860
rect 23799 23820 24400 23848
rect 23799 23817 23811 23820
rect 23753 23811 23811 23817
rect 24394 23808 24400 23820
rect 24452 23808 24458 23860
rect 25958 23848 25964 23860
rect 25919 23820 25964 23848
rect 25958 23808 25964 23820
rect 26016 23808 26022 23860
rect 32122 23808 32128 23860
rect 32180 23848 32186 23860
rect 32217 23851 32275 23857
rect 32217 23848 32229 23851
rect 32180 23820 32229 23848
rect 32180 23808 32186 23820
rect 32217 23817 32229 23820
rect 32263 23817 32275 23851
rect 34514 23848 34520 23860
rect 34475 23820 34520 23848
rect 32217 23811 32275 23817
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 41046 23848 41052 23860
rect 41007 23820 41052 23848
rect 41046 23808 41052 23820
rect 41104 23808 41110 23860
rect 19613 23783 19671 23789
rect 16868 23752 19334 23780
rect 19306 23724 19334 23752
rect 19613 23749 19625 23783
rect 19659 23780 19671 23783
rect 20070 23780 20076 23792
rect 19659 23752 20076 23780
rect 19659 23749 19671 23752
rect 19613 23743 19671 23749
rect 20070 23740 20076 23752
rect 20128 23740 20134 23792
rect 26786 23740 26792 23792
rect 26844 23780 26850 23792
rect 40310 23780 40316 23792
rect 26844 23752 40316 23780
rect 26844 23740 26850 23752
rect 40310 23740 40316 23752
rect 40368 23740 40374 23792
rect 47486 23780 47492 23792
rect 40420 23752 47492 23780
rect 14918 23712 14924 23724
rect 14879 23684 14924 23712
rect 14918 23672 14924 23684
rect 14976 23672 14982 23724
rect 15286 23672 15292 23724
rect 15344 23712 15350 23724
rect 15565 23715 15623 23721
rect 15565 23712 15577 23715
rect 15344 23684 15577 23712
rect 15344 23672 15350 23684
rect 15565 23681 15577 23684
rect 15611 23681 15623 23715
rect 15565 23675 15623 23681
rect 17405 23715 17463 23721
rect 17405 23681 17417 23715
rect 17451 23712 17463 23715
rect 17954 23712 17960 23724
rect 17451 23684 17960 23712
rect 17451 23681 17463 23684
rect 17405 23675 17463 23681
rect 17954 23672 17960 23684
rect 18012 23712 18018 23724
rect 18417 23715 18475 23721
rect 18417 23712 18429 23715
rect 18012 23684 18429 23712
rect 18012 23672 18018 23684
rect 18417 23681 18429 23684
rect 18463 23681 18475 23715
rect 19306 23684 19340 23724
rect 18417 23675 18475 23681
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 23106 23672 23112 23724
rect 23164 23712 23170 23724
rect 23569 23715 23627 23721
rect 23569 23712 23581 23715
rect 23164 23684 23581 23712
rect 23164 23672 23170 23684
rect 23569 23681 23581 23684
rect 23615 23712 23627 23715
rect 24305 23715 24363 23721
rect 24305 23712 24317 23715
rect 23615 23684 24317 23712
rect 23615 23681 23627 23684
rect 23569 23675 23627 23681
rect 24305 23681 24317 23684
rect 24351 23681 24363 23715
rect 24305 23675 24363 23681
rect 24394 23672 24400 23724
rect 24452 23712 24458 23724
rect 25869 23715 25927 23721
rect 25869 23712 25881 23715
rect 24452 23684 25881 23712
rect 24452 23672 24458 23684
rect 25869 23681 25881 23684
rect 25915 23712 25927 23715
rect 26970 23712 26976 23724
rect 25915 23684 26976 23712
rect 25915 23681 25927 23684
rect 25869 23675 25927 23681
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 28626 23672 28632 23724
rect 28684 23712 28690 23724
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 28684 23684 32137 23712
rect 28684 23672 28690 23684
rect 32125 23681 32137 23684
rect 32171 23712 32183 23715
rect 32490 23712 32496 23724
rect 32171 23684 32496 23712
rect 32171 23681 32183 23684
rect 32125 23675 32183 23681
rect 32490 23672 32496 23684
rect 32548 23672 32554 23724
rect 34425 23715 34483 23721
rect 34425 23681 34437 23715
rect 34471 23712 34483 23715
rect 35253 23715 35311 23721
rect 35253 23712 35265 23715
rect 34471 23684 35265 23712
rect 34471 23681 34483 23684
rect 34425 23675 34483 23681
rect 35253 23681 35265 23684
rect 35299 23712 35311 23715
rect 35342 23712 35348 23724
rect 35299 23684 35348 23712
rect 35299 23681 35311 23684
rect 35253 23675 35311 23681
rect 35342 23672 35348 23684
rect 35400 23672 35406 23724
rect 39666 23712 39672 23724
rect 39627 23684 39672 23712
rect 39666 23672 39672 23684
rect 39724 23672 39730 23724
rect 40420 23712 40448 23752
rect 47486 23740 47492 23752
rect 47544 23740 47550 23792
rect 39776 23684 40448 23712
rect 40681 23715 40739 23721
rect 13173 23647 13231 23653
rect 13173 23613 13185 23647
rect 13219 23613 13231 23647
rect 13173 23607 13231 23613
rect 13906 23604 13912 23656
rect 13964 23644 13970 23656
rect 14936 23644 14964 23672
rect 13964 23616 14964 23644
rect 15105 23647 15163 23653
rect 13964 23604 13970 23616
rect 15105 23613 15117 23647
rect 15151 23644 15163 23647
rect 16390 23644 16396 23656
rect 15151 23616 16396 23644
rect 15151 23613 15163 23616
rect 15105 23607 15163 23613
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 18141 23647 18199 23653
rect 18141 23613 18153 23647
rect 18187 23644 18199 23647
rect 19058 23644 19064 23656
rect 18187 23616 19064 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 19058 23604 19064 23616
rect 19116 23604 19122 23656
rect 19429 23647 19487 23653
rect 19429 23613 19441 23647
rect 19475 23628 19487 23647
rect 20806 23644 20812 23656
rect 19475 23613 19564 23628
rect 20767 23616 20812 23644
rect 19429 23607 19564 23613
rect 19444 23600 19564 23607
rect 20806 23604 20812 23616
rect 20864 23604 20870 23656
rect 36265 23647 36323 23653
rect 36265 23613 36277 23647
rect 36311 23613 36323 23647
rect 36265 23607 36323 23613
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 19536 23576 19564 23600
rect 27154 23576 27160 23588
rect 2087 23548 17724 23576
rect 19536 23548 19748 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 14277 23511 14335 23517
rect 14277 23508 14289 23511
rect 13872 23480 14289 23508
rect 13872 23468 13878 23480
rect 14277 23477 14289 23480
rect 14323 23508 14335 23511
rect 14918 23508 14924 23520
rect 14323 23480 14924 23508
rect 14323 23477 14335 23480
rect 14277 23471 14335 23477
rect 14918 23468 14924 23480
rect 14976 23468 14982 23520
rect 15657 23511 15715 23517
rect 15657 23477 15669 23511
rect 15703 23508 15715 23511
rect 17126 23508 17132 23520
rect 15703 23480 17132 23508
rect 15703 23477 15715 23480
rect 15657 23471 15715 23477
rect 17126 23468 17132 23480
rect 17184 23468 17190 23520
rect 17696 23508 17724 23548
rect 19334 23508 19340 23520
rect 17696 23480 19340 23508
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 19720 23508 19748 23548
rect 24412 23548 27160 23576
rect 24412 23508 24440 23548
rect 27154 23536 27160 23548
rect 27212 23536 27218 23588
rect 35986 23536 35992 23588
rect 36044 23576 36050 23588
rect 36280 23576 36308 23607
rect 39390 23604 39396 23656
rect 39448 23644 39454 23656
rect 39577 23647 39635 23653
rect 39577 23644 39589 23647
rect 39448 23616 39589 23644
rect 39448 23604 39454 23616
rect 39577 23613 39589 23616
rect 39623 23613 39635 23647
rect 39577 23607 39635 23613
rect 39776 23576 39804 23684
rect 40681 23681 40693 23715
rect 40727 23712 40739 23715
rect 42610 23712 42616 23724
rect 40727 23684 42616 23712
rect 40727 23681 40739 23684
rect 40681 23675 40739 23681
rect 42610 23672 42616 23684
rect 42668 23672 42674 23724
rect 43254 23712 43260 23724
rect 43215 23684 43260 23712
rect 43254 23672 43260 23684
rect 43312 23672 43318 23724
rect 43441 23715 43499 23721
rect 43441 23681 43453 23715
rect 43487 23712 43499 23715
rect 43898 23712 43904 23724
rect 43487 23684 43904 23712
rect 43487 23681 43499 23684
rect 43441 23675 43499 23681
rect 43898 23672 43904 23684
rect 43956 23672 43962 23724
rect 44082 23712 44088 23724
rect 44043 23684 44088 23712
rect 44082 23672 44088 23684
rect 44140 23672 44146 23724
rect 44269 23715 44327 23721
rect 44269 23681 44281 23715
rect 44315 23681 44327 23715
rect 45738 23712 45744 23724
rect 45699 23684 45744 23712
rect 44269 23675 44327 23681
rect 40589 23647 40647 23653
rect 40589 23644 40601 23647
rect 40052 23616 40601 23644
rect 40052 23585 40080 23616
rect 40589 23613 40601 23616
rect 40635 23613 40647 23647
rect 40589 23607 40647 23613
rect 43625 23647 43683 23653
rect 43625 23613 43637 23647
rect 43671 23644 43683 23647
rect 44284 23644 44312 23675
rect 45738 23672 45744 23684
rect 45796 23672 45802 23724
rect 47026 23672 47032 23724
rect 47084 23712 47090 23724
rect 47581 23715 47639 23721
rect 47581 23712 47593 23715
rect 47084 23684 47593 23712
rect 47084 23672 47090 23684
rect 47581 23681 47593 23684
rect 47627 23681 47639 23715
rect 47581 23675 47639 23681
rect 46198 23644 46204 23656
rect 43671 23616 44312 23644
rect 46159 23616 46204 23644
rect 43671 23613 43683 23616
rect 43625 23607 43683 23613
rect 46198 23604 46204 23616
rect 46256 23604 46262 23656
rect 46477 23647 46535 23653
rect 46477 23613 46489 23647
rect 46523 23613 46535 23647
rect 46477 23607 46535 23613
rect 36044 23548 39804 23576
rect 40037 23579 40095 23585
rect 36044 23536 36050 23548
rect 40037 23545 40049 23579
rect 40083 23545 40095 23579
rect 40037 23539 40095 23545
rect 45646 23536 45652 23588
rect 45704 23576 45710 23588
rect 46492 23576 46520 23607
rect 45704 23548 46520 23576
rect 45704 23536 45710 23548
rect 19720 23480 24440 23508
rect 24489 23511 24547 23517
rect 24489 23477 24501 23511
rect 24535 23508 24547 23511
rect 24578 23508 24584 23520
rect 24535 23480 24584 23508
rect 24535 23477 24547 23480
rect 24489 23471 24547 23477
rect 24578 23468 24584 23480
rect 24636 23468 24642 23520
rect 43806 23468 43812 23520
rect 43864 23508 43870 23520
rect 44085 23511 44143 23517
rect 44085 23508 44097 23511
rect 43864 23480 44097 23508
rect 43864 23468 43870 23480
rect 44085 23477 44097 23480
rect 44131 23477 44143 23511
rect 44085 23471 44143 23477
rect 45557 23511 45615 23517
rect 45557 23477 45569 23511
rect 45603 23508 45615 23511
rect 46934 23508 46940 23520
rect 45603 23480 46940 23508
rect 45603 23477 45615 23480
rect 45557 23471 45615 23477
rect 46934 23468 46940 23480
rect 46992 23468 46998 23520
rect 47670 23508 47676 23520
rect 47631 23480 47676 23508
rect 47670 23468 47676 23480
rect 47728 23468 47734 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 11330 23304 11336 23316
rect 11291 23276 11336 23304
rect 11330 23264 11336 23276
rect 11388 23264 11394 23316
rect 11974 23264 11980 23316
rect 12032 23304 12038 23316
rect 12161 23307 12219 23313
rect 12161 23304 12173 23307
rect 12032 23276 12173 23304
rect 12032 23264 12038 23276
rect 12161 23273 12173 23276
rect 12207 23273 12219 23307
rect 12161 23267 12219 23273
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 13081 23307 13139 23313
rect 13081 23304 13093 23307
rect 12308 23276 13093 23304
rect 12308 23264 12314 23276
rect 13081 23273 13093 23276
rect 13127 23273 13139 23307
rect 13081 23267 13139 23273
rect 13265 23307 13323 23313
rect 13265 23273 13277 23307
rect 13311 23304 13323 23307
rect 14550 23304 14556 23316
rect 13311 23276 14556 23304
rect 13311 23273 13323 23276
rect 13265 23267 13323 23273
rect 14550 23264 14556 23276
rect 14608 23264 14614 23316
rect 14734 23264 14740 23316
rect 14792 23304 14798 23316
rect 16850 23304 16856 23316
rect 14792 23276 16856 23304
rect 14792 23264 14798 23276
rect 16850 23264 16856 23276
rect 16908 23264 16914 23316
rect 19242 23264 19248 23316
rect 19300 23304 19306 23316
rect 20625 23307 20683 23313
rect 20625 23304 20637 23307
rect 19300 23276 20637 23304
rect 19300 23264 19306 23276
rect 20625 23273 20637 23276
rect 20671 23304 20683 23307
rect 21818 23304 21824 23316
rect 20671 23276 21824 23304
rect 20671 23273 20683 23276
rect 20625 23267 20683 23273
rect 21818 23264 21824 23276
rect 21876 23264 21882 23316
rect 22002 23264 22008 23316
rect 22060 23304 22066 23316
rect 22554 23304 22560 23316
rect 22060 23276 22560 23304
rect 22060 23264 22066 23276
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 22646 23264 22652 23316
rect 22704 23304 22710 23316
rect 25685 23307 25743 23313
rect 25685 23304 25697 23307
rect 22704 23276 25697 23304
rect 22704 23264 22710 23276
rect 25685 23273 25697 23276
rect 25731 23304 25743 23307
rect 25866 23304 25872 23316
rect 25731 23276 25872 23304
rect 25731 23273 25743 23276
rect 25685 23267 25743 23273
rect 25866 23264 25872 23276
rect 25924 23264 25930 23316
rect 35710 23264 35716 23316
rect 35768 23304 35774 23316
rect 42334 23304 42340 23316
rect 35768 23276 42340 23304
rect 35768 23264 35774 23276
rect 42334 23264 42340 23276
rect 42392 23264 42398 23316
rect 6886 23208 16528 23236
rect 3602 23128 3608 23180
rect 3660 23168 3666 23180
rect 6886 23168 6914 23208
rect 14090 23168 14096 23180
rect 3660 23140 6914 23168
rect 14051 23140 14096 23168
rect 3660 23128 3666 23140
rect 14090 23128 14096 23140
rect 14148 23128 14154 23180
rect 15746 23168 15752 23180
rect 15707 23140 15752 23168
rect 15746 23128 15752 23140
rect 15804 23128 15810 23180
rect 16390 23168 16396 23180
rect 16351 23140 16396 23168
rect 16390 23128 16396 23140
rect 16448 23128 16454 23180
rect 16500 23168 16528 23208
rect 19334 23196 19340 23248
rect 19392 23236 19398 23248
rect 20530 23236 20536 23248
rect 19392 23208 20536 23236
rect 19392 23196 19398 23208
rect 20530 23196 20536 23208
rect 20588 23236 20594 23248
rect 42521 23239 42579 23245
rect 20588 23208 42288 23236
rect 20588 23196 20594 23208
rect 30653 23171 30711 23177
rect 30653 23168 30665 23171
rect 16500 23140 30665 23168
rect 30653 23137 30665 23140
rect 30699 23137 30711 23171
rect 35710 23168 35716 23180
rect 35671 23140 35716 23168
rect 30653 23131 30711 23137
rect 35710 23128 35716 23140
rect 35768 23128 35774 23180
rect 40494 23168 40500 23180
rect 40455 23140 40500 23168
rect 40494 23128 40500 23140
rect 40552 23128 40558 23180
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23100 9919 23103
rect 9950 23100 9956 23112
rect 9907 23072 9956 23100
rect 9907 23069 9919 23072
rect 9861 23063 9919 23069
rect 9950 23060 9956 23072
rect 10008 23060 10014 23112
rect 10689 23103 10747 23109
rect 10689 23069 10701 23103
rect 10735 23100 10747 23103
rect 11054 23100 11060 23112
rect 10735 23072 11060 23100
rect 10735 23069 10747 23072
rect 10689 23063 10747 23069
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 11606 23100 11612 23112
rect 11567 23072 11612 23100
rect 11606 23060 11612 23072
rect 11664 23060 11670 23112
rect 12069 23103 12127 23109
rect 12069 23069 12081 23103
rect 12115 23100 12127 23103
rect 12115 23072 14136 23100
rect 12115 23069 12127 23072
rect 12069 23063 12127 23069
rect 11333 23035 11391 23041
rect 11333 23001 11345 23035
rect 11379 23032 11391 23035
rect 11790 23032 11796 23044
rect 11379 23004 11796 23032
rect 11379 23001 11391 23004
rect 11333 22995 11391 23001
rect 11790 22992 11796 23004
rect 11848 23032 11854 23044
rect 12897 23035 12955 23041
rect 12897 23032 12909 23035
rect 11848 23004 12909 23032
rect 11848 22992 11854 23004
rect 12897 23001 12909 23004
rect 12943 23001 12955 23035
rect 12897 22995 12955 23001
rect 9858 22964 9864 22976
rect 9819 22936 9864 22964
rect 9858 22924 9864 22936
rect 9916 22924 9922 22976
rect 10778 22964 10784 22976
rect 10739 22936 10784 22964
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 11517 22967 11575 22973
rect 11517 22933 11529 22967
rect 11563 22964 11575 22967
rect 12250 22964 12256 22976
rect 11563 22936 12256 22964
rect 11563 22933 11575 22936
rect 11517 22927 11575 22933
rect 12250 22924 12256 22936
rect 12308 22924 12314 22976
rect 13078 22924 13084 22976
rect 13136 22973 13142 22976
rect 13136 22967 13155 22973
rect 13143 22933 13155 22967
rect 14108 22964 14136 23072
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19392 23072 19437 23100
rect 19392 23060 19398 23072
rect 20070 23060 20076 23112
rect 20128 23100 20134 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20128 23072 20453 23100
rect 20128 23060 20134 23072
rect 20441 23069 20453 23072
rect 20487 23100 20499 23103
rect 21358 23100 21364 23112
rect 20487 23072 21364 23100
rect 20487 23069 20499 23072
rect 20441 23063 20499 23069
rect 21358 23060 21364 23072
rect 21416 23060 21422 23112
rect 22830 23100 22836 23112
rect 22791 23072 22836 23100
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 23474 23100 23480 23112
rect 23435 23072 23480 23100
rect 23474 23060 23480 23072
rect 23532 23060 23538 23112
rect 25498 23100 25504 23112
rect 25411 23072 25504 23100
rect 25498 23060 25504 23072
rect 25556 23060 25562 23112
rect 28258 23100 28264 23112
rect 28219 23072 28264 23100
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 30190 23100 30196 23112
rect 30151 23072 30196 23100
rect 30190 23060 30196 23072
rect 30248 23060 30254 23112
rect 33134 23060 33140 23112
rect 33192 23100 33198 23112
rect 33689 23103 33747 23109
rect 33689 23100 33701 23103
rect 33192 23072 33701 23100
rect 33192 23060 33198 23072
rect 33689 23069 33701 23072
rect 33735 23100 33747 23103
rect 35161 23103 35219 23109
rect 33735 23072 35112 23100
rect 33735 23069 33747 23072
rect 33689 23063 33747 23069
rect 14274 23032 14280 23044
rect 14235 23004 14280 23032
rect 14274 22992 14280 23004
rect 14332 22992 14338 23044
rect 14458 22992 14464 23044
rect 14516 23032 14522 23044
rect 15286 23032 15292 23044
rect 14516 23004 15292 23032
rect 14516 22992 14522 23004
rect 15286 22992 15292 23004
rect 15344 22992 15350 23044
rect 15470 22992 15476 23044
rect 15528 23032 15534 23044
rect 16669 23035 16727 23041
rect 16669 23032 16681 23035
rect 15528 23004 16681 23032
rect 15528 22992 15534 23004
rect 16669 23001 16681 23004
rect 16715 23001 16727 23035
rect 16669 22995 16727 23001
rect 17126 22992 17132 23044
rect 17184 22992 17190 23044
rect 18414 22992 18420 23044
rect 18472 23032 18478 23044
rect 19889 23035 19947 23041
rect 19889 23032 19901 23035
rect 18472 23004 19901 23032
rect 18472 22992 18478 23004
rect 19889 23001 19901 23004
rect 19935 23032 19947 23035
rect 20714 23032 20720 23044
rect 19935 23004 20720 23032
rect 19935 23001 19947 23004
rect 19889 22995 19947 23001
rect 20714 22992 20720 23004
rect 20772 22992 20778 23044
rect 22554 22992 22560 23044
rect 22612 23032 22618 23044
rect 25516 23032 25544 23060
rect 22612 23004 25544 23032
rect 30377 23035 30435 23041
rect 22612 22992 22618 23004
rect 30377 23001 30389 23035
rect 30423 23032 30435 23035
rect 32214 23032 32220 23044
rect 30423 23004 32220 23032
rect 30423 23001 30435 23004
rect 30377 22995 30435 23001
rect 32214 22992 32220 23004
rect 32272 22992 32278 23044
rect 16574 22964 16580 22976
rect 14108 22936 16580 22964
rect 13136 22927 13155 22933
rect 13136 22924 13142 22927
rect 16574 22924 16580 22936
rect 16632 22924 16638 22976
rect 16850 22924 16856 22976
rect 16908 22964 16914 22976
rect 18141 22967 18199 22973
rect 18141 22964 18153 22967
rect 16908 22936 18153 22964
rect 16908 22924 16914 22936
rect 18141 22933 18153 22936
rect 18187 22933 18199 22967
rect 22922 22964 22928 22976
rect 22883 22936 22928 22964
rect 18141 22927 18199 22933
rect 22922 22924 22928 22936
rect 22980 22924 22986 22976
rect 23382 22924 23388 22976
rect 23440 22964 23446 22976
rect 23569 22967 23627 22973
rect 23569 22964 23581 22967
rect 23440 22936 23581 22964
rect 23440 22924 23446 22936
rect 23569 22933 23581 22936
rect 23615 22933 23627 22967
rect 23569 22927 23627 22933
rect 28353 22967 28411 22973
rect 28353 22933 28365 22967
rect 28399 22964 28411 22967
rect 28718 22964 28724 22976
rect 28399 22936 28724 22964
rect 28399 22933 28411 22936
rect 28353 22927 28411 22933
rect 28718 22924 28724 22936
rect 28776 22924 28782 22976
rect 33778 22964 33784 22976
rect 33739 22936 33784 22964
rect 33778 22924 33784 22936
rect 33836 22924 33842 22976
rect 35084 22964 35112 23072
rect 35161 23069 35173 23103
rect 35207 23100 35219 23103
rect 35342 23100 35348 23112
rect 35207 23072 35348 23100
rect 35207 23069 35219 23072
rect 35161 23063 35219 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 39850 23100 39856 23112
rect 39811 23072 39856 23100
rect 39850 23060 39856 23072
rect 39908 23060 39914 23112
rect 42260 23109 42288 23208
rect 42521 23205 42533 23239
rect 42567 23236 42579 23239
rect 45922 23236 45928 23248
rect 42567 23208 45928 23236
rect 42567 23205 42579 23208
rect 42521 23199 42579 23205
rect 42245 23103 42303 23109
rect 42245 23069 42257 23103
rect 42291 23100 42303 23103
rect 42426 23100 42432 23112
rect 42291 23072 42432 23100
rect 42291 23069 42303 23072
rect 42245 23063 42303 23069
rect 42426 23060 42432 23072
rect 42484 23060 42490 23112
rect 39482 22992 39488 23044
rect 39540 23032 39546 23044
rect 40037 23035 40095 23041
rect 40037 23032 40049 23035
rect 39540 23004 40049 23032
rect 39540 22992 39546 23004
rect 40037 23001 40049 23004
rect 40083 23001 40095 23035
rect 40037 22995 40095 23001
rect 39574 22964 39580 22976
rect 35084 22936 39580 22964
rect 39574 22924 39580 22936
rect 39632 22964 39638 22976
rect 42536 22964 42564 23199
rect 45922 23196 45928 23208
rect 45980 23196 45986 23248
rect 46382 23196 46388 23248
rect 46440 23196 46446 23248
rect 43622 23168 43628 23180
rect 43583 23140 43628 23168
rect 43622 23128 43628 23140
rect 43680 23128 43686 23180
rect 46293 23171 46351 23177
rect 46293 23137 46305 23171
rect 46339 23168 46351 23171
rect 46400 23168 46428 23196
rect 46339 23140 46428 23168
rect 46477 23171 46535 23177
rect 46339 23137 46351 23140
rect 46293 23131 46351 23137
rect 46477 23137 46489 23171
rect 46523 23168 46535 23171
rect 47670 23168 47676 23180
rect 46523 23140 47676 23168
rect 46523 23137 46535 23140
rect 46477 23131 46535 23137
rect 47670 23128 47676 23140
rect 47728 23128 47734 23180
rect 48133 23171 48191 23177
rect 48133 23137 48145 23171
rect 48179 23168 48191 23171
rect 48222 23168 48228 23180
rect 48179 23140 48228 23168
rect 48179 23137 48191 23140
rect 48133 23131 48191 23137
rect 48222 23128 48228 23140
rect 48280 23128 48286 23180
rect 43806 23100 43812 23112
rect 43767 23072 43812 23100
rect 43806 23060 43812 23072
rect 43864 23060 43870 23112
rect 45833 23103 45891 23109
rect 45833 23069 45845 23103
rect 45879 23100 45891 23103
rect 45879 23072 46336 23100
rect 45879 23069 45891 23072
rect 45833 23063 45891 23069
rect 44453 23035 44511 23041
rect 44453 23001 44465 23035
rect 44499 23032 44511 23035
rect 45554 23032 45560 23044
rect 44499 23004 45560 23032
rect 44499 23001 44511 23004
rect 44453 22995 44511 23001
rect 45554 22992 45560 23004
rect 45612 23032 45618 23044
rect 46308 23032 46336 23072
rect 47762 23032 47768 23044
rect 45612 23004 45784 23032
rect 46308 23004 47768 23032
rect 45612 22992 45618 23004
rect 39632 22936 42564 22964
rect 39632 22924 39638 22936
rect 45370 22924 45376 22976
rect 45428 22964 45434 22976
rect 45649 22967 45707 22973
rect 45649 22964 45661 22967
rect 45428 22936 45661 22964
rect 45428 22924 45434 22936
rect 45649 22933 45661 22936
rect 45695 22933 45707 22967
rect 45756 22964 45784 23004
rect 47762 22992 47768 23004
rect 47820 22992 47826 23044
rect 46290 22964 46296 22976
rect 45756 22936 46296 22964
rect 45649 22927 45707 22933
rect 46290 22924 46296 22936
rect 46348 22924 46354 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 9950 22720 9956 22772
rect 10008 22760 10014 22772
rect 10873 22763 10931 22769
rect 10873 22760 10885 22763
rect 10008 22732 10885 22760
rect 10008 22720 10014 22732
rect 10873 22729 10885 22732
rect 10919 22729 10931 22763
rect 11882 22760 11888 22772
rect 11795 22732 11888 22760
rect 10873 22723 10931 22729
rect 11882 22720 11888 22732
rect 11940 22760 11946 22772
rect 12250 22760 12256 22772
rect 11940 22732 12256 22760
rect 11940 22720 11946 22732
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 13541 22763 13599 22769
rect 13541 22729 13553 22763
rect 13587 22760 13599 22763
rect 14303 22763 14361 22769
rect 13587 22732 14228 22760
rect 13587 22729 13599 22732
rect 13541 22723 13599 22729
rect 11238 22692 11244 22704
rect 8220 22664 11244 22692
rect 8220 22633 8248 22664
rect 11238 22652 11244 22664
rect 11296 22692 11302 22704
rect 11517 22695 11575 22701
rect 11517 22692 11529 22695
rect 11296 22664 11529 22692
rect 11296 22652 11302 22664
rect 11517 22661 11529 22664
rect 11563 22661 11575 22695
rect 11517 22655 11575 22661
rect 11733 22695 11791 22701
rect 11733 22661 11745 22695
rect 11779 22692 11791 22695
rect 12158 22692 12164 22704
rect 11779 22664 12164 22692
rect 11779 22661 11791 22664
rect 11733 22655 11791 22661
rect 12158 22652 12164 22664
rect 12216 22652 12222 22704
rect 14093 22695 14151 22701
rect 14093 22661 14105 22695
rect 14139 22661 14151 22695
rect 14200 22692 14228 22732
rect 14303 22729 14315 22763
rect 14349 22760 14361 22763
rect 14734 22760 14740 22772
rect 14349 22732 14740 22760
rect 14349 22729 14361 22732
rect 14303 22723 14361 22729
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 22002 22760 22008 22772
rect 14844 22732 22008 22760
rect 14458 22692 14464 22704
rect 14200 22664 14464 22692
rect 14093 22655 14151 22661
rect 8205 22627 8263 22633
rect 8205 22593 8217 22627
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 11330 22624 11336 22636
rect 10735 22596 11336 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 11330 22584 11336 22596
rect 11388 22584 11394 22636
rect 12529 22627 12587 22633
rect 12529 22593 12541 22627
rect 12575 22624 12587 22627
rect 13357 22627 13415 22633
rect 13357 22624 13369 22627
rect 12575 22596 13369 22624
rect 12575 22593 12587 22596
rect 12529 22587 12587 22593
rect 13357 22593 13369 22596
rect 13403 22624 13415 22627
rect 13814 22624 13820 22636
rect 13403 22596 13820 22624
rect 13403 22593 13415 22596
rect 13357 22587 13415 22593
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 14108 22624 14136 22655
rect 14458 22652 14464 22664
rect 14516 22652 14522 22704
rect 14844 22624 14872 22732
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 32214 22760 32220 22772
rect 25148 22732 31754 22760
rect 32175 22732 32220 22760
rect 21913 22695 21971 22701
rect 21913 22692 21925 22695
rect 20746 22664 21925 22692
rect 21913 22661 21925 22664
rect 21959 22661 21971 22695
rect 21913 22655 21971 22661
rect 22922 22652 22928 22704
rect 22980 22692 22986 22704
rect 25148 22701 25176 22732
rect 23477 22695 23535 22701
rect 23477 22692 23489 22695
rect 22980 22664 23489 22692
rect 22980 22652 22986 22664
rect 23477 22661 23489 22664
rect 23523 22661 23535 22695
rect 23477 22655 23535 22661
rect 25133 22695 25191 22701
rect 25133 22661 25145 22695
rect 25179 22661 25191 22695
rect 28258 22692 28264 22704
rect 25133 22655 25191 22661
rect 25976 22664 28264 22692
rect 14108 22596 14872 22624
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22624 15163 22627
rect 15838 22624 15844 22636
rect 15151 22596 15844 22624
rect 15151 22593 15163 22596
rect 15105 22587 15163 22593
rect 15838 22584 15844 22596
rect 15896 22624 15902 22636
rect 16850 22624 16856 22636
rect 15896 22596 16856 22624
rect 15896 22584 15902 22596
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 21818 22624 21824 22636
rect 21779 22596 21824 22624
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 25976 22633 26004 22664
rect 28258 22652 28264 22664
rect 28316 22652 28322 22704
rect 29638 22652 29644 22704
rect 29696 22652 29702 22704
rect 31726 22692 31754 22732
rect 32214 22720 32220 22732
rect 32272 22720 32278 22772
rect 37274 22760 37280 22772
rect 32324 22732 37280 22760
rect 32324 22692 32352 22732
rect 37274 22720 37280 22732
rect 37332 22720 37338 22772
rect 39482 22760 39488 22772
rect 39443 22732 39488 22760
rect 39482 22720 39488 22732
rect 39540 22720 39546 22772
rect 41892 22732 46888 22760
rect 33778 22692 33784 22704
rect 31726 22664 32352 22692
rect 33739 22664 33784 22692
rect 33778 22652 33784 22664
rect 33836 22652 33842 22704
rect 41892 22701 41920 22732
rect 41877 22695 41935 22701
rect 41877 22661 41889 22695
rect 41923 22661 41935 22695
rect 41877 22655 41935 22661
rect 43349 22695 43407 22701
rect 43349 22661 43361 22695
rect 43395 22692 43407 22695
rect 43990 22692 43996 22704
rect 43395 22664 43996 22692
rect 43395 22661 43407 22664
rect 43349 22655 43407 22661
rect 43990 22652 43996 22664
rect 44048 22652 44054 22704
rect 45370 22692 45376 22704
rect 45331 22664 45376 22692
rect 45370 22652 45376 22664
rect 45428 22652 45434 22704
rect 25961 22627 26019 22633
rect 25961 22624 25973 22627
rect 25884 22596 25973 22624
rect 8386 22556 8392 22568
rect 8347 22528 8392 22556
rect 8386 22516 8392 22528
rect 8444 22516 8450 22568
rect 8665 22559 8723 22565
rect 8665 22525 8677 22559
rect 8711 22525 8723 22559
rect 15194 22556 15200 22568
rect 15155 22528 15200 22556
rect 8665 22519 8723 22525
rect 3694 22448 3700 22500
rect 3752 22488 3758 22500
rect 8680 22488 8708 22519
rect 15194 22516 15200 22528
rect 15252 22516 15258 22568
rect 15470 22556 15476 22568
rect 15431 22528 15476 22556
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 17034 22556 17040 22568
rect 16995 22528 17040 22556
rect 17034 22516 17040 22528
rect 17092 22516 17098 22568
rect 18690 22556 18696 22568
rect 18651 22528 18696 22556
rect 18690 22516 18696 22528
rect 18748 22516 18754 22568
rect 19245 22559 19303 22565
rect 19245 22525 19257 22559
rect 19291 22556 19303 22559
rect 19521 22559 19579 22565
rect 19291 22528 19380 22556
rect 19291 22525 19303 22528
rect 19245 22519 19303 22525
rect 3752 22460 8708 22488
rect 3752 22448 3758 22460
rect 11054 22448 11060 22500
rect 11112 22488 11118 22500
rect 11112 22460 12020 22488
rect 11112 22448 11118 22460
rect 11992 22432 12020 22460
rect 13078 22448 13084 22500
rect 13136 22488 13142 22500
rect 15654 22488 15660 22500
rect 13136 22460 15660 22488
rect 13136 22448 13142 22460
rect 11698 22420 11704 22432
rect 11659 22392 11704 22420
rect 11698 22380 11704 22392
rect 11756 22380 11762 22432
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 12342 22420 12348 22432
rect 12032 22392 12348 22420
rect 12032 22380 12038 22392
rect 12342 22380 12348 22392
rect 12400 22420 12406 22432
rect 14292 22429 14320 22460
rect 15654 22448 15660 22460
rect 15712 22448 15718 22500
rect 19352 22432 19380 22528
rect 19521 22525 19533 22559
rect 19567 22556 19579 22559
rect 19978 22556 19984 22568
rect 19567 22528 19984 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 19978 22516 19984 22528
rect 20036 22516 20042 22568
rect 21266 22556 21272 22568
rect 21227 22528 21272 22556
rect 21266 22516 21272 22528
rect 21324 22516 21330 22568
rect 23290 22556 23296 22568
rect 23251 22528 23296 22556
rect 23290 22516 23296 22528
rect 23348 22516 23354 22568
rect 23106 22448 23112 22500
rect 23164 22488 23170 22500
rect 25884 22488 25912 22596
rect 25961 22593 25973 22596
rect 26007 22593 26019 22627
rect 25961 22587 26019 22593
rect 27065 22627 27123 22633
rect 27065 22593 27077 22627
rect 27111 22624 27123 22627
rect 27338 22624 27344 22636
rect 27111 22596 27344 22624
rect 27111 22593 27123 22596
rect 27065 22587 27123 22593
rect 27338 22584 27344 22596
rect 27396 22584 27402 22636
rect 27893 22627 27951 22633
rect 27893 22593 27905 22627
rect 27939 22624 27951 22627
rect 28718 22624 28724 22636
rect 27939 22596 28212 22624
rect 28679 22596 28724 22624
rect 27939 22593 27951 22596
rect 27893 22587 27951 22593
rect 27982 22556 27988 22568
rect 27943 22528 27988 22556
rect 27982 22516 27988 22528
rect 28040 22516 28046 22568
rect 23164 22460 25912 22488
rect 23164 22448 23170 22460
rect 12713 22423 12771 22429
rect 12713 22420 12725 22423
rect 12400 22392 12725 22420
rect 12400 22380 12406 22392
rect 12713 22389 12725 22392
rect 12759 22389 12771 22423
rect 12713 22383 12771 22389
rect 14277 22423 14335 22429
rect 14277 22389 14289 22423
rect 14323 22389 14335 22423
rect 14458 22420 14464 22432
rect 14419 22392 14464 22420
rect 14277 22383 14335 22389
rect 14458 22380 14464 22392
rect 14516 22380 14522 22432
rect 19334 22380 19340 22432
rect 19392 22380 19398 22432
rect 25958 22420 25964 22432
rect 25919 22392 25964 22420
rect 25958 22380 25964 22392
rect 26016 22380 26022 22432
rect 27062 22380 27068 22432
rect 27120 22420 27126 22432
rect 27157 22423 27215 22429
rect 27157 22420 27169 22423
rect 27120 22392 27169 22420
rect 27120 22380 27126 22392
rect 27157 22389 27169 22392
rect 27203 22389 27215 22423
rect 28184 22420 28212 22596
rect 28718 22584 28724 22596
rect 28776 22584 28782 22636
rect 32125 22627 32183 22633
rect 32125 22593 32137 22627
rect 32171 22624 32183 22627
rect 33134 22624 33140 22636
rect 32171 22596 33140 22624
rect 32171 22593 32183 22596
rect 32125 22587 32183 22593
rect 33134 22584 33140 22596
rect 33192 22584 33198 22636
rect 39393 22627 39451 22633
rect 39393 22593 39405 22627
rect 39439 22624 39451 22627
rect 39574 22624 39580 22636
rect 39439 22596 39580 22624
rect 39439 22593 39451 22596
rect 39393 22587 39451 22593
rect 39574 22584 39580 22596
rect 39632 22584 39638 22636
rect 40034 22624 40040 22636
rect 39995 22596 40040 22624
rect 40034 22584 40040 22596
rect 40092 22584 40098 22636
rect 42426 22624 42432 22636
rect 42387 22596 42432 22624
rect 42426 22584 42432 22596
rect 42484 22584 42490 22636
rect 43530 22624 43536 22636
rect 43491 22596 43536 22624
rect 43530 22584 43536 22596
rect 43588 22584 43594 22636
rect 43622 22584 43628 22636
rect 43680 22624 43686 22636
rect 43680 22596 43725 22624
rect 43680 22584 43686 22596
rect 43898 22584 43904 22636
rect 43956 22624 43962 22636
rect 44085 22627 44143 22633
rect 44085 22624 44097 22627
rect 43956 22596 44097 22624
rect 43956 22584 43962 22596
rect 44085 22593 44097 22596
rect 44131 22593 44143 22627
rect 44266 22624 44272 22636
rect 44227 22596 44272 22624
rect 44085 22587 44143 22593
rect 44266 22584 44272 22596
rect 44324 22584 44330 22636
rect 28261 22559 28319 22565
rect 28261 22525 28273 22559
rect 28307 22556 28319 22559
rect 28997 22559 29055 22565
rect 28997 22556 29009 22559
rect 28307 22528 29009 22556
rect 28307 22525 28319 22528
rect 28261 22519 28319 22525
rect 28997 22525 29009 22528
rect 29043 22525 29055 22559
rect 28997 22519 29055 22525
rect 29086 22516 29092 22568
rect 29144 22556 29150 22568
rect 33597 22559 33655 22565
rect 33597 22556 33609 22559
rect 29144 22528 33609 22556
rect 29144 22516 29150 22528
rect 33597 22525 33609 22528
rect 33643 22525 33655 22559
rect 33597 22519 33655 22525
rect 35437 22559 35495 22565
rect 35437 22525 35449 22559
rect 35483 22525 35495 22559
rect 40218 22556 40224 22568
rect 40179 22528 40224 22556
rect 35437 22519 35495 22525
rect 35452 22488 35480 22519
rect 40218 22516 40224 22528
rect 40276 22516 40282 22568
rect 42705 22559 42763 22565
rect 42705 22525 42717 22559
rect 42751 22556 42763 22559
rect 45189 22559 45247 22565
rect 42751 22528 44404 22556
rect 42751 22525 42763 22528
rect 42705 22519 42763 22525
rect 42518 22488 42524 22500
rect 35452 22460 42524 22488
rect 42518 22448 42524 22460
rect 42576 22448 42582 22500
rect 42610 22448 42616 22500
rect 42668 22488 42674 22500
rect 43349 22491 43407 22497
rect 43349 22488 43361 22491
rect 42668 22460 43361 22488
rect 42668 22448 42674 22460
rect 43349 22457 43361 22460
rect 43395 22457 43407 22491
rect 44082 22488 44088 22500
rect 44043 22460 44088 22488
rect 43349 22451 43407 22457
rect 44082 22448 44088 22460
rect 44140 22448 44146 22500
rect 44376 22488 44404 22528
rect 45189 22525 45201 22559
rect 45235 22556 45247 22559
rect 45554 22556 45560 22568
rect 45235 22528 45560 22556
rect 45235 22525 45247 22528
rect 45189 22519 45247 22525
rect 45554 22516 45560 22528
rect 45612 22516 45618 22568
rect 46860 22565 46888 22732
rect 47670 22720 47676 22772
rect 47728 22760 47734 22772
rect 47949 22763 48007 22769
rect 47949 22760 47961 22763
rect 47728 22732 47961 22760
rect 47728 22720 47734 22732
rect 47949 22729 47961 22732
rect 47995 22729 48007 22763
rect 47949 22723 48007 22729
rect 46934 22652 46940 22704
rect 46992 22692 46998 22704
rect 47765 22695 47823 22701
rect 47765 22692 47777 22695
rect 46992 22664 47777 22692
rect 46992 22652 46998 22664
rect 47765 22661 47777 22664
rect 47811 22661 47823 22695
rect 47765 22655 47823 22661
rect 47118 22584 47124 22636
rect 47176 22624 47182 22636
rect 47578 22624 47584 22636
rect 47176 22596 47584 22624
rect 47176 22584 47182 22596
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 47854 22624 47860 22636
rect 47815 22596 47860 22624
rect 47854 22584 47860 22596
rect 47912 22584 47918 22636
rect 46845 22559 46903 22565
rect 46845 22525 46857 22559
rect 46891 22556 46903 22559
rect 47210 22556 47216 22568
rect 46891 22528 47216 22556
rect 46891 22525 46903 22528
rect 46845 22519 46903 22525
rect 47210 22516 47216 22528
rect 47268 22516 47274 22568
rect 47486 22488 47492 22500
rect 44376 22460 47492 22488
rect 47486 22448 47492 22460
rect 47544 22448 47550 22500
rect 30190 22420 30196 22432
rect 28184 22392 30196 22420
rect 27157 22383 27215 22389
rect 30190 22380 30196 22392
rect 30248 22420 30254 22432
rect 30469 22423 30527 22429
rect 30469 22420 30481 22423
rect 30248 22392 30481 22420
rect 30248 22380 30254 22392
rect 30469 22389 30481 22392
rect 30515 22389 30527 22423
rect 30469 22383 30527 22389
rect 43254 22380 43260 22432
rect 43312 22420 43318 22432
rect 44266 22420 44272 22432
rect 43312 22392 44272 22420
rect 43312 22380 43318 22392
rect 44266 22380 44272 22392
rect 44324 22380 44330 22432
rect 48130 22420 48136 22432
rect 48091 22392 48136 22420
rect 48130 22380 48136 22392
rect 48188 22380 48194 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8386 22216 8392 22228
rect 8343 22188 8392 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8386 22176 8392 22188
rect 8444 22176 8450 22228
rect 9756 22219 9814 22225
rect 9756 22185 9768 22219
rect 9802 22216 9814 22219
rect 11701 22219 11759 22225
rect 11701 22216 11713 22219
rect 9802 22188 11713 22216
rect 9802 22185 9814 22188
rect 9756 22179 9814 22185
rect 11701 22185 11713 22188
rect 11747 22185 11759 22219
rect 11701 22179 11759 22185
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 15105 22219 15163 22225
rect 15105 22216 15117 22219
rect 14332 22188 15117 22216
rect 14332 22176 14338 22188
rect 15105 22185 15117 22188
rect 15151 22185 15163 22219
rect 15105 22179 15163 22185
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 16945 22219 17003 22225
rect 16945 22216 16957 22219
rect 16632 22188 16957 22216
rect 16632 22176 16638 22188
rect 16945 22185 16957 22188
rect 16991 22185 17003 22219
rect 16945 22179 17003 22185
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 20622 22216 20628 22228
rect 18288 22188 20628 22216
rect 18288 22176 18294 22188
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 21266 22176 21272 22228
rect 21324 22216 21330 22228
rect 39850 22216 39856 22228
rect 21324 22188 39856 22216
rect 21324 22176 21330 22188
rect 39850 22176 39856 22188
rect 39908 22176 39914 22228
rect 40126 22216 40132 22228
rect 40087 22188 40132 22216
rect 40126 22176 40132 22188
rect 40184 22176 40190 22228
rect 40218 22176 40224 22228
rect 40276 22216 40282 22228
rect 40957 22219 41015 22225
rect 40957 22216 40969 22219
rect 40276 22188 40969 22216
rect 40276 22176 40282 22188
rect 40957 22185 40969 22188
rect 41003 22185 41015 22219
rect 40957 22179 41015 22185
rect 43257 22219 43315 22225
rect 43257 22185 43269 22219
rect 43303 22216 43315 22219
rect 43530 22216 43536 22228
rect 43303 22188 43536 22216
rect 43303 22185 43315 22188
rect 43257 22179 43315 22185
rect 43530 22176 43536 22188
rect 43588 22176 43594 22228
rect 44450 22176 44456 22228
rect 44508 22216 44514 22228
rect 48038 22216 48044 22228
rect 44508 22188 48044 22216
rect 44508 22176 44514 22188
rect 48038 22176 48044 22188
rect 48096 22176 48102 22228
rect 11238 22148 11244 22160
rect 11199 22120 11244 22148
rect 11238 22108 11244 22120
rect 11296 22148 11302 22160
rect 12253 22151 12311 22157
rect 12253 22148 12265 22151
rect 11296 22120 12265 22148
rect 11296 22108 11302 22120
rect 12253 22117 12265 22120
rect 12299 22117 12311 22151
rect 12253 22111 12311 22117
rect 14918 22108 14924 22160
rect 14976 22148 14982 22160
rect 20070 22148 20076 22160
rect 14976 22120 20076 22148
rect 14976 22108 14982 22120
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 20441 22151 20499 22157
rect 20441 22148 20453 22151
rect 20364 22120 20453 22148
rect 9493 22083 9551 22089
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9858 22080 9864 22092
rect 9539 22052 9864 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 9858 22040 9864 22052
rect 9916 22040 9922 22092
rect 11330 22040 11336 22092
rect 11388 22080 11394 22092
rect 17586 22080 17592 22092
rect 11388 22052 14136 22080
rect 11388 22040 11394 22052
rect 14108 22024 14136 22052
rect 15028 22052 17592 22080
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 22012 8263 22015
rect 8938 22012 8944 22024
rect 8251 21984 8944 22012
rect 8251 21981 8263 21984
rect 8205 21975 8263 21981
rect 8938 21972 8944 21984
rect 8996 21972 9002 22024
rect 11882 22012 11888 22024
rect 11843 21984 11888 22012
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 22012 12403 22015
rect 12802 22012 12808 22024
rect 12391 21984 12808 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 14090 22012 14096 22024
rect 14051 21984 14096 22012
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 15028 22021 15056 22052
rect 17586 22040 17592 22052
rect 17644 22040 17650 22092
rect 19886 22080 19892 22092
rect 19847 22052 19892 22080
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 21981 15071 22015
rect 15013 21975 15071 21981
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 22012 16083 22015
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16071 21984 16865 22012
rect 16071 21981 16083 21984
rect 16025 21975 16083 21981
rect 16853 21981 16865 21984
rect 16899 22012 16911 22015
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 16899 21984 17785 22012
rect 16899 21981 16911 21984
rect 16853 21975 16911 21981
rect 17773 21981 17785 21984
rect 17819 22012 17831 22015
rect 17954 22012 17960 22024
rect 17819 21984 17960 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 19337 22015 19395 22021
rect 19337 21981 19349 22015
rect 19383 22012 19395 22015
rect 19426 22012 19432 22024
rect 19383 21984 19432 22012
rect 19383 21981 19395 21984
rect 19337 21975 19395 21981
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 19628 21984 20024 22012
rect 10778 21904 10784 21956
rect 10836 21904 10842 21956
rect 12894 21944 12900 21956
rect 12807 21916 12900 21944
rect 12894 21904 12900 21916
rect 12952 21944 12958 21956
rect 14458 21944 14464 21956
rect 12952 21916 14464 21944
rect 12952 21904 12958 21916
rect 14458 21904 14464 21916
rect 14516 21904 14522 21956
rect 18325 21947 18383 21953
rect 18325 21913 18337 21947
rect 18371 21944 18383 21947
rect 19058 21944 19064 21956
rect 18371 21916 19064 21944
rect 18371 21913 18383 21916
rect 18325 21907 18383 21913
rect 19058 21904 19064 21916
rect 19116 21944 19122 21956
rect 19628 21944 19656 21984
rect 19116 21916 19656 21944
rect 19996 21944 20024 21984
rect 20070 21972 20076 22024
rect 20128 22012 20134 22024
rect 20364 22012 20392 22120
rect 20441 22117 20453 22120
rect 20487 22117 20499 22151
rect 21284 22148 21312 22176
rect 20441 22111 20499 22117
rect 20548 22120 21312 22148
rect 20128 21984 20392 22012
rect 20441 22015 20499 22021
rect 20128 21972 20134 21984
rect 20441 21981 20453 22015
rect 20487 22012 20499 22015
rect 20548 22012 20576 22120
rect 21358 22108 21364 22160
rect 21416 22148 21422 22160
rect 21416 22120 22140 22148
rect 21416 22108 21422 22120
rect 21082 22080 21088 22092
rect 20732 22052 21088 22080
rect 20487 21984 20576 22012
rect 20487 21981 20499 21984
rect 20441 21975 20499 21981
rect 20622 21972 20628 22024
rect 20680 22012 20686 22024
rect 20732 22021 20760 22052
rect 21082 22040 21088 22052
rect 21140 22040 21146 22092
rect 21249 22083 21307 22089
rect 21249 22049 21261 22083
rect 21295 22080 21307 22083
rect 22112 22080 22140 22120
rect 27982 22108 27988 22160
rect 28040 22148 28046 22160
rect 28905 22151 28963 22157
rect 28905 22148 28917 22151
rect 28040 22120 28917 22148
rect 28040 22108 28046 22120
rect 28905 22117 28917 22120
rect 28951 22117 28963 22151
rect 28905 22111 28963 22117
rect 43162 22108 43168 22160
rect 43220 22148 43226 22160
rect 43898 22148 43904 22160
rect 43220 22120 43904 22148
rect 43220 22108 43226 22120
rect 43898 22108 43904 22120
rect 43956 22108 43962 22160
rect 45388 22120 45554 22148
rect 21295 22052 22048 22080
rect 22112 22052 22876 22080
rect 21295 22049 21307 22052
rect 21249 22043 21307 22049
rect 20717 22015 20775 22021
rect 20717 22012 20729 22015
rect 20680 21984 20729 22012
rect 20680 21972 20686 21984
rect 20717 21981 20729 21984
rect 20763 21981 20775 22015
rect 20717 21975 20775 21981
rect 20990 21972 20996 22024
rect 21048 22012 21054 22024
rect 22020 22021 22048 22052
rect 21453 22015 21511 22021
rect 21453 22012 21465 22015
rect 21048 21984 21465 22012
rect 21048 21972 21054 21984
rect 21453 21981 21465 21984
rect 21499 21981 21511 22015
rect 21453 21975 21511 21981
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22848 22021 22876 22052
rect 25958 22040 25964 22092
rect 26016 22080 26022 22092
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 26016 22052 26065 22080
rect 26016 22040 26022 22052
rect 26053 22049 26065 22052
rect 26099 22049 26111 22083
rect 26053 22043 26111 22049
rect 26694 22040 26700 22092
rect 26752 22080 26758 22092
rect 27338 22080 27344 22092
rect 26752 22052 27344 22080
rect 26752 22040 26758 22052
rect 27338 22040 27344 22052
rect 27396 22080 27402 22092
rect 29638 22080 29644 22092
rect 27396 22052 29500 22080
rect 29599 22052 29644 22080
rect 27396 22040 27402 22052
rect 29472 22024 29500 22052
rect 29638 22040 29644 22052
rect 29696 22040 29702 22092
rect 30006 22040 30012 22092
rect 30064 22080 30070 22092
rect 31570 22080 31576 22092
rect 30064 22052 31576 22080
rect 30064 22040 30070 22052
rect 31570 22040 31576 22052
rect 31628 22080 31634 22092
rect 32585 22083 32643 22089
rect 32585 22080 32597 22083
rect 31628 22052 32597 22080
rect 31628 22040 31634 22052
rect 32585 22049 32597 22052
rect 32631 22049 32643 22083
rect 45388 22080 45416 22120
rect 32585 22043 32643 22049
rect 33888 22052 44496 22080
rect 22189 22015 22247 22021
rect 22189 22012 22201 22015
rect 22152 21984 22201 22012
rect 22152 21972 22158 21984
rect 22189 21981 22201 21984
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 23569 22015 23627 22021
rect 23569 22012 23581 22015
rect 22833 21975 22891 21981
rect 23400 21984 23581 22012
rect 20898 21944 20904 21956
rect 19996 21916 20904 21944
rect 19116 21904 19122 21916
rect 20898 21904 20904 21916
rect 20956 21904 20962 21956
rect 21174 21944 21180 21956
rect 21087 21916 21180 21944
rect 21174 21904 21180 21916
rect 21232 21944 21238 21956
rect 23290 21944 23296 21956
rect 21232 21916 23296 21944
rect 21232 21904 21238 21916
rect 23290 21904 23296 21916
rect 23348 21904 23354 21956
rect 11606 21836 11612 21888
rect 11664 21876 11670 21888
rect 11882 21876 11888 21888
rect 11664 21848 11888 21876
rect 11664 21836 11670 21848
rect 11882 21836 11888 21848
rect 11940 21876 11946 21888
rect 12989 21879 13047 21885
rect 12989 21876 13001 21879
rect 11940 21848 13001 21876
rect 11940 21836 11946 21848
rect 12989 21845 13001 21848
rect 13035 21845 13047 21879
rect 12989 21839 13047 21845
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13964 21848 14289 21876
rect 13964 21836 13970 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 16206 21876 16212 21888
rect 16167 21848 16212 21876
rect 14277 21839 14335 21845
rect 16206 21836 16212 21848
rect 16264 21836 16270 21888
rect 20530 21836 20536 21888
rect 20588 21876 20594 21888
rect 20625 21879 20683 21885
rect 20625 21876 20637 21879
rect 20588 21848 20637 21876
rect 20588 21836 20594 21848
rect 20625 21845 20637 21848
rect 20671 21845 20683 21879
rect 20625 21839 20683 21845
rect 20806 21836 20812 21888
rect 20864 21876 20870 21888
rect 21361 21879 21419 21885
rect 21361 21876 21373 21879
rect 20864 21848 21373 21876
rect 20864 21836 20870 21848
rect 21361 21845 21373 21848
rect 21407 21845 21419 21879
rect 21361 21839 21419 21845
rect 22097 21879 22155 21885
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22554 21876 22560 21888
rect 22143 21848 22560 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22554 21836 22560 21848
rect 22612 21836 22618 21888
rect 23017 21879 23075 21885
rect 23017 21845 23029 21879
rect 23063 21876 23075 21879
rect 23400 21876 23428 21984
rect 23569 21981 23581 21984
rect 23615 22012 23627 22015
rect 25409 22015 25467 22021
rect 25409 22012 25421 22015
rect 23615 21984 25421 22012
rect 23615 21981 23627 21984
rect 23569 21975 23627 21981
rect 25409 21981 25421 21984
rect 25455 22012 25467 22015
rect 25455 21984 26004 22012
rect 25455 21981 25467 21984
rect 25409 21975 25467 21981
rect 23658 21876 23664 21888
rect 23063 21848 23428 21876
rect 23619 21848 23664 21876
rect 23063 21845 23075 21848
rect 23017 21839 23075 21845
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 25498 21876 25504 21888
rect 25459 21848 25504 21876
rect 25498 21836 25504 21848
rect 25556 21836 25562 21888
rect 25976 21876 26004 21984
rect 28166 21972 28172 22024
rect 28224 22012 28230 22024
rect 28721 22015 28779 22021
rect 28721 22012 28733 22015
rect 28224 21984 28733 22012
rect 28224 21972 28230 21984
rect 28721 21981 28733 21984
rect 28767 22012 28779 22015
rect 29178 22012 29184 22024
rect 28767 21984 29184 22012
rect 28767 21981 28779 21984
rect 28721 21975 28779 21981
rect 29178 21972 29184 21984
rect 29236 21972 29242 22024
rect 29454 21972 29460 22024
rect 29512 22012 29518 22024
rect 29549 22015 29607 22021
rect 29549 22012 29561 22015
rect 29512 21984 29561 22012
rect 29512 21972 29518 21984
rect 29549 21981 29561 21984
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 26326 21944 26332 21956
rect 26287 21916 26332 21944
rect 26326 21904 26332 21916
rect 26384 21904 26390 21956
rect 27062 21904 27068 21956
rect 27120 21904 27126 21956
rect 28353 21947 28411 21953
rect 28353 21944 28365 21947
rect 27816 21916 28365 21944
rect 26694 21876 26700 21888
rect 25976 21848 26700 21876
rect 26694 21836 26700 21848
rect 26752 21836 26758 21888
rect 27154 21836 27160 21888
rect 27212 21876 27218 21888
rect 27816 21885 27844 21916
rect 28353 21913 28365 21916
rect 28399 21913 28411 21947
rect 28353 21907 28411 21913
rect 28537 21947 28595 21953
rect 28537 21913 28549 21947
rect 28583 21944 28595 21947
rect 28994 21944 29000 21956
rect 28583 21916 29000 21944
rect 28583 21913 28595 21916
rect 28537 21907 28595 21913
rect 28994 21904 29000 21916
rect 29052 21904 29058 21956
rect 32309 21947 32367 21953
rect 32309 21913 32321 21947
rect 32355 21913 32367 21947
rect 32309 21907 32367 21913
rect 27801 21879 27859 21885
rect 27801 21876 27813 21879
rect 27212 21848 27813 21876
rect 27212 21836 27218 21848
rect 27801 21845 27813 21848
rect 27847 21845 27859 21879
rect 27801 21839 27859 21845
rect 28629 21879 28687 21885
rect 28629 21845 28641 21879
rect 28675 21876 28687 21879
rect 28718 21876 28724 21888
rect 28675 21848 28724 21876
rect 28675 21845 28687 21848
rect 28629 21839 28687 21845
rect 28718 21836 28724 21848
rect 28776 21876 28782 21888
rect 29086 21876 29092 21888
rect 28776 21848 29092 21876
rect 28776 21836 28782 21848
rect 29086 21836 29092 21848
rect 29144 21836 29150 21888
rect 32324 21876 32352 21907
rect 32398 21904 32404 21956
rect 32456 21944 32462 21956
rect 32456 21916 32501 21944
rect 32456 21904 32462 21916
rect 33888 21876 33916 22052
rect 33962 21972 33968 22024
rect 34020 22012 34026 22024
rect 34149 22015 34207 22021
rect 34149 22012 34161 22015
rect 34020 21984 34161 22012
rect 34020 21972 34026 21984
rect 34149 21981 34161 21984
rect 34195 21981 34207 22015
rect 40034 22012 40040 22024
rect 39995 21984 40040 22012
rect 34149 21975 34207 21981
rect 40034 21972 40040 21984
rect 40092 21972 40098 22024
rect 41141 22015 41199 22021
rect 41141 21981 41153 22015
rect 41187 21981 41199 22015
rect 43162 22012 43168 22024
rect 43123 21984 43168 22012
rect 41141 21975 41199 21981
rect 34054 21904 34060 21956
rect 34112 21944 34118 21956
rect 34793 21947 34851 21953
rect 34793 21944 34805 21947
rect 34112 21916 34805 21944
rect 34112 21904 34118 21916
rect 34793 21913 34805 21916
rect 34839 21913 34851 21947
rect 34793 21907 34851 21913
rect 34885 21947 34943 21953
rect 34885 21913 34897 21947
rect 34931 21913 34943 21947
rect 35802 21944 35808 21956
rect 35763 21916 35808 21944
rect 34885 21907 34943 21913
rect 32324 21848 33916 21876
rect 33965 21879 34023 21885
rect 33965 21845 33977 21879
rect 34011 21876 34023 21879
rect 34900 21876 34928 21907
rect 35802 21904 35808 21916
rect 35860 21904 35866 21956
rect 41156 21944 41184 21975
rect 43162 21972 43168 21984
rect 43220 21972 43226 22024
rect 43254 21972 43260 22024
rect 43312 22012 43318 22024
rect 43349 22015 43407 22021
rect 43349 22012 43361 22015
rect 43312 21984 43361 22012
rect 43312 21972 43318 21984
rect 43349 21981 43361 21984
rect 43395 21981 43407 22015
rect 43349 21975 43407 21981
rect 43898 21944 43904 21956
rect 40512 21916 41184 21944
rect 43859 21916 43904 21944
rect 40512 21885 40540 21916
rect 43898 21904 43904 21916
rect 43956 21904 43962 21956
rect 43990 21904 43996 21956
rect 44048 21944 44054 21956
rect 44085 21947 44143 21953
rect 44085 21944 44097 21947
rect 44048 21916 44097 21944
rect 44048 21904 44054 21916
rect 44085 21913 44097 21916
rect 44131 21913 44143 21947
rect 44468 21944 44496 22052
rect 45020 22052 45416 22080
rect 45526 22080 45554 22120
rect 47394 22080 47400 22092
rect 45526 22052 47400 22080
rect 45020 22021 45048 22052
rect 47394 22040 47400 22052
rect 47452 22080 47458 22092
rect 47670 22080 47676 22092
rect 47452 22052 47676 22080
rect 47452 22040 47458 22052
rect 47670 22040 47676 22052
rect 47728 22040 47734 22092
rect 45005 22015 45063 22021
rect 45005 21981 45017 22015
rect 45051 21981 45063 22015
rect 45186 22012 45192 22024
rect 45147 21984 45192 22012
rect 45005 21975 45063 21981
rect 45186 21972 45192 21984
rect 45244 21972 45250 22024
rect 45278 21972 45284 22024
rect 45336 22012 45342 22024
rect 45649 22015 45707 22021
rect 45649 22012 45661 22015
rect 45336 21984 45661 22012
rect 45336 21972 45342 21984
rect 45649 21981 45661 21984
rect 45695 21981 45707 22015
rect 45649 21975 45707 21981
rect 48038 21972 48044 22024
rect 48096 22012 48102 22024
rect 48133 22015 48191 22021
rect 48133 22012 48145 22015
rect 48096 21984 48145 22012
rect 48096 21972 48102 21984
rect 48133 21981 48145 21984
rect 48179 21981 48191 22015
rect 48133 21975 48191 21981
rect 45554 21944 45560 21956
rect 44468 21916 45560 21944
rect 44085 21907 44143 21913
rect 45554 21904 45560 21916
rect 45612 21904 45618 21956
rect 45833 21947 45891 21953
rect 45833 21913 45845 21947
rect 45879 21913 45891 21947
rect 45833 21907 45891 21913
rect 34011 21848 34928 21876
rect 40497 21879 40555 21885
rect 34011 21845 34023 21848
rect 33965 21839 34023 21845
rect 40497 21845 40509 21879
rect 40543 21845 40555 21879
rect 44266 21876 44272 21888
rect 44227 21848 44272 21876
rect 40497 21839 40555 21845
rect 44266 21836 44272 21848
rect 44324 21836 44330 21888
rect 45189 21879 45247 21885
rect 45189 21845 45201 21879
rect 45235 21876 45247 21879
rect 45462 21876 45468 21888
rect 45235 21848 45468 21876
rect 45235 21845 45247 21848
rect 45189 21839 45247 21845
rect 45462 21836 45468 21848
rect 45520 21836 45526 21888
rect 45848 21876 45876 21907
rect 47118 21904 47124 21956
rect 47176 21944 47182 21956
rect 47489 21947 47547 21953
rect 47489 21944 47501 21947
rect 47176 21916 47501 21944
rect 47176 21904 47182 21916
rect 47489 21913 47501 21916
rect 47535 21913 47547 21947
rect 47489 21907 47547 21913
rect 47949 21879 48007 21885
rect 47949 21876 47961 21879
rect 45848 21848 47961 21876
rect 47949 21845 47961 21848
rect 47995 21845 48007 21879
rect 47949 21839 48007 21845
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12158 21672 12164 21684
rect 11931 21644 12164 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 12647 21675 12705 21681
rect 12647 21641 12659 21675
rect 12693 21672 12705 21675
rect 12894 21672 12900 21684
rect 12693 21644 12900 21672
rect 12693 21641 12705 21644
rect 12647 21635 12705 21641
rect 12894 21632 12900 21644
rect 12952 21632 12958 21684
rect 16025 21675 16083 21681
rect 16025 21641 16037 21675
rect 16071 21672 16083 21675
rect 17034 21672 17040 21684
rect 16071 21644 17040 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 19521 21675 19579 21681
rect 19521 21672 19533 21675
rect 19392 21644 19533 21672
rect 19392 21632 19398 21644
rect 19521 21641 19533 21644
rect 19567 21641 19579 21675
rect 19521 21635 19579 21641
rect 19978 21632 19984 21684
rect 20036 21672 20042 21684
rect 20165 21675 20223 21681
rect 20165 21672 20177 21675
rect 20036 21644 20177 21672
rect 20036 21632 20042 21644
rect 20165 21641 20177 21644
rect 20211 21641 20223 21675
rect 20165 21635 20223 21641
rect 20993 21675 21051 21681
rect 20993 21641 21005 21675
rect 21039 21672 21051 21675
rect 21266 21672 21272 21684
rect 21039 21644 21272 21672
rect 21039 21641 21051 21644
rect 20993 21635 21051 21641
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 21726 21632 21732 21684
rect 21784 21672 21790 21684
rect 21784 21644 31754 21672
rect 21784 21632 21790 21644
rect 11422 21604 11428 21616
rect 8312 21576 11428 21604
rect 8312 21545 8340 21576
rect 11422 21564 11428 21576
rect 11480 21564 11486 21616
rect 12434 21604 12440 21616
rect 11808 21576 12440 21604
rect 8297 21539 8355 21545
rect 8297 21505 8309 21539
rect 8343 21505 8355 21539
rect 11698 21536 11704 21548
rect 11611 21508 11704 21536
rect 8297 21499 8355 21505
rect 11698 21496 11704 21508
rect 11756 21536 11762 21548
rect 11808 21536 11836 21576
rect 12434 21564 12440 21576
rect 12492 21604 12498 21616
rect 20717 21607 20775 21613
rect 12492 21576 12537 21604
rect 12492 21564 12498 21576
rect 20717 21573 20729 21607
rect 20763 21604 20775 21607
rect 21174 21604 21180 21616
rect 20763 21576 21180 21604
rect 20763 21573 20775 21576
rect 20717 21567 20775 21573
rect 21174 21564 21180 21576
rect 21232 21564 21238 21616
rect 22554 21604 22560 21616
rect 22515 21576 22560 21604
rect 22554 21564 22560 21576
rect 22612 21564 22618 21616
rect 25498 21564 25504 21616
rect 25556 21564 25562 21616
rect 27985 21607 28043 21613
rect 27985 21573 27997 21607
rect 28031 21573 28043 21607
rect 27985 21567 28043 21573
rect 11756 21508 11836 21536
rect 11756 21496 11762 21508
rect 11882 21496 11888 21548
rect 11940 21536 11946 21548
rect 11977 21539 12035 21545
rect 11977 21536 11989 21539
rect 11940 21508 11989 21536
rect 11940 21496 11946 21508
rect 11977 21505 11989 21508
rect 12023 21536 12035 21539
rect 12342 21536 12348 21548
rect 12023 21508 12348 21536
rect 12023 21505 12035 21508
rect 11977 21499 12035 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21505 13783 21539
rect 14918 21536 14924 21548
rect 14879 21508 14924 21536
rect 13725 21499 13783 21505
rect 8481 21471 8539 21477
rect 8481 21437 8493 21471
rect 8527 21468 8539 21471
rect 9030 21468 9036 21480
rect 8527 21440 9036 21468
rect 8527 21437 8539 21440
rect 8481 21431 8539 21437
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 9125 21471 9183 21477
rect 9125 21437 9137 21471
rect 9171 21437 9183 21471
rect 13740 21468 13768 21499
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21536 15991 21539
rect 16206 21536 16212 21548
rect 15979 21508 16212 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 15948 21468 15976 21499
rect 16206 21496 16212 21508
rect 16264 21496 16270 21548
rect 17310 21536 17316 21548
rect 17271 21508 17316 21536
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18141 21539 18199 21545
rect 18141 21536 18153 21539
rect 18012 21508 18153 21536
rect 18012 21496 18018 21508
rect 18141 21505 18153 21508
rect 18187 21505 18199 21539
rect 19426 21536 19432 21548
rect 19387 21508 19432 21536
rect 18141 21499 18199 21505
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 20070 21536 20076 21548
rect 20031 21508 20076 21536
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21505 20315 21539
rect 20257 21499 20315 21505
rect 9125 21431 9183 21437
rect 11348 21440 15976 21468
rect 17405 21471 17463 21477
rect 7926 21360 7932 21412
rect 7984 21400 7990 21412
rect 9140 21400 9168 21431
rect 7984 21372 9168 21400
rect 7984 21360 7990 21372
rect 8938 21292 8944 21344
rect 8996 21332 9002 21344
rect 11348 21332 11376 21440
rect 17405 21437 17417 21471
rect 17451 21468 17463 21471
rect 18230 21468 18236 21480
rect 17451 21440 18236 21468
rect 17451 21437 17463 21440
rect 17405 21431 17463 21437
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 18417 21471 18475 21477
rect 18417 21437 18429 21471
rect 18463 21468 18475 21471
rect 18598 21468 18604 21480
rect 18463 21440 18604 21468
rect 18463 21437 18475 21440
rect 18417 21431 18475 21437
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 20272 21468 20300 21499
rect 20806 21496 20812 21548
rect 20864 21536 20870 21548
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20864 21508 20913 21536
rect 20864 21496 20870 21508
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21505 21143 21539
rect 21085 21499 21143 21505
rect 20530 21468 20536 21480
rect 20272 21440 20536 21468
rect 20530 21428 20536 21440
rect 20588 21468 20594 21480
rect 20990 21468 20996 21480
rect 20588 21440 20996 21468
rect 20588 21428 20594 21440
rect 20990 21428 20996 21440
rect 21048 21428 21054 21480
rect 12802 21400 12808 21412
rect 12763 21372 12808 21400
rect 12802 21360 12808 21372
rect 12860 21360 12866 21412
rect 14090 21360 14096 21412
rect 14148 21400 14154 21412
rect 14148 21372 18368 21400
rect 14148 21360 14154 21372
rect 11514 21332 11520 21344
rect 8996 21304 11376 21332
rect 11475 21304 11520 21332
rect 8996 21292 9002 21304
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 12158 21292 12164 21344
rect 12216 21332 12222 21344
rect 12621 21335 12679 21341
rect 12621 21332 12633 21335
rect 12216 21304 12633 21332
rect 12216 21292 12222 21304
rect 12621 21301 12633 21304
rect 12667 21301 12679 21335
rect 12621 21295 12679 21301
rect 13817 21335 13875 21341
rect 13817 21301 13829 21335
rect 13863 21332 13875 21335
rect 14274 21332 14280 21344
rect 13863 21304 14280 21332
rect 13863 21301 13875 21304
rect 13817 21295 13875 21301
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 15105 21335 15163 21341
rect 15105 21332 15117 21335
rect 14424 21304 15117 21332
rect 14424 21292 14430 21304
rect 15105 21301 15117 21304
rect 15151 21301 15163 21335
rect 15105 21295 15163 21301
rect 17681 21335 17739 21341
rect 17681 21301 17693 21335
rect 17727 21332 17739 21335
rect 18230 21332 18236 21344
rect 17727 21304 18236 21332
rect 17727 21301 17739 21304
rect 17681 21295 17739 21301
rect 18230 21292 18236 21304
rect 18288 21292 18294 21344
rect 18340 21332 18368 21372
rect 20622 21360 20628 21412
rect 20680 21400 20686 21412
rect 21100 21400 21128 21499
rect 23658 21496 23664 21548
rect 23716 21496 23722 21548
rect 27154 21536 27160 21548
rect 27115 21508 27160 21536
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 28000 21536 28028 21567
rect 28166 21564 28172 21616
rect 28224 21613 28230 21616
rect 28224 21607 28243 21613
rect 28231 21573 28243 21607
rect 28224 21567 28243 21573
rect 28224 21564 28230 21567
rect 28718 21564 28724 21616
rect 28776 21604 28782 21616
rect 28776 21576 29040 21604
rect 28776 21564 28782 21576
rect 28552 21536 28672 21542
rect 28813 21539 28871 21545
rect 28813 21536 28825 21539
rect 28000 21514 28825 21536
rect 28000 21508 28580 21514
rect 28644 21508 28825 21514
rect 28813 21505 28825 21508
rect 28859 21536 28871 21539
rect 28902 21536 28908 21548
rect 28859 21508 28908 21536
rect 28859 21505 28871 21508
rect 28813 21499 28871 21505
rect 28902 21496 28908 21508
rect 28960 21496 28966 21548
rect 29012 21545 29040 21576
rect 29178 21570 29184 21616
rect 29104 21567 29184 21570
rect 29089 21564 29184 21567
rect 29236 21564 29242 21616
rect 30282 21564 30288 21616
rect 30340 21604 30346 21616
rect 30653 21607 30711 21613
rect 30653 21604 30665 21607
rect 30340 21576 30665 21604
rect 30340 21564 30346 21576
rect 30653 21573 30665 21576
rect 30699 21604 30711 21607
rect 31570 21604 31576 21616
rect 30699 21576 31432 21604
rect 31531 21576 31576 21604
rect 30699 21573 30711 21576
rect 30653 21567 30711 21573
rect 29089 21561 29224 21564
rect 28997 21539 29055 21545
rect 28997 21505 29009 21539
rect 29043 21505 29055 21539
rect 29089 21527 29101 21561
rect 29135 21542 29224 21561
rect 29135 21527 29147 21542
rect 29089 21521 29147 21527
rect 29549 21539 29607 21545
rect 28997 21499 29055 21505
rect 29549 21505 29561 21539
rect 29595 21505 29607 21539
rect 29730 21536 29736 21548
rect 29691 21508 29736 21536
rect 29549 21499 29607 21505
rect 22278 21468 22284 21480
rect 22239 21440 22284 21468
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 23290 21428 23296 21480
rect 23348 21468 23354 21480
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23348 21440 24041 21468
rect 23348 21428 23354 21440
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 24118 21428 24124 21480
rect 24176 21468 24182 21480
rect 24489 21471 24547 21477
rect 24489 21468 24501 21471
rect 24176 21440 24501 21468
rect 24176 21428 24182 21440
rect 24489 21437 24501 21440
rect 24535 21437 24547 21471
rect 24489 21431 24547 21437
rect 24765 21471 24823 21477
rect 24765 21437 24777 21471
rect 24811 21468 24823 21471
rect 25314 21468 25320 21480
rect 24811 21440 25320 21468
rect 24811 21437 24823 21440
rect 24765 21431 24823 21437
rect 25314 21428 25320 21440
rect 25372 21428 25378 21480
rect 27249 21471 27307 21477
rect 27249 21437 27261 21471
rect 27295 21468 27307 21471
rect 27295 21440 28396 21468
rect 27295 21437 27307 21440
rect 27249 21431 27307 21437
rect 28368 21412 28396 21440
rect 20680 21372 21128 21400
rect 21192 21372 21588 21400
rect 20680 21360 20686 21372
rect 21192 21332 21220 21372
rect 18340 21304 21220 21332
rect 21269 21335 21327 21341
rect 21269 21301 21281 21335
rect 21315 21332 21327 21335
rect 21450 21332 21456 21344
rect 21315 21304 21456 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 21450 21292 21456 21304
rect 21508 21292 21514 21344
rect 21560 21332 21588 21372
rect 26326 21360 26332 21412
rect 26384 21400 26390 21412
rect 27525 21403 27583 21409
rect 27525 21400 27537 21403
rect 26384 21372 27537 21400
rect 26384 21360 26390 21372
rect 27525 21369 27537 21372
rect 27571 21369 27583 21403
rect 28350 21400 28356 21412
rect 28311 21372 28356 21400
rect 27525 21363 27583 21369
rect 28350 21360 28356 21372
rect 28408 21360 28414 21412
rect 28813 21403 28871 21409
rect 28813 21369 28825 21403
rect 28859 21400 28871 21403
rect 29564 21400 29592 21499
rect 29730 21496 29736 21508
rect 29788 21496 29794 21548
rect 31404 21536 31432 21576
rect 31570 21564 31576 21576
rect 31628 21564 31634 21616
rect 31726 21604 31754 21644
rect 32398 21632 32404 21684
rect 32456 21672 32462 21684
rect 33045 21675 33103 21681
rect 33045 21672 33057 21675
rect 32456 21644 33057 21672
rect 32456 21632 32462 21644
rect 33045 21641 33057 21644
rect 33091 21641 33103 21675
rect 33962 21672 33968 21684
rect 33923 21644 33968 21672
rect 33045 21635 33103 21641
rect 33962 21632 33968 21644
rect 34020 21632 34026 21684
rect 42702 21672 42708 21684
rect 34992 21644 42708 21672
rect 34992 21604 35020 21644
rect 42702 21632 42708 21644
rect 42760 21632 42766 21684
rect 46106 21672 46112 21684
rect 43180 21644 46112 21672
rect 31726 21576 35020 21604
rect 35066 21564 35072 21616
rect 35124 21604 35130 21616
rect 36354 21604 36360 21616
rect 35124 21576 36360 21604
rect 35124 21564 35130 21576
rect 36354 21564 36360 21576
rect 36412 21564 36418 21616
rect 38378 21564 38384 21616
rect 38436 21604 38442 21616
rect 43180 21604 43208 21644
rect 46106 21632 46112 21644
rect 46164 21632 46170 21684
rect 47762 21632 47768 21684
rect 47820 21672 47826 21684
rect 48133 21675 48191 21681
rect 48133 21672 48145 21675
rect 47820 21644 48145 21672
rect 47820 21632 47826 21644
rect 48133 21641 48145 21644
rect 48179 21641 48191 21675
rect 48133 21635 48191 21641
rect 38436 21576 43208 21604
rect 45005 21607 45063 21613
rect 38436 21564 38442 21576
rect 45005 21573 45017 21607
rect 45051 21604 45063 21607
rect 45094 21604 45100 21616
rect 45051 21576 45100 21604
rect 45051 21573 45063 21576
rect 45005 21567 45063 21573
rect 45094 21564 45100 21576
rect 45152 21564 45158 21616
rect 45186 21564 45192 21616
rect 45244 21604 45250 21616
rect 47670 21604 47676 21616
rect 45244 21576 47676 21604
rect 45244 21564 45250 21576
rect 47670 21564 47676 21576
rect 47728 21564 47734 21616
rect 32125 21539 32183 21545
rect 32125 21536 32137 21539
rect 31404 21508 32137 21536
rect 32125 21505 32137 21508
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 33229 21539 33287 21545
rect 33229 21505 33241 21539
rect 33275 21505 33287 21539
rect 33229 21499 33287 21505
rect 34425 21539 34483 21545
rect 34425 21505 34437 21539
rect 34471 21536 34483 21539
rect 34790 21536 34796 21548
rect 34471 21508 34796 21536
rect 34471 21505 34483 21508
rect 34425 21499 34483 21505
rect 30561 21471 30619 21477
rect 30561 21437 30573 21471
rect 30607 21437 30619 21471
rect 30561 21431 30619 21437
rect 32585 21471 32643 21477
rect 32585 21437 32597 21471
rect 32631 21468 32643 21471
rect 33244 21468 33272 21499
rect 34790 21496 34796 21508
rect 34848 21496 34854 21548
rect 39942 21536 39948 21548
rect 39903 21508 39948 21536
rect 39942 21496 39948 21508
rect 40000 21496 40006 21548
rect 40126 21536 40132 21548
rect 40087 21508 40132 21536
rect 40126 21496 40132 21508
rect 40184 21496 40190 21548
rect 42886 21496 42892 21548
rect 42944 21536 42950 21548
rect 43165 21539 43223 21545
rect 43165 21536 43177 21539
rect 42944 21508 43177 21536
rect 42944 21496 42950 21508
rect 43165 21505 43177 21508
rect 43211 21536 43223 21539
rect 43254 21536 43260 21548
rect 43211 21508 43260 21536
rect 43211 21505 43223 21508
rect 43165 21499 43223 21505
rect 43254 21496 43260 21508
rect 43312 21496 43318 21548
rect 43349 21539 43407 21545
rect 43349 21505 43361 21539
rect 43395 21536 43407 21539
rect 43530 21536 43536 21548
rect 43395 21508 43536 21536
rect 43395 21505 43407 21508
rect 43349 21499 43407 21505
rect 43530 21496 43536 21508
rect 43588 21496 43594 21548
rect 44174 21496 44180 21548
rect 44232 21536 44238 21548
rect 44269 21539 44327 21545
rect 44269 21536 44281 21539
rect 44232 21508 44281 21536
rect 44232 21496 44238 21508
rect 44269 21505 44281 21508
rect 44315 21505 44327 21539
rect 44269 21499 44327 21505
rect 44542 21496 44548 21548
rect 44600 21496 44606 21548
rect 46198 21536 46204 21548
rect 46159 21508 46204 21536
rect 46198 21496 46204 21508
rect 46256 21496 46262 21548
rect 47026 21536 47032 21548
rect 46308 21508 47032 21536
rect 34977 21471 35035 21477
rect 34977 21468 34989 21471
rect 32631 21440 33272 21468
rect 33336 21440 34989 21468
rect 32631 21437 32643 21440
rect 32585 21431 32643 21437
rect 28859 21372 29592 21400
rect 30576 21400 30604 21431
rect 30576 21372 32628 21400
rect 28859 21369 28871 21372
rect 28813 21363 28871 21369
rect 22002 21332 22008 21344
rect 21560 21304 22008 21332
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 26234 21332 26240 21344
rect 26195 21304 26240 21332
rect 26234 21292 26240 21304
rect 26292 21332 26298 21344
rect 28169 21335 28227 21341
rect 28169 21332 28181 21335
rect 26292 21304 28181 21332
rect 26292 21292 26298 21304
rect 28169 21301 28181 21304
rect 28215 21332 28227 21335
rect 28718 21332 28724 21344
rect 28215 21304 28724 21332
rect 28215 21301 28227 21304
rect 28169 21295 28227 21301
rect 28718 21292 28724 21304
rect 28776 21292 28782 21344
rect 28994 21292 29000 21344
rect 29052 21332 29058 21344
rect 29549 21335 29607 21341
rect 29549 21332 29561 21335
rect 29052 21304 29561 21332
rect 29052 21292 29058 21304
rect 29549 21301 29561 21304
rect 29595 21301 29607 21335
rect 32398 21332 32404 21344
rect 32359 21304 32404 21332
rect 29549 21295 29607 21301
rect 32398 21292 32404 21304
rect 32456 21292 32462 21344
rect 32600 21332 32628 21372
rect 33336 21332 33364 21440
rect 34977 21437 34989 21440
rect 35023 21437 35035 21471
rect 35802 21468 35808 21480
rect 35715 21440 35808 21468
rect 34977 21431 35035 21437
rect 33594 21332 33600 21344
rect 32600 21304 33364 21332
rect 33555 21304 33600 21332
rect 33594 21292 33600 21304
rect 33652 21332 33658 21344
rect 34149 21335 34207 21341
rect 34149 21332 34161 21335
rect 33652 21304 34161 21332
rect 33652 21292 33658 21304
rect 34149 21301 34161 21304
rect 34195 21301 34207 21335
rect 34992 21332 35020 21431
rect 35802 21428 35808 21440
rect 35860 21468 35866 21480
rect 43898 21468 43904 21480
rect 35860 21440 43904 21468
rect 35860 21428 35866 21440
rect 43898 21428 43904 21440
rect 43956 21428 43962 21480
rect 44450 21428 44456 21480
rect 44508 21468 44514 21480
rect 46308 21468 46336 21508
rect 47026 21496 47032 21508
rect 47084 21496 47090 21548
rect 47578 21536 47584 21548
rect 47539 21508 47584 21536
rect 47578 21496 47584 21508
rect 47636 21496 47642 21548
rect 46474 21468 46480 21480
rect 44508 21440 46336 21468
rect 46435 21440 46480 21468
rect 44508 21428 44514 21440
rect 46474 21428 46480 21440
rect 46532 21428 46538 21480
rect 47854 21468 47860 21480
rect 47815 21440 47860 21468
rect 47854 21428 47860 21440
rect 47912 21428 47918 21480
rect 36998 21360 37004 21412
rect 37056 21400 37062 21412
rect 46014 21400 46020 21412
rect 37056 21372 46020 21400
rect 37056 21360 37062 21372
rect 46014 21360 46020 21372
rect 46072 21360 46078 21412
rect 38378 21332 38384 21344
rect 34992 21304 38384 21332
rect 34149 21295 34207 21301
rect 38378 21292 38384 21304
rect 38436 21292 38442 21344
rect 40037 21335 40095 21341
rect 40037 21301 40049 21335
rect 40083 21332 40095 21335
rect 40126 21332 40132 21344
rect 40083 21304 40132 21332
rect 40083 21301 40095 21304
rect 40037 21295 40095 21301
rect 40126 21292 40132 21304
rect 40184 21292 40190 21344
rect 43165 21335 43223 21341
rect 43165 21301 43177 21335
rect 43211 21332 43223 21335
rect 43622 21332 43628 21344
rect 43211 21304 43628 21332
rect 43211 21301 43223 21304
rect 43165 21295 43223 21301
rect 43622 21292 43628 21304
rect 43680 21292 43686 21344
rect 45462 21292 45468 21344
rect 45520 21332 45526 21344
rect 47673 21335 47731 21341
rect 47673 21332 47685 21335
rect 45520 21304 47685 21332
rect 45520 21292 45526 21304
rect 47673 21301 47685 21304
rect 47719 21301 47731 21335
rect 47673 21295 47731 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 9030 21128 9036 21140
rect 8991 21100 9036 21128
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 11348 21100 17264 21128
rect 2866 21020 2872 21072
rect 2924 21060 2930 21072
rect 11348 21060 11376 21100
rect 11514 21060 11520 21072
rect 2924 21032 11376 21060
rect 11475 21032 11520 21060
rect 2924 21020 2930 21032
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 17236 21060 17264 21100
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 20622 21128 20628 21140
rect 19392 21100 20628 21128
rect 19392 21088 19398 21100
rect 20622 21088 20628 21100
rect 20680 21128 20686 21140
rect 20809 21131 20867 21137
rect 20809 21128 20821 21131
rect 20680 21100 20821 21128
rect 20680 21088 20686 21100
rect 20809 21097 20821 21100
rect 20855 21097 20867 21131
rect 20990 21128 20996 21140
rect 20951 21100 20996 21128
rect 20809 21091 20867 21097
rect 20990 21088 20996 21100
rect 21048 21088 21054 21140
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 22373 21131 22431 21137
rect 22373 21128 22385 21131
rect 22336 21100 22385 21128
rect 22336 21088 22342 21100
rect 22373 21097 22385 21100
rect 22419 21097 22431 21131
rect 25314 21128 25320 21140
rect 25275 21100 25320 21128
rect 22373 21091 22431 21097
rect 25314 21088 25320 21100
rect 25372 21088 25378 21140
rect 31110 21088 31116 21140
rect 31168 21128 31174 21140
rect 46474 21128 46480 21140
rect 31168 21100 46480 21128
rect 31168 21088 31174 21100
rect 46474 21088 46480 21100
rect 46532 21088 46538 21140
rect 47210 21088 47216 21140
rect 47268 21128 47274 21140
rect 47854 21128 47860 21140
rect 47268 21100 47860 21128
rect 47268 21088 47274 21100
rect 47854 21088 47860 21100
rect 47912 21088 47918 21140
rect 33594 21060 33600 21072
rect 11808 21032 14596 21060
rect 17236 21032 33600 21060
rect 11701 20995 11759 21001
rect 11701 20992 11713 20995
rect 10796 20964 11713 20992
rect 8938 20924 8944 20936
rect 8899 20896 8944 20924
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 10796 20933 10824 20964
rect 11701 20961 11713 20964
rect 11747 20961 11759 20995
rect 11701 20955 11759 20961
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20893 10839 20927
rect 11808 20924 11836 21032
rect 14274 20992 14280 21004
rect 14235 20964 14280 20992
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 14568 21001 14596 21032
rect 33594 21020 33600 21032
rect 33652 21020 33658 21072
rect 43165 21063 43223 21069
rect 43165 21029 43177 21063
rect 43211 21060 43223 21063
rect 43714 21060 43720 21072
rect 43211 21032 43720 21060
rect 43211 21029 43223 21032
rect 43165 21023 43223 21029
rect 43714 21020 43720 21032
rect 43772 21020 43778 21072
rect 46934 21060 46940 21072
rect 45664 21032 46940 21060
rect 14553 20995 14611 21001
rect 14553 20961 14565 20995
rect 14599 20961 14611 20995
rect 14553 20955 14611 20961
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20992 16451 20995
rect 17310 20992 17316 21004
rect 16439 20964 17316 20992
rect 16439 20961 16451 20964
rect 16393 20955 16451 20961
rect 17310 20952 17316 20964
rect 17368 20992 17374 21004
rect 17954 20992 17960 21004
rect 17368 20964 17816 20992
rect 17915 20964 17960 20992
rect 17368 20952 17374 20964
rect 14090 20924 14096 20936
rect 10781 20887 10839 20893
rect 11164 20896 11836 20924
rect 14051 20896 14096 20924
rect 14 20816 20 20868
rect 72 20856 78 20868
rect 11164 20856 11192 20896
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 17788 20924 17816 20964
rect 17954 20952 17960 20964
rect 18012 20952 18018 21004
rect 21450 20992 21456 21004
rect 21411 20964 21456 20992
rect 21450 20952 21456 20964
rect 21508 20952 21514 21004
rect 21821 20995 21879 21001
rect 21821 20961 21833 20995
rect 21867 20992 21879 20995
rect 22094 20992 22100 21004
rect 21867 20964 22100 20992
rect 21867 20961 21879 20964
rect 21821 20955 21879 20961
rect 22094 20952 22100 20964
rect 22152 20992 22158 21004
rect 24857 20995 24915 21001
rect 24857 20992 24869 20995
rect 22152 20964 24869 20992
rect 22152 20952 22158 20964
rect 24857 20961 24869 20964
rect 24903 20992 24915 20995
rect 28166 20992 28172 21004
rect 24903 20964 28172 20992
rect 24903 20961 24915 20964
rect 24857 20955 24915 20961
rect 28166 20952 28172 20964
rect 28224 20952 28230 21004
rect 28534 20952 28540 21004
rect 28592 20992 28598 21004
rect 34054 20992 34060 21004
rect 28592 20964 32536 20992
rect 28592 20952 28598 20964
rect 19334 20924 19340 20936
rect 17788 20896 19340 20924
rect 19334 20884 19340 20896
rect 19392 20884 19398 20936
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19484 20896 19577 20924
rect 19484 20884 19490 20896
rect 21358 20884 21364 20936
rect 21416 20924 21422 20936
rect 21637 20927 21695 20933
rect 21637 20924 21649 20927
rect 21416 20896 21649 20924
rect 21416 20884 21422 20896
rect 21637 20893 21649 20896
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20893 22615 20927
rect 22557 20887 22615 20893
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 23198 20924 23204 20936
rect 23155 20896 23204 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 72 20828 11192 20856
rect 11241 20859 11299 20865
rect 72 20816 78 20828
rect 11241 20825 11253 20859
rect 11287 20856 11299 20859
rect 12802 20856 12808 20868
rect 11287 20828 12808 20856
rect 11287 20825 11299 20828
rect 11241 20819 11299 20825
rect 12802 20816 12808 20828
rect 12860 20816 12866 20868
rect 16574 20856 16580 20868
rect 16535 20828 16580 20856
rect 16574 20816 16580 20828
rect 16632 20816 16638 20868
rect 19242 20816 19248 20868
rect 19300 20856 19306 20868
rect 19444 20856 19472 20884
rect 20625 20859 20683 20865
rect 19300 20828 20576 20856
rect 19300 20816 19306 20828
rect 10597 20791 10655 20797
rect 10597 20757 10609 20791
rect 10643 20788 10655 20791
rect 11790 20788 11796 20800
rect 10643 20760 11796 20788
rect 10643 20757 10655 20760
rect 10597 20751 10655 20757
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 19484 20760 19625 20788
rect 19484 20748 19490 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 20548 20788 20576 20828
rect 20625 20825 20637 20859
rect 20671 20856 20683 20859
rect 20714 20856 20720 20868
rect 20671 20828 20720 20856
rect 20671 20825 20683 20828
rect 20625 20819 20683 20825
rect 20714 20816 20720 20828
rect 20772 20816 20778 20868
rect 20841 20859 20899 20865
rect 20841 20825 20853 20859
rect 20887 20856 20899 20859
rect 20990 20856 20996 20868
rect 20887 20828 20996 20856
rect 20887 20825 20899 20828
rect 20841 20819 20899 20825
rect 20990 20816 20996 20828
rect 21048 20816 21054 20868
rect 22572 20856 22600 20887
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 26234 20924 26240 20936
rect 24995 20896 26240 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 28258 20924 28264 20936
rect 28219 20896 28264 20924
rect 28258 20884 28264 20896
rect 28316 20884 28322 20936
rect 29454 20884 29460 20936
rect 29512 20924 29518 20936
rect 29549 20927 29607 20933
rect 29549 20924 29561 20927
rect 29512 20896 29561 20924
rect 29512 20884 29518 20896
rect 29549 20893 29561 20896
rect 29595 20893 29607 20927
rect 29549 20887 29607 20893
rect 30374 20884 30380 20936
rect 30432 20924 30438 20936
rect 30837 20927 30895 20933
rect 30837 20924 30849 20927
rect 30432 20896 30849 20924
rect 30432 20884 30438 20896
rect 30837 20893 30849 20896
rect 30883 20893 30895 20927
rect 32508 20924 32536 20964
rect 32784 20964 34060 20992
rect 32784 20924 32812 20964
rect 34054 20952 34060 20964
rect 34112 20952 34118 21004
rect 43254 20992 43260 21004
rect 42536 20964 43260 20992
rect 33134 20924 33140 20936
rect 32508 20896 32812 20924
rect 33095 20896 33140 20924
rect 30837 20887 30895 20893
rect 33134 20884 33140 20896
rect 33192 20884 33198 20936
rect 42536 20933 42564 20964
rect 43254 20952 43260 20964
rect 43312 20952 43318 21004
rect 43346 20952 43352 21004
rect 43404 20992 43410 21004
rect 43622 20992 43628 21004
rect 43404 20964 43449 20992
rect 43583 20964 43628 20992
rect 43404 20952 43410 20964
rect 43622 20952 43628 20964
rect 43680 20952 43686 21004
rect 42521 20927 42579 20933
rect 42521 20893 42533 20927
rect 42567 20893 42579 20927
rect 42521 20887 42579 20893
rect 42705 20927 42763 20933
rect 42705 20893 42717 20927
rect 42751 20893 42763 20927
rect 43438 20924 43444 20936
rect 43399 20896 43444 20924
rect 42705 20887 42763 20893
rect 28442 20856 28448 20868
rect 22066 20828 23336 20856
rect 28403 20828 28448 20856
rect 22066 20788 22094 20828
rect 23308 20800 23336 20828
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 31018 20856 31024 20868
rect 30979 20828 31024 20856
rect 31018 20816 31024 20828
rect 31076 20816 31082 20868
rect 32677 20859 32735 20865
rect 32677 20825 32689 20859
rect 32723 20856 32735 20859
rect 36998 20856 37004 20868
rect 32723 20828 37004 20856
rect 32723 20825 32735 20828
rect 32677 20819 32735 20825
rect 36998 20816 37004 20828
rect 37056 20816 37062 20868
rect 42720 20856 42748 20887
rect 43438 20884 43444 20896
rect 43496 20884 43502 20936
rect 43533 20927 43591 20933
rect 43533 20893 43545 20927
rect 43579 20893 43591 20927
rect 43533 20887 43591 20893
rect 42978 20856 42984 20868
rect 42720 20828 42984 20856
rect 42978 20816 42984 20828
rect 43036 20856 43042 20868
rect 43548 20856 43576 20887
rect 43898 20884 43904 20936
rect 43956 20924 43962 20936
rect 44177 20927 44235 20933
rect 44177 20924 44189 20927
rect 43956 20896 44189 20924
rect 43956 20884 43962 20896
rect 44177 20893 44189 20896
rect 44223 20893 44235 20927
rect 44177 20887 44235 20893
rect 44361 20927 44419 20933
rect 44361 20893 44373 20927
rect 44407 20893 44419 20927
rect 45462 20924 45468 20936
rect 45423 20896 45468 20924
rect 44361 20887 44419 20893
rect 43036 20828 43576 20856
rect 43036 20816 43042 20828
rect 43990 20816 43996 20868
rect 44048 20856 44054 20868
rect 44376 20856 44404 20887
rect 45462 20884 45468 20896
rect 45520 20884 45526 20936
rect 45664 20933 45692 21032
rect 46934 21020 46940 21032
rect 46992 21060 46998 21072
rect 47578 21060 47584 21072
rect 46992 21032 47584 21060
rect 46992 21020 46998 21032
rect 47578 21020 47584 21032
rect 47636 21020 47642 21072
rect 46293 20995 46351 21001
rect 46293 20961 46305 20995
rect 46339 20992 46351 20995
rect 47854 20992 47860 21004
rect 46339 20964 47860 20992
rect 46339 20961 46351 20964
rect 46293 20955 46351 20961
rect 47854 20952 47860 20964
rect 47912 20952 47918 21004
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 45649 20927 45707 20933
rect 45649 20893 45661 20927
rect 45695 20893 45707 20927
rect 45649 20887 45707 20893
rect 46474 20856 46480 20868
rect 44048 20828 44404 20856
rect 46435 20828 46480 20856
rect 44048 20816 44054 20828
rect 46474 20816 46480 20828
rect 46532 20816 46538 20868
rect 23290 20788 23296 20800
rect 20548 20760 22094 20788
rect 23251 20760 23296 20788
rect 19613 20751 19671 20757
rect 23290 20748 23296 20760
rect 23348 20748 23354 20800
rect 29641 20791 29699 20797
rect 29641 20757 29653 20791
rect 29687 20788 29699 20791
rect 29730 20788 29736 20800
rect 29687 20760 29736 20788
rect 29687 20757 29699 20760
rect 29641 20751 29699 20757
rect 29730 20748 29736 20760
rect 29788 20748 29794 20800
rect 33226 20788 33232 20800
rect 33187 20760 33232 20788
rect 33226 20748 33232 20760
rect 33284 20748 33290 20800
rect 42705 20791 42763 20797
rect 42705 20757 42717 20791
rect 42751 20788 42763 20791
rect 43070 20788 43076 20800
rect 42751 20760 43076 20788
rect 42751 20757 42763 20760
rect 42705 20751 42763 20757
rect 43070 20748 43076 20760
rect 43128 20748 43134 20800
rect 43438 20748 43444 20800
rect 43496 20788 43502 20800
rect 44082 20788 44088 20800
rect 43496 20760 44088 20788
rect 43496 20748 43502 20760
rect 44082 20748 44088 20760
rect 44140 20788 44146 20800
rect 44269 20791 44327 20797
rect 44269 20788 44281 20791
rect 44140 20760 44281 20788
rect 44140 20748 44146 20760
rect 44269 20757 44281 20760
rect 44315 20757 44327 20791
rect 45830 20788 45836 20800
rect 45791 20760 45836 20788
rect 44269 20751 44327 20757
rect 45830 20748 45836 20760
rect 45888 20748 45894 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 3016 20556 15332 20584
rect 3016 20544 3022 20556
rect 11790 20516 11796 20528
rect 11751 20488 11796 20516
rect 11790 20476 11796 20488
rect 11848 20476 11854 20528
rect 12066 20476 12072 20528
rect 12124 20516 12130 20528
rect 15304 20516 15332 20556
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 16761 20587 16819 20593
rect 16761 20584 16773 20587
rect 16632 20556 16773 20584
rect 16632 20544 16638 20556
rect 16761 20553 16773 20556
rect 16807 20553 16819 20587
rect 16761 20547 16819 20553
rect 19150 20544 19156 20596
rect 19208 20584 19214 20596
rect 21818 20584 21824 20596
rect 19208 20556 21824 20584
rect 19208 20544 19214 20556
rect 21818 20544 21824 20556
rect 21876 20544 21882 20596
rect 23106 20544 23112 20596
rect 23164 20584 23170 20596
rect 23293 20587 23351 20593
rect 23293 20584 23305 20587
rect 23164 20556 23305 20584
rect 23164 20544 23170 20556
rect 23293 20553 23305 20556
rect 23339 20553 23351 20587
rect 45649 20587 45707 20593
rect 23293 20547 23351 20553
rect 26896 20556 45600 20584
rect 17954 20516 17960 20528
rect 12124 20488 12282 20516
rect 15304 20488 17960 20516
rect 12124 20476 12130 20488
rect 17954 20476 17960 20488
rect 18012 20476 18018 20528
rect 18230 20516 18236 20528
rect 18191 20488 18236 20516
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 18966 20476 18972 20528
rect 19024 20476 19030 20528
rect 16206 20408 16212 20460
rect 16264 20448 16270 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16264 20420 16681 20448
rect 16264 20408 16270 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 16816 20420 17325 20448
rect 16816 20408 16822 20420
rect 17313 20417 17325 20420
rect 17359 20448 17371 20451
rect 17862 20448 17868 20460
rect 17359 20420 17868 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 20441 20451 20499 20457
rect 20441 20417 20453 20451
rect 20487 20448 20499 20451
rect 20806 20448 20812 20460
rect 20487 20420 20812 20448
rect 20487 20417 20499 20420
rect 20441 20411 20499 20417
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 21836 20457 21864 20544
rect 22002 20476 22008 20528
rect 22060 20516 22066 20528
rect 24118 20516 24124 20528
rect 22060 20476 22094 20516
rect 24079 20488 24124 20516
rect 24118 20476 24124 20488
rect 24176 20476 24182 20528
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20417 21879 20451
rect 22066 20448 22094 20476
rect 23109 20451 23167 20457
rect 23109 20448 23121 20451
rect 22066 20420 23121 20448
rect 21821 20411 21879 20417
rect 23109 20417 23121 20420
rect 23155 20448 23167 20451
rect 23198 20448 23204 20460
rect 23155 20420 23204 20448
rect 23155 20417 23167 20420
rect 23109 20411 23167 20417
rect 23198 20408 23204 20420
rect 23256 20408 23262 20460
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23845 20451 23903 20457
rect 23845 20448 23857 20451
rect 23348 20420 23857 20448
rect 23348 20408 23354 20420
rect 23845 20417 23857 20420
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 10686 20340 10692 20392
rect 10744 20380 10750 20392
rect 11517 20383 11575 20389
rect 11517 20380 11529 20383
rect 10744 20352 11529 20380
rect 10744 20340 10750 20352
rect 11517 20349 11529 20352
rect 11563 20349 11575 20383
rect 11517 20343 11575 20349
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 13265 20383 13323 20389
rect 13265 20380 13277 20383
rect 12492 20352 13277 20380
rect 12492 20340 12498 20352
rect 13265 20349 13277 20352
rect 13311 20380 13323 20383
rect 14277 20383 14335 20389
rect 14277 20380 14289 20383
rect 13311 20352 14289 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 14277 20349 14289 20352
rect 14323 20349 14335 20383
rect 14277 20343 14335 20349
rect 14461 20383 14519 20389
rect 14461 20349 14473 20383
rect 14507 20380 14519 20383
rect 15470 20380 15476 20392
rect 14507 20352 15476 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 16114 20380 16120 20392
rect 16075 20352 16120 20380
rect 16114 20340 16120 20352
rect 16172 20340 16178 20392
rect 17954 20380 17960 20392
rect 17915 20352 17960 20380
rect 17954 20340 17960 20352
rect 18012 20340 18018 20392
rect 18598 20340 18604 20392
rect 18656 20380 18662 20392
rect 20530 20380 20536 20392
rect 18656 20352 19840 20380
rect 20491 20352 20536 20380
rect 18656 20340 18662 20352
rect 19334 20272 19340 20324
rect 19392 20312 19398 20324
rect 19705 20315 19763 20321
rect 19705 20312 19717 20315
rect 19392 20284 19717 20312
rect 19392 20272 19398 20284
rect 19705 20281 19717 20284
rect 19751 20281 19763 20315
rect 19812 20312 19840 20352
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 26896 20312 26924 20556
rect 28721 20519 28779 20525
rect 28721 20485 28733 20519
rect 28767 20516 28779 20519
rect 28994 20516 29000 20528
rect 28767 20488 29000 20516
rect 28767 20485 28779 20488
rect 28721 20479 28779 20485
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 29730 20476 29736 20528
rect 29788 20476 29794 20528
rect 32953 20519 33011 20525
rect 32953 20485 32965 20519
rect 32999 20516 33011 20519
rect 33226 20516 33232 20528
rect 32999 20488 33232 20516
rect 32999 20485 33011 20488
rect 32953 20479 33011 20485
rect 33226 20476 33232 20488
rect 33284 20476 33290 20528
rect 43254 20476 43260 20528
rect 43312 20516 43318 20528
rect 44913 20519 44971 20525
rect 44913 20516 44925 20519
rect 43312 20488 44925 20516
rect 43312 20476 43318 20488
rect 44913 20485 44925 20488
rect 44959 20485 44971 20519
rect 44913 20479 44971 20485
rect 28442 20448 28448 20460
rect 28403 20420 28448 20448
rect 28442 20408 28448 20420
rect 28500 20408 28506 20460
rect 32122 20448 32128 20460
rect 32083 20420 32128 20448
rect 32122 20408 32128 20420
rect 32180 20408 32186 20460
rect 43070 20448 43076 20460
rect 43031 20420 43076 20448
rect 43070 20408 43076 20420
rect 43128 20408 43134 20460
rect 43438 20448 43444 20460
rect 43399 20420 43444 20448
rect 43438 20408 43444 20420
rect 43496 20408 43502 20460
rect 44358 20408 44364 20460
rect 44416 20448 44422 20460
rect 44545 20451 44603 20457
rect 44545 20448 44557 20451
rect 44416 20420 44557 20448
rect 44416 20408 44422 20420
rect 44545 20417 44557 20420
rect 44591 20417 44603 20451
rect 44726 20448 44732 20460
rect 44687 20420 44732 20448
rect 44545 20411 44603 20417
rect 44726 20408 44732 20420
rect 44784 20408 44790 20460
rect 45572 20457 45600 20556
rect 45649 20553 45661 20587
rect 45695 20584 45707 20587
rect 46474 20584 46480 20596
rect 45695 20556 46480 20584
rect 45695 20553 45707 20556
rect 45649 20547 45707 20553
rect 46474 20544 46480 20556
rect 46532 20544 46538 20596
rect 48038 20584 48044 20596
rect 47999 20556 48044 20584
rect 48038 20544 48044 20556
rect 48096 20544 48102 20596
rect 45557 20451 45615 20457
rect 45557 20417 45569 20451
rect 45603 20417 45615 20451
rect 45557 20411 45615 20417
rect 45830 20408 45836 20460
rect 45888 20448 45894 20460
rect 46201 20451 46259 20457
rect 46201 20448 46213 20451
rect 45888 20420 46213 20448
rect 45888 20408 45894 20420
rect 46201 20417 46213 20420
rect 46247 20417 46259 20451
rect 46201 20411 46259 20417
rect 47394 20408 47400 20460
rect 47452 20448 47458 20460
rect 47581 20451 47639 20457
rect 47581 20448 47593 20451
rect 47452 20420 47593 20448
rect 47452 20408 47458 20420
rect 47581 20417 47593 20420
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 29086 20340 29092 20392
rect 29144 20380 29150 20392
rect 30193 20383 30251 20389
rect 30193 20380 30205 20383
rect 29144 20352 30205 20380
rect 29144 20340 29150 20352
rect 30193 20349 30205 20352
rect 30239 20380 30251 20383
rect 32769 20383 32827 20389
rect 32769 20380 32781 20383
rect 30239 20352 32781 20380
rect 30239 20349 30251 20352
rect 30193 20343 30251 20349
rect 32769 20349 32781 20352
rect 32815 20349 32827 20383
rect 34422 20380 34428 20392
rect 34383 20352 34428 20380
rect 32769 20343 32827 20349
rect 34422 20340 34428 20352
rect 34480 20340 34486 20392
rect 43898 20340 43904 20392
rect 43956 20380 43962 20392
rect 43993 20383 44051 20389
rect 43993 20380 44005 20383
rect 43956 20352 44005 20380
rect 43956 20340 43962 20352
rect 43993 20349 44005 20352
rect 44039 20349 44051 20383
rect 43993 20343 44051 20349
rect 45738 20340 45744 20392
rect 45796 20380 45802 20392
rect 46477 20383 46535 20389
rect 46477 20380 46489 20383
rect 45796 20352 46489 20380
rect 45796 20340 45802 20352
rect 46477 20349 46489 20352
rect 46523 20349 46535 20383
rect 46477 20343 46535 20349
rect 19812 20284 26924 20312
rect 19705 20275 19763 20281
rect 17034 20204 17040 20256
rect 17092 20244 17098 20256
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 17092 20216 17417 20244
rect 17092 20204 17098 20216
rect 17405 20213 17417 20216
rect 17451 20213 17463 20247
rect 17405 20207 17463 20213
rect 19886 20204 19892 20256
rect 19944 20244 19950 20256
rect 20809 20247 20867 20253
rect 20809 20244 20821 20247
rect 19944 20216 20821 20244
rect 19944 20204 19950 20216
rect 20809 20213 20821 20216
rect 20855 20213 20867 20247
rect 21910 20244 21916 20256
rect 21871 20216 21916 20244
rect 20809 20207 20867 20213
rect 21910 20204 21916 20216
rect 21968 20204 21974 20256
rect 32214 20244 32220 20256
rect 32175 20216 32220 20244
rect 32214 20204 32220 20216
rect 32272 20204 32278 20256
rect 47670 20244 47676 20256
rect 47631 20216 47676 20244
rect 47670 20204 47676 20216
rect 47728 20204 47734 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 3418 20000 3424 20052
rect 3476 20040 3482 20052
rect 27246 20040 27252 20052
rect 3476 20012 27252 20040
rect 3476 20000 3482 20012
rect 27246 20000 27252 20012
rect 27304 20000 27310 20052
rect 28626 20000 28632 20052
rect 28684 20040 28690 20052
rect 28813 20043 28871 20049
rect 28813 20040 28825 20043
rect 28684 20012 28825 20040
rect 28684 20000 28690 20012
rect 28813 20009 28825 20012
rect 28859 20009 28871 20043
rect 28813 20003 28871 20009
rect 30745 20043 30803 20049
rect 30745 20009 30757 20043
rect 30791 20040 30803 20043
rect 31018 20040 31024 20052
rect 30791 20012 31024 20040
rect 30791 20009 30803 20012
rect 30745 20003 30803 20009
rect 31018 20000 31024 20012
rect 31076 20000 31082 20052
rect 42978 20040 42984 20052
rect 42939 20012 42984 20040
rect 42978 20000 42984 20012
rect 43036 20000 43042 20052
rect 43346 20000 43352 20052
rect 43404 20040 43410 20052
rect 43809 20043 43867 20049
rect 43809 20040 43821 20043
rect 43404 20012 43821 20040
rect 43404 20000 43410 20012
rect 43809 20009 43821 20012
rect 43855 20009 43867 20043
rect 43809 20003 43867 20009
rect 47854 20000 47860 20052
rect 47912 20040 47918 20052
rect 48041 20043 48099 20049
rect 48041 20040 48053 20043
rect 47912 20012 48053 20040
rect 47912 20000 47918 20012
rect 48041 20009 48053 20012
rect 48087 20009 48099 20043
rect 48041 20003 48099 20009
rect 10686 19972 10692 19984
rect 10647 19944 10692 19972
rect 10686 19932 10692 19944
rect 10744 19932 10750 19984
rect 12066 19972 12072 19984
rect 12027 19944 12072 19972
rect 12066 19932 12072 19944
rect 12124 19932 12130 19984
rect 15470 19972 15476 19984
rect 15431 19944 15476 19972
rect 15470 19932 15476 19944
rect 15528 19932 15534 19984
rect 23290 19932 23296 19984
rect 23348 19972 23354 19984
rect 23753 19975 23811 19981
rect 23753 19972 23765 19975
rect 23348 19944 23765 19972
rect 23348 19932 23354 19944
rect 23753 19941 23765 19944
rect 23799 19941 23811 19975
rect 23753 19935 23811 19941
rect 27338 19932 27344 19984
rect 27396 19972 27402 19984
rect 43533 19975 43591 19981
rect 27396 19944 41414 19972
rect 27396 19932 27402 19944
rect 16850 19904 16856 19916
rect 16811 19876 16856 19904
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 17034 19904 17040 19916
rect 16995 19876 17040 19904
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 19484 19876 19625 19904
rect 19484 19864 19490 19876
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 19886 19904 19892 19916
rect 19847 19876 19892 19904
rect 19613 19867 19671 19873
rect 19886 19864 19892 19876
rect 19944 19864 19950 19916
rect 19978 19864 19984 19916
rect 20036 19904 20042 19916
rect 20036 19876 26924 19904
rect 20036 19864 20042 19876
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19836 11299 19839
rect 11330 19836 11336 19848
rect 11287 19808 11336 19836
rect 11287 19805 11299 19808
rect 11241 19799 11299 19805
rect 10704 19768 10732 19799
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 11974 19836 11980 19848
rect 11935 19808 11980 19836
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19805 12863 19839
rect 14366 19836 14372 19848
rect 14327 19808 14372 19836
rect 12805 19799 12863 19805
rect 10870 19768 10876 19780
rect 10704 19740 10876 19768
rect 10870 19728 10876 19740
rect 10928 19768 10934 19780
rect 12820 19768 12848 19799
rect 14366 19796 14372 19808
rect 14424 19836 14430 19848
rect 15102 19836 15108 19848
rect 14424 19808 15108 19836
rect 14424 19796 14430 19808
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19836 15439 19839
rect 16758 19836 16764 19848
rect 15427 19808 16764 19836
rect 15427 19805 15439 19808
rect 15381 19799 15439 19805
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 22002 19836 22008 19848
rect 21963 19808 22008 19836
rect 22002 19796 22008 19808
rect 22060 19796 22066 19848
rect 23382 19796 23388 19848
rect 23440 19796 23446 19848
rect 26326 19796 26332 19848
rect 26384 19836 26390 19848
rect 26789 19839 26847 19845
rect 26789 19836 26801 19839
rect 26384 19808 26801 19836
rect 26384 19796 26390 19808
rect 26789 19805 26801 19808
rect 26835 19805 26847 19839
rect 26896 19836 26924 19876
rect 27246 19864 27252 19916
rect 27304 19904 27310 19916
rect 31757 19907 31815 19913
rect 31757 19904 31769 19907
rect 27304 19876 31769 19904
rect 27304 19864 27310 19876
rect 31757 19873 31769 19876
rect 31803 19873 31815 19907
rect 31757 19867 31815 19873
rect 27338 19836 27344 19848
rect 26896 19808 27344 19836
rect 26789 19799 26847 19805
rect 27338 19796 27344 19808
rect 27396 19796 27402 19848
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19805 28687 19839
rect 28629 19799 28687 19805
rect 13262 19768 13268 19780
rect 10928 19740 13268 19768
rect 10928 19728 10934 19740
rect 11440 19709 11468 19740
rect 13262 19728 13268 19740
rect 13320 19728 13326 19780
rect 18693 19771 18751 19777
rect 18693 19737 18705 19771
rect 18739 19768 18751 19771
rect 19978 19768 19984 19780
rect 18739 19740 19984 19768
rect 18739 19737 18751 19740
rect 18693 19731 18751 19737
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 21910 19768 21916 19780
rect 21114 19740 21916 19768
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 22278 19768 22284 19780
rect 22239 19740 22284 19768
rect 22278 19728 22284 19740
rect 22336 19728 22342 19780
rect 24578 19728 24584 19780
rect 24636 19768 24642 19780
rect 28644 19768 28672 19799
rect 30466 19796 30472 19848
rect 30524 19836 30530 19848
rect 30653 19839 30711 19845
rect 30653 19836 30665 19839
rect 30524 19808 30665 19836
rect 30524 19796 30530 19808
rect 30653 19805 30665 19808
rect 30699 19805 30711 19839
rect 31294 19836 31300 19848
rect 31255 19808 31300 19836
rect 30653 19799 30711 19805
rect 31294 19796 31300 19808
rect 31352 19796 31358 19848
rect 24636 19740 28672 19768
rect 31481 19771 31539 19777
rect 24636 19728 24642 19740
rect 31481 19737 31493 19771
rect 31527 19768 31539 19771
rect 41386 19768 41414 19944
rect 43533 19941 43545 19975
rect 43579 19972 43591 19975
rect 44174 19972 44180 19984
rect 43579 19944 44180 19972
rect 43579 19941 43591 19944
rect 43533 19935 43591 19941
rect 44174 19932 44180 19944
rect 44232 19932 44238 19984
rect 43898 19864 43904 19916
rect 43956 19904 43962 19916
rect 45557 19907 45615 19913
rect 45557 19904 45569 19907
rect 43956 19876 45569 19904
rect 43956 19864 43962 19876
rect 45557 19873 45569 19876
rect 45603 19873 45615 19907
rect 45738 19904 45744 19916
rect 45699 19876 45744 19904
rect 45557 19867 45615 19873
rect 45738 19864 45744 19876
rect 45796 19864 45802 19916
rect 46934 19904 46940 19916
rect 46895 19876 46940 19904
rect 46934 19864 46940 19876
rect 46992 19904 46998 19916
rect 47118 19904 47124 19916
rect 46992 19876 47124 19904
rect 46992 19864 46998 19876
rect 47118 19864 47124 19876
rect 47176 19864 47182 19916
rect 42886 19836 42892 19848
rect 42847 19808 42892 19836
rect 42886 19796 42892 19808
rect 42944 19796 42950 19848
rect 43070 19836 43076 19848
rect 43031 19808 43076 19836
rect 43070 19796 43076 19808
rect 43128 19836 43134 19848
rect 43530 19836 43536 19848
rect 43128 19808 43536 19836
rect 43128 19796 43134 19808
rect 43530 19796 43536 19808
rect 43588 19796 43594 19848
rect 43806 19836 43812 19848
rect 43767 19808 43812 19836
rect 43806 19796 43812 19808
rect 43864 19796 43870 19848
rect 43990 19836 43996 19848
rect 43951 19808 43996 19836
rect 43990 19796 43996 19808
rect 44048 19796 44054 19848
rect 46566 19768 46572 19780
rect 31527 19740 31754 19768
rect 41386 19740 46572 19768
rect 31527 19737 31539 19740
rect 31481 19731 31539 19737
rect 11425 19703 11483 19709
rect 11425 19669 11437 19703
rect 11471 19669 11483 19703
rect 11425 19663 11483 19669
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 12989 19703 13047 19709
rect 12989 19700 13001 19703
rect 12952 19672 13001 19700
rect 12952 19660 12958 19672
rect 12989 19669 13001 19672
rect 13035 19669 13047 19703
rect 14458 19700 14464 19712
rect 14419 19672 14464 19700
rect 12989 19663 13047 19669
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 21361 19703 21419 19709
rect 21361 19700 21373 19703
rect 20680 19672 21373 19700
rect 20680 19660 20686 19672
rect 21361 19669 21373 19672
rect 21407 19669 21419 19703
rect 21361 19663 21419 19669
rect 26605 19703 26663 19709
rect 26605 19669 26617 19703
rect 26651 19700 26663 19703
rect 27062 19700 27068 19712
rect 26651 19672 27068 19700
rect 26651 19669 26663 19672
rect 26605 19663 26663 19669
rect 27062 19660 27068 19672
rect 27120 19660 27126 19712
rect 31726 19700 31754 19740
rect 46566 19728 46572 19740
rect 46624 19728 46630 19780
rect 32214 19700 32220 19712
rect 31726 19672 32220 19700
rect 32214 19660 32220 19672
rect 32272 19660 32278 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 14090 19456 14096 19508
rect 14148 19496 14154 19508
rect 14645 19499 14703 19505
rect 14645 19496 14657 19499
rect 14148 19468 14657 19496
rect 14148 19456 14154 19468
rect 14645 19465 14657 19468
rect 14691 19496 14703 19499
rect 14691 19468 15148 19496
rect 14691 19465 14703 19468
rect 14645 19459 14703 19465
rect 14458 19428 14464 19440
rect 14398 19400 14464 19428
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 15120 19437 15148 19468
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18417 19499 18475 19505
rect 18417 19496 18429 19499
rect 18012 19468 18429 19496
rect 18012 19456 18018 19468
rect 18417 19465 18429 19468
rect 18463 19465 18475 19499
rect 18417 19459 18475 19465
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 19024 19468 19073 19496
rect 19024 19456 19030 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 22278 19456 22284 19508
rect 22336 19496 22342 19508
rect 22925 19499 22983 19505
rect 22925 19496 22937 19499
rect 22336 19468 22937 19496
rect 22336 19456 22342 19468
rect 22925 19465 22937 19468
rect 22971 19465 22983 19499
rect 26326 19496 26332 19508
rect 26287 19468 26332 19496
rect 22925 19459 22983 19465
rect 26326 19456 26332 19468
rect 26384 19456 26390 19508
rect 31113 19499 31171 19505
rect 31113 19465 31125 19499
rect 31159 19496 31171 19499
rect 31294 19496 31300 19508
rect 31159 19468 31300 19496
rect 31159 19465 31171 19468
rect 31113 19459 31171 19465
rect 31294 19456 31300 19468
rect 31352 19496 31358 19508
rect 31938 19496 31944 19508
rect 31352 19468 31944 19496
rect 31352 19456 31358 19468
rect 31938 19456 31944 19468
rect 31996 19456 32002 19508
rect 43438 19496 43444 19508
rect 43399 19468 43444 19496
rect 43438 19456 43444 19468
rect 43496 19456 43502 19508
rect 44269 19499 44327 19505
rect 44269 19465 44281 19499
rect 44315 19496 44327 19499
rect 44542 19496 44548 19508
rect 44315 19468 44548 19496
rect 44315 19465 44327 19468
rect 44269 19459 44327 19465
rect 44542 19456 44548 19468
rect 44600 19456 44606 19508
rect 46014 19456 46020 19508
rect 46072 19496 46078 19508
rect 46753 19499 46811 19505
rect 46753 19496 46765 19499
rect 46072 19468 46765 19496
rect 46072 19456 46078 19468
rect 46753 19465 46765 19468
rect 46799 19496 46811 19499
rect 47302 19496 47308 19508
rect 46799 19468 47308 19496
rect 46799 19465 46811 19468
rect 46753 19459 46811 19465
rect 47302 19456 47308 19468
rect 47360 19456 47366 19508
rect 15105 19431 15163 19437
rect 15105 19397 15117 19431
rect 15151 19397 15163 19431
rect 15105 19391 15163 19397
rect 15289 19431 15347 19437
rect 15289 19397 15301 19431
rect 15335 19428 15347 19431
rect 16850 19428 16856 19440
rect 15335 19400 16856 19428
rect 15335 19397 15347 19400
rect 15289 19391 15347 19397
rect 16850 19388 16856 19400
rect 16908 19388 16914 19440
rect 19334 19428 19340 19440
rect 18340 19400 19340 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 10870 19360 10876 19372
rect 10831 19332 10876 19360
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 11974 19360 11980 19372
rect 11563 19332 11980 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12894 19360 12900 19372
rect 12855 19332 12900 19360
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 14734 19320 14740 19372
rect 14792 19360 14798 19372
rect 18340 19369 18368 19400
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 22002 19388 22008 19440
rect 22060 19428 22066 19440
rect 34054 19428 34060 19440
rect 22060 19400 34060 19428
rect 22060 19388 22066 19400
rect 34054 19388 34060 19400
rect 34112 19388 34118 19440
rect 46382 19388 46388 19440
rect 46440 19428 46446 19440
rect 46661 19431 46719 19437
rect 46661 19428 46673 19431
rect 46440 19400 46673 19428
rect 46440 19388 46446 19400
rect 46661 19397 46673 19400
rect 46707 19397 46719 19431
rect 46661 19391 46719 19397
rect 46937 19431 46995 19437
rect 46937 19397 46949 19431
rect 46983 19428 46995 19431
rect 47394 19428 47400 19440
rect 46983 19400 47400 19428
rect 46983 19397 46995 19400
rect 46937 19391 46995 19397
rect 47394 19388 47400 19400
rect 47452 19388 47458 19440
rect 15381 19363 15439 19369
rect 15381 19360 15393 19363
rect 14792 19332 15393 19360
rect 14792 19320 14798 19332
rect 15381 19329 15393 19332
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19329 18383 19363
rect 18325 19323 18383 19329
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19360 19027 19363
rect 19150 19360 19156 19372
rect 19015 19332 19156 19360
rect 19015 19329 19027 19332
rect 18969 19323 19027 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 13170 19292 13176 19304
rect 13131 19264 13176 19292
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 14366 19252 14372 19304
rect 14424 19292 14430 19304
rect 15488 19292 15516 19323
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 22833 19363 22891 19369
rect 22833 19329 22845 19363
rect 22879 19360 22891 19363
rect 23290 19360 23296 19372
rect 22879 19332 23296 19360
rect 22879 19329 22891 19332
rect 22833 19323 22891 19329
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 26142 19360 26148 19372
rect 26103 19332 26148 19360
rect 26142 19320 26148 19332
rect 26200 19320 26206 19372
rect 26510 19320 26516 19372
rect 26568 19360 26574 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26568 19332 26985 19360
rect 26568 19320 26574 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 28169 19363 28227 19369
rect 28169 19329 28181 19363
rect 28215 19329 28227 19363
rect 28169 19323 28227 19329
rect 15654 19292 15660 19304
rect 14424 19264 15516 19292
rect 15615 19264 15660 19292
rect 14424 19252 14430 19264
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 19058 19252 19064 19304
rect 19116 19292 19122 19304
rect 19518 19292 19524 19304
rect 19116 19264 19524 19292
rect 19116 19252 19122 19264
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 25590 19252 25596 19304
rect 25648 19292 25654 19304
rect 25961 19295 26019 19301
rect 25961 19292 25973 19295
rect 25648 19264 25973 19292
rect 25648 19252 25654 19264
rect 25961 19261 25973 19264
rect 26007 19261 26019 19295
rect 28184 19292 28212 19323
rect 28258 19320 28264 19372
rect 28316 19360 28322 19372
rect 28626 19360 28632 19372
rect 28316 19332 28361 19360
rect 28460 19332 28632 19360
rect 28316 19320 28322 19332
rect 28460 19292 28488 19332
rect 28626 19320 28632 19332
rect 28684 19360 28690 19372
rect 28813 19363 28871 19369
rect 28813 19360 28825 19363
rect 28684 19332 28825 19360
rect 28684 19320 28690 19332
rect 28813 19329 28825 19332
rect 28859 19329 28871 19363
rect 28813 19323 28871 19329
rect 31202 19320 31208 19372
rect 31260 19360 31266 19372
rect 31297 19363 31355 19369
rect 31297 19360 31309 19363
rect 31260 19332 31309 19360
rect 31260 19320 31266 19332
rect 31297 19329 31309 19332
rect 31343 19329 31355 19363
rect 32122 19360 32128 19372
rect 32083 19332 32128 19360
rect 31297 19323 31355 19329
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 43346 19360 43352 19372
rect 43307 19332 43352 19360
rect 43346 19320 43352 19332
rect 43404 19320 43410 19372
rect 43533 19363 43591 19369
rect 43533 19329 43545 19363
rect 43579 19360 43591 19363
rect 44082 19360 44088 19372
rect 43579 19332 44088 19360
rect 43579 19329 43591 19332
rect 43533 19323 43591 19329
rect 44082 19320 44088 19332
rect 44140 19320 44146 19372
rect 44266 19360 44272 19372
rect 44227 19332 44272 19360
rect 44266 19320 44272 19332
rect 44324 19320 44330 19372
rect 46569 19363 46627 19369
rect 46569 19329 46581 19363
rect 46615 19360 46627 19363
rect 46750 19360 46756 19372
rect 46615 19332 46756 19360
rect 46615 19329 46627 19332
rect 46569 19323 46627 19329
rect 46750 19320 46756 19332
rect 46808 19320 46814 19372
rect 28184 19264 28488 19292
rect 25961 19255 26019 19261
rect 35342 19184 35348 19236
rect 35400 19224 35406 19236
rect 46385 19227 46443 19233
rect 46385 19224 46397 19227
rect 35400 19196 46397 19224
rect 35400 19184 35406 19196
rect 46385 19193 46397 19196
rect 46431 19224 46443 19227
rect 47026 19224 47032 19236
rect 46431 19196 47032 19224
rect 46431 19193 46443 19196
rect 46385 19187 46443 19193
rect 47026 19184 47032 19196
rect 47084 19184 47090 19236
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 10689 19159 10747 19165
rect 10689 19156 10701 19159
rect 10468 19128 10701 19156
rect 10468 19116 10474 19128
rect 10689 19125 10701 19128
rect 10735 19125 10747 19159
rect 10689 19119 10747 19125
rect 11609 19159 11667 19165
rect 11609 19125 11621 19159
rect 11655 19156 11667 19159
rect 11698 19156 11704 19168
rect 11655 19128 11704 19156
rect 11655 19125 11667 19128
rect 11609 19119 11667 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 26786 19116 26792 19168
rect 26844 19156 26850 19168
rect 26973 19159 27031 19165
rect 26973 19156 26985 19159
rect 26844 19128 26985 19156
rect 26844 19116 26850 19128
rect 26973 19125 26985 19128
rect 27019 19125 27031 19159
rect 28902 19156 28908 19168
rect 28863 19128 28908 19156
rect 26973 19119 27031 19125
rect 28902 19116 28908 19128
rect 28960 19116 28966 19168
rect 32214 19156 32220 19168
rect 32175 19128 32220 19156
rect 32214 19116 32220 19128
rect 32272 19116 32278 19168
rect 47762 19156 47768 19168
rect 47723 19128 47768 19156
rect 47762 19116 47768 19128
rect 47820 19116 47826 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 4982 18912 4988 18964
rect 5040 18952 5046 18964
rect 28994 18952 29000 18964
rect 5040 18924 29000 18952
rect 5040 18912 5046 18924
rect 28994 18912 29000 18924
rect 29052 18952 29058 18964
rect 33781 18955 33839 18961
rect 29052 18924 30144 18952
rect 29052 18912 29058 18924
rect 12897 18887 12955 18893
rect 12897 18853 12909 18887
rect 12943 18884 12955 18887
rect 13170 18884 13176 18896
rect 12943 18856 13176 18884
rect 12943 18853 12955 18856
rect 12897 18847 12955 18853
rect 13170 18844 13176 18856
rect 13228 18844 13234 18896
rect 13814 18844 13820 18896
rect 13872 18884 13878 18896
rect 22370 18884 22376 18896
rect 13872 18856 22376 18884
rect 13872 18844 13878 18856
rect 22370 18844 22376 18856
rect 22428 18844 22434 18896
rect 10410 18816 10416 18828
rect 10371 18788 10416 18816
rect 10410 18776 10416 18788
rect 10468 18776 10474 18828
rect 15013 18819 15071 18825
rect 15013 18816 15025 18819
rect 13372 18788 15025 18816
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 2188 18720 6914 18748
rect 2188 18708 2194 18720
rect 6886 18612 6914 18720
rect 12342 18708 12348 18760
rect 12400 18748 12406 18760
rect 13372 18757 13400 18788
rect 15013 18785 15025 18788
rect 15059 18785 15071 18819
rect 23106 18816 23112 18828
rect 15013 18779 15071 18785
rect 21744 18788 23112 18816
rect 13081 18751 13139 18757
rect 13081 18748 13093 18751
rect 12400 18720 13093 18748
rect 12400 18708 12406 18720
rect 13081 18717 13093 18720
rect 13127 18717 13139 18751
rect 13081 18711 13139 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 14090 18748 14096 18760
rect 13587 18720 14096 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 14734 18748 14740 18760
rect 14691 18720 14740 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 19518 18748 19524 18760
rect 19475 18720 19524 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 19518 18708 19524 18720
rect 19576 18748 19582 18760
rect 20806 18748 20812 18760
rect 19576 18720 20812 18748
rect 19576 18708 19582 18720
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 10689 18683 10747 18689
rect 10689 18649 10701 18683
rect 10735 18680 10747 18683
rect 10962 18680 10968 18692
rect 10735 18652 10968 18680
rect 10735 18649 10747 18652
rect 10689 18643 10747 18649
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 11698 18640 11704 18692
rect 11756 18640 11762 18692
rect 14458 18680 14464 18692
rect 11992 18652 12434 18680
rect 14419 18652 14464 18680
rect 11992 18612 12020 18652
rect 12158 18612 12164 18624
rect 6886 18584 12020 18612
rect 12119 18584 12164 18612
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 12406 18612 12434 18652
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 21744 18680 21772 18788
rect 23106 18776 23112 18788
rect 23164 18816 23170 18828
rect 23164 18788 23244 18816
rect 23164 18776 23170 18788
rect 21818 18708 21824 18760
rect 21876 18748 21882 18760
rect 23216 18757 23244 18788
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24486 18816 24492 18828
rect 23716 18788 24492 18816
rect 23716 18776 23722 18788
rect 24486 18776 24492 18788
rect 24544 18816 24550 18828
rect 24544 18788 24716 18816
rect 24544 18776 24550 18788
rect 23201 18751 23259 18757
rect 21876 18720 23152 18748
rect 21876 18708 21882 18720
rect 22005 18683 22063 18689
rect 22005 18680 22017 18683
rect 19392 18652 19656 18680
rect 21744 18652 22017 18680
rect 19392 18640 19398 18652
rect 13354 18612 13360 18624
rect 12406 18584 13360 18612
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 14737 18615 14795 18621
rect 14737 18612 14749 18615
rect 14424 18584 14749 18612
rect 14424 18572 14430 18584
rect 14737 18581 14749 18584
rect 14783 18581 14795 18615
rect 14737 18575 14795 18581
rect 14829 18615 14887 18621
rect 14829 18581 14841 18615
rect 14875 18612 14887 18615
rect 14918 18612 14924 18624
rect 14875 18584 14924 18612
rect 14875 18581 14887 18584
rect 14829 18575 14887 18581
rect 14918 18572 14924 18584
rect 14976 18572 14982 18624
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 16758 18612 16764 18624
rect 15068 18584 16764 18612
rect 15068 18572 15074 18584
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 19521 18615 19579 18621
rect 19521 18612 19533 18615
rect 19484 18584 19533 18612
rect 19484 18572 19490 18584
rect 19521 18581 19533 18584
rect 19567 18581 19579 18615
rect 19628 18612 19656 18652
rect 22005 18649 22017 18652
rect 22051 18649 22063 18683
rect 23124 18680 23152 18720
rect 23201 18717 23213 18751
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 24397 18751 24455 18757
rect 24397 18717 24409 18751
rect 24443 18748 24455 18751
rect 24578 18748 24584 18760
rect 24443 18720 24584 18748
rect 24443 18717 24455 18720
rect 24397 18711 24455 18717
rect 24578 18708 24584 18720
rect 24636 18708 24642 18760
rect 24688 18748 24716 18788
rect 25590 18776 25596 18828
rect 25648 18816 25654 18828
rect 25869 18819 25927 18825
rect 25869 18816 25881 18819
rect 25648 18788 25881 18816
rect 25648 18776 25654 18788
rect 25869 18785 25881 18788
rect 25915 18785 25927 18819
rect 26786 18816 26792 18828
rect 26747 18788 26792 18816
rect 25869 18779 25927 18785
rect 26786 18776 26792 18788
rect 26844 18776 26850 18828
rect 27062 18816 27068 18828
rect 27023 18788 27068 18816
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 30116 18760 30144 18924
rect 33781 18921 33793 18955
rect 33827 18952 33839 18955
rect 35342 18952 35348 18964
rect 33827 18924 35348 18952
rect 33827 18921 33839 18924
rect 33781 18915 33839 18921
rect 35342 18912 35348 18924
rect 35400 18912 35406 18964
rect 31389 18819 31447 18825
rect 31389 18785 31401 18819
rect 31435 18816 31447 18819
rect 32214 18816 32220 18828
rect 31435 18788 32220 18816
rect 31435 18785 31447 18788
rect 31389 18779 31447 18785
rect 32214 18776 32220 18788
rect 32272 18776 32278 18828
rect 32306 18776 32312 18828
rect 32364 18816 32370 18828
rect 46293 18819 46351 18825
rect 32364 18788 32409 18816
rect 32364 18776 32370 18788
rect 46293 18785 46305 18819
rect 46339 18816 46351 18819
rect 47762 18816 47768 18828
rect 46339 18788 47768 18816
rect 46339 18785 46351 18788
rect 46293 18779 46351 18785
rect 47762 18776 47768 18788
rect 47820 18776 47826 18828
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 25958 18748 25964 18760
rect 24688 18720 25964 18748
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18748 29975 18751
rect 30006 18748 30012 18760
rect 29963 18720 30012 18748
rect 29963 18717 29975 18720
rect 29917 18711 29975 18717
rect 30006 18708 30012 18720
rect 30064 18708 30070 18760
rect 30098 18708 30104 18760
rect 30156 18748 30162 18760
rect 30156 18720 30249 18748
rect 30156 18708 30162 18720
rect 31110 18708 31116 18760
rect 31168 18748 31174 18760
rect 31205 18751 31263 18757
rect 31205 18748 31217 18751
rect 31168 18720 31217 18748
rect 31168 18708 31174 18720
rect 31205 18717 31217 18720
rect 31251 18717 31263 18751
rect 33502 18748 33508 18760
rect 33415 18720 33508 18748
rect 31205 18711 31263 18717
rect 33502 18708 33508 18720
rect 33560 18748 33566 18760
rect 35526 18748 35532 18760
rect 33560 18720 35532 18748
rect 33560 18708 33566 18720
rect 35526 18708 35532 18720
rect 35584 18708 35590 18760
rect 45830 18748 45836 18760
rect 45791 18720 45836 18748
rect 45830 18708 45836 18720
rect 45888 18708 45894 18760
rect 28902 18680 28908 18692
rect 23124 18652 27476 18680
rect 28290 18652 28908 18680
rect 22005 18643 22063 18649
rect 19978 18612 19984 18624
rect 19628 18584 19984 18612
rect 19521 18575 19579 18581
rect 19978 18572 19984 18584
rect 20036 18612 20042 18624
rect 22097 18615 22155 18621
rect 22097 18612 22109 18615
rect 20036 18584 22109 18612
rect 20036 18572 20042 18584
rect 22097 18581 22109 18584
rect 22143 18581 22155 18615
rect 22097 18575 22155 18581
rect 23290 18572 23296 18624
rect 23348 18612 23354 18624
rect 23385 18615 23443 18621
rect 23385 18612 23397 18615
rect 23348 18584 23397 18612
rect 23348 18572 23354 18584
rect 23385 18581 23397 18584
rect 23431 18581 23443 18615
rect 23385 18575 23443 18581
rect 24581 18615 24639 18621
rect 24581 18581 24593 18615
rect 24627 18612 24639 18615
rect 24762 18612 24768 18624
rect 24627 18584 24768 18612
rect 24627 18581 24639 18584
rect 24581 18575 24639 18581
rect 24762 18572 24768 18584
rect 24820 18572 24826 18624
rect 26329 18615 26387 18621
rect 26329 18581 26341 18615
rect 26375 18612 26387 18615
rect 27246 18612 27252 18624
rect 26375 18584 27252 18612
rect 26375 18581 26387 18584
rect 26329 18575 26387 18581
rect 27246 18572 27252 18584
rect 27304 18572 27310 18624
rect 27448 18612 27476 18652
rect 28902 18640 28908 18652
rect 28960 18640 28966 18692
rect 34606 18680 34612 18692
rect 29012 18652 34612 18680
rect 28537 18615 28595 18621
rect 28537 18612 28549 18615
rect 27448 18584 28549 18612
rect 28537 18581 28549 18584
rect 28583 18612 28595 18615
rect 29012 18612 29040 18652
rect 34606 18640 34612 18652
rect 34664 18640 34670 18692
rect 46477 18683 46535 18689
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 47670 18680 47676 18692
rect 46523 18652 47676 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 47670 18640 47676 18652
rect 47728 18640 47734 18692
rect 28583 18584 29040 18612
rect 30101 18615 30159 18621
rect 28583 18581 28595 18584
rect 28537 18575 28595 18581
rect 30101 18581 30113 18615
rect 30147 18612 30159 18615
rect 30190 18612 30196 18624
rect 30147 18584 30196 18612
rect 30147 18581 30159 18584
rect 30101 18575 30159 18581
rect 30190 18572 30196 18584
rect 30248 18572 30254 18624
rect 33965 18615 34023 18621
rect 33965 18581 33977 18615
rect 34011 18612 34023 18615
rect 34790 18612 34796 18624
rect 34011 18584 34796 18612
rect 34011 18581 34023 18584
rect 33965 18575 34023 18581
rect 34790 18572 34796 18584
rect 34848 18572 34854 18624
rect 45646 18612 45652 18624
rect 45607 18584 45652 18612
rect 45646 18572 45652 18584
rect 45704 18572 45710 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 47670 18408 47676 18420
rect 3476 18380 31754 18408
rect 47631 18380 47676 18408
rect 3476 18368 3482 18380
rect 12342 18340 12348 18352
rect 10520 18312 12348 18340
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 10520 18213 10548 18312
rect 12342 18300 12348 18312
rect 12400 18300 12406 18352
rect 14458 18300 14464 18352
rect 14516 18340 14522 18352
rect 16850 18340 16856 18352
rect 14516 18312 16856 18340
rect 14516 18300 14522 18312
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 11514 18272 11520 18284
rect 10643 18244 11520 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 11514 18232 11520 18244
rect 11572 18272 11578 18284
rect 12158 18272 12164 18284
rect 11572 18244 12164 18272
rect 11572 18232 11578 18244
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 13262 18272 13268 18284
rect 13223 18244 13268 18272
rect 13262 18232 13268 18244
rect 13320 18232 13326 18284
rect 14752 18281 14780 18312
rect 16850 18300 16856 18312
rect 16908 18300 16914 18352
rect 19426 18300 19432 18352
rect 19484 18340 19490 18352
rect 19613 18343 19671 18349
rect 19613 18340 19625 18343
rect 19484 18312 19625 18340
rect 19484 18300 19490 18312
rect 19613 18309 19625 18312
rect 19659 18309 19671 18343
rect 19613 18303 19671 18309
rect 23934 18300 23940 18352
rect 23992 18340 23998 18352
rect 25498 18340 25504 18352
rect 23992 18312 25504 18340
rect 23992 18300 23998 18312
rect 25498 18300 25504 18312
rect 25556 18340 25562 18352
rect 25593 18343 25651 18349
rect 25593 18340 25605 18343
rect 25556 18312 25605 18340
rect 25556 18300 25562 18312
rect 25593 18309 25605 18312
rect 25639 18340 25651 18343
rect 25961 18343 26019 18349
rect 25639 18312 25912 18340
rect 25639 18309 25651 18312
rect 25593 18303 25651 18309
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18241 13967 18275
rect 13909 18235 13967 18241
rect 14093 18275 14151 18281
rect 14093 18241 14105 18275
rect 14139 18272 14151 18275
rect 14737 18275 14795 18281
rect 14139 18244 14688 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 10505 18207 10563 18213
rect 10505 18173 10517 18207
rect 10551 18173 10563 18207
rect 10962 18204 10968 18216
rect 10923 18176 10968 18204
rect 10505 18167 10563 18173
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 13814 18204 13820 18216
rect 12406 18176 13820 18204
rect 1581 18139 1639 18145
rect 1581 18105 1593 18139
rect 1627 18136 1639 18139
rect 12406 18136 12434 18176
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 13924 18204 13952 18235
rect 14660 18216 14688 18244
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 15102 18232 15108 18284
rect 15160 18272 15166 18284
rect 15654 18272 15660 18284
rect 15160 18244 15660 18272
rect 15160 18232 15166 18244
rect 15654 18232 15660 18244
rect 15712 18272 15718 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15712 18244 15945 18272
rect 15712 18232 15718 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 16758 18272 16764 18284
rect 16719 18244 16764 18272
rect 15933 18235 15991 18241
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 16945 18275 17003 18281
rect 16945 18241 16957 18275
rect 16991 18272 17003 18275
rect 17034 18272 17040 18284
rect 16991 18244 17040 18272
rect 16991 18241 17003 18244
rect 16945 18235 17003 18241
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18272 18843 18275
rect 19334 18272 19340 18284
rect 18831 18244 19340 18272
rect 18831 18241 18843 18244
rect 18785 18235 18843 18241
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 21818 18272 21824 18284
rect 21779 18244 21824 18272
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 23842 18272 23848 18284
rect 23339 18244 23848 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 24210 18232 24216 18284
rect 24268 18272 24274 18284
rect 24762 18272 24768 18284
rect 24268 18244 24313 18272
rect 24723 18244 24768 18272
rect 24268 18232 24274 18244
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 25682 18232 25688 18284
rect 25740 18272 25746 18284
rect 25777 18275 25835 18281
rect 25777 18272 25789 18275
rect 25740 18244 25789 18272
rect 25740 18232 25746 18244
rect 25777 18241 25789 18244
rect 25823 18241 25835 18275
rect 25884 18272 25912 18312
rect 25961 18309 25973 18343
rect 26007 18340 26019 18343
rect 26142 18340 26148 18352
rect 26007 18312 26148 18340
rect 26007 18309 26019 18312
rect 25961 18303 26019 18309
rect 26142 18300 26148 18312
rect 26200 18300 26206 18352
rect 27246 18340 27252 18352
rect 27207 18312 27252 18340
rect 27246 18300 27252 18312
rect 27304 18300 27310 18352
rect 28258 18300 28264 18352
rect 28316 18300 28322 18352
rect 30006 18340 30012 18352
rect 29967 18312 30012 18340
rect 30006 18300 30012 18312
rect 30064 18300 30070 18352
rect 30098 18300 30104 18352
rect 30156 18340 30162 18352
rect 30193 18343 30251 18349
rect 30193 18340 30205 18343
rect 30156 18312 30205 18340
rect 30156 18300 30162 18312
rect 30193 18309 30205 18312
rect 30239 18309 30251 18343
rect 31202 18340 31208 18352
rect 31163 18312 31208 18340
rect 30193 18303 30251 18309
rect 31202 18300 31208 18312
rect 31260 18300 31266 18352
rect 31726 18340 31754 18380
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 32306 18340 32312 18352
rect 31726 18312 32312 18340
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 32493 18343 32551 18349
rect 32493 18309 32505 18343
rect 32539 18340 32551 18343
rect 33502 18340 33508 18352
rect 32539 18312 33508 18340
rect 32539 18309 32551 18312
rect 32493 18303 32551 18309
rect 33502 18300 33508 18312
rect 33560 18300 33566 18352
rect 43898 18340 43904 18352
rect 43364 18312 43904 18340
rect 26418 18272 26424 18284
rect 25884 18244 26424 18272
rect 25777 18235 25835 18241
rect 26418 18232 26424 18244
rect 26476 18232 26482 18284
rect 30377 18275 30435 18281
rect 30377 18241 30389 18275
rect 30423 18272 30435 18275
rect 31021 18275 31079 18281
rect 31021 18272 31033 18275
rect 30423 18244 31033 18272
rect 30423 18241 30435 18244
rect 30377 18235 30435 18241
rect 31021 18241 31033 18244
rect 31067 18241 31079 18275
rect 34790 18272 34796 18284
rect 34751 18244 34796 18272
rect 31021 18235 31079 18241
rect 34790 18232 34796 18244
rect 34848 18232 34854 18284
rect 43364 18281 43392 18312
rect 43898 18300 43904 18312
rect 43956 18300 43962 18352
rect 43349 18275 43407 18281
rect 43349 18241 43361 18275
rect 43395 18241 43407 18275
rect 46014 18272 46020 18284
rect 45975 18244 46020 18272
rect 43349 18235 43407 18241
rect 46014 18232 46020 18244
rect 46072 18232 46078 18284
rect 46382 18272 46388 18284
rect 46343 18244 46388 18272
rect 46382 18232 46388 18244
rect 46440 18232 46446 18284
rect 46750 18272 46756 18284
rect 46711 18244 46756 18272
rect 46750 18232 46756 18244
rect 46808 18232 46814 18284
rect 47026 18272 47032 18284
rect 46939 18244 47032 18272
rect 47026 18232 47032 18244
rect 47084 18232 47090 18284
rect 47578 18272 47584 18284
rect 47539 18244 47584 18272
rect 47578 18232 47584 18244
rect 47636 18232 47642 18284
rect 14550 18204 14556 18216
rect 13924 18176 14556 18204
rect 14550 18164 14556 18176
rect 14608 18164 14614 18216
rect 14642 18164 14648 18216
rect 14700 18204 14706 18216
rect 14700 18176 14793 18204
rect 14700 18164 14706 18176
rect 14918 18164 14924 18216
rect 14976 18204 14982 18216
rect 16776 18204 16804 18232
rect 19429 18207 19487 18213
rect 14976 18176 15608 18204
rect 16776 18176 19380 18204
rect 14976 18164 14982 18176
rect 1627 18108 12434 18136
rect 13357 18139 13415 18145
rect 1627 18105 1639 18108
rect 1581 18099 1639 18105
rect 13357 18105 13369 18139
rect 13403 18136 13415 18139
rect 15010 18136 15016 18148
rect 13403 18108 15016 18136
rect 13403 18105 13415 18108
rect 13357 18099 13415 18105
rect 15010 18096 15016 18108
rect 15068 18096 15074 18148
rect 15580 18136 15608 18176
rect 17129 18139 17187 18145
rect 17129 18136 17141 18139
rect 15580 18108 17141 18136
rect 17129 18105 17141 18108
rect 17175 18105 17187 18139
rect 17129 18099 17187 18105
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 13909 18071 13967 18077
rect 13909 18068 13921 18071
rect 13872 18040 13921 18068
rect 13872 18028 13878 18040
rect 13909 18037 13921 18040
rect 13955 18037 13967 18071
rect 13909 18031 13967 18037
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 15470 18068 15476 18080
rect 15151 18040 15476 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 16574 18068 16580 18080
rect 16071 18040 16580 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 18785 18071 18843 18077
rect 18785 18037 18797 18071
rect 18831 18068 18843 18071
rect 19242 18068 19248 18080
rect 18831 18040 19248 18068
rect 18831 18037 18843 18040
rect 18785 18031 18843 18037
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19352 18068 19380 18176
rect 19429 18173 19441 18207
rect 19475 18204 19487 18207
rect 20622 18204 20628 18216
rect 19475 18176 20628 18204
rect 19475 18173 19487 18176
rect 19429 18167 19487 18173
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 21266 18204 21272 18216
rect 21227 18176 21272 18204
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 23382 18204 23388 18216
rect 22152 18176 23388 18204
rect 22152 18164 22158 18176
rect 23382 18164 23388 18176
rect 23440 18204 23446 18216
rect 23934 18204 23940 18216
rect 23440 18176 23796 18204
rect 23895 18176 23940 18204
rect 23440 18164 23446 18176
rect 23768 18136 23796 18176
rect 23934 18164 23940 18176
rect 23992 18164 23998 18216
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18173 24087 18207
rect 24029 18167 24087 18173
rect 24121 18207 24179 18213
rect 24121 18173 24133 18207
rect 24167 18204 24179 18207
rect 24486 18204 24492 18216
rect 24167 18176 24492 18204
rect 24167 18173 24179 18176
rect 24121 18167 24179 18173
rect 24044 18136 24072 18167
rect 24486 18164 24492 18176
rect 24544 18164 24550 18216
rect 26970 18204 26976 18216
rect 26931 18176 26976 18204
rect 26970 18164 26976 18176
rect 27028 18164 27034 18216
rect 30282 18164 30288 18216
rect 30340 18204 30346 18216
rect 30837 18207 30895 18213
rect 30837 18204 30849 18207
rect 30340 18176 30849 18204
rect 30340 18164 30346 18176
rect 30837 18173 30849 18176
rect 30883 18173 30895 18207
rect 30837 18167 30895 18173
rect 31938 18164 31944 18216
rect 31996 18204 32002 18216
rect 32309 18207 32367 18213
rect 32309 18204 32321 18207
rect 31996 18176 32321 18204
rect 31996 18164 32002 18176
rect 32309 18173 32321 18176
rect 32355 18173 32367 18207
rect 34054 18204 34060 18216
rect 34015 18176 34060 18204
rect 32309 18167 32367 18173
rect 34054 18164 34060 18176
rect 34112 18164 34118 18216
rect 43530 18204 43536 18216
rect 43491 18176 43536 18204
rect 43530 18164 43536 18176
rect 43588 18164 43594 18216
rect 45186 18204 45192 18216
rect 45147 18176 45192 18204
rect 45186 18164 45192 18176
rect 45244 18164 45250 18216
rect 47044 18204 47072 18232
rect 47854 18204 47860 18216
rect 47044 18176 47860 18204
rect 47854 18164 47860 18176
rect 47912 18164 47918 18216
rect 25682 18136 25688 18148
rect 23768 18108 25688 18136
rect 25682 18096 25688 18108
rect 25740 18096 25746 18148
rect 28721 18139 28779 18145
rect 28721 18105 28733 18139
rect 28767 18136 28779 18139
rect 30374 18136 30380 18148
rect 28767 18108 30380 18136
rect 28767 18105 28779 18108
rect 28721 18099 28779 18105
rect 22646 18068 22652 18080
rect 19352 18040 22652 18068
rect 22646 18028 22652 18040
rect 22704 18028 22710 18080
rect 23109 18071 23167 18077
rect 23109 18037 23121 18071
rect 23155 18068 23167 18071
rect 23474 18068 23480 18080
rect 23155 18040 23480 18068
rect 23155 18037 23167 18040
rect 23109 18031 23167 18037
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 23753 18071 23811 18077
rect 23753 18037 23765 18071
rect 23799 18068 23811 18071
rect 24670 18068 24676 18080
rect 23799 18040 24676 18068
rect 23799 18037 23811 18040
rect 23753 18031 23811 18037
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 24854 18068 24860 18080
rect 24815 18040 24860 18068
rect 24854 18028 24860 18040
rect 24912 18028 24918 18080
rect 25958 18028 25964 18080
rect 26016 18068 26022 18080
rect 28736 18068 28764 18099
rect 30374 18096 30380 18108
rect 30432 18096 30438 18148
rect 35526 18096 35532 18148
rect 35584 18136 35590 18148
rect 46750 18136 46756 18148
rect 35584 18108 46756 18136
rect 35584 18096 35590 18108
rect 46750 18096 46756 18108
rect 46808 18096 46814 18148
rect 26016 18040 28764 18068
rect 26016 18028 26022 18040
rect 33134 18028 33140 18080
rect 33192 18068 33198 18080
rect 34609 18071 34667 18077
rect 34609 18068 34621 18071
rect 33192 18040 34621 18068
rect 33192 18028 33198 18040
rect 34609 18037 34621 18040
rect 34655 18037 34667 18071
rect 46290 18068 46296 18080
rect 46251 18040 46296 18068
rect 34609 18031 34667 18037
rect 46290 18028 46296 18040
rect 46348 18028 46354 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 14366 17824 14372 17876
rect 14424 17864 14430 17876
rect 14553 17867 14611 17873
rect 14553 17864 14565 17867
rect 14424 17836 14565 17864
rect 14424 17824 14430 17836
rect 14553 17833 14565 17836
rect 14599 17833 14611 17867
rect 14553 17827 14611 17833
rect 14568 17796 14596 17827
rect 14642 17824 14648 17876
rect 14700 17864 14706 17876
rect 14737 17867 14795 17873
rect 14737 17864 14749 17867
rect 14700 17836 14749 17864
rect 14700 17824 14706 17836
rect 14737 17833 14749 17836
rect 14783 17833 14795 17867
rect 14737 17827 14795 17833
rect 16850 17824 16856 17876
rect 16908 17864 16914 17876
rect 16945 17867 17003 17873
rect 16945 17864 16957 17867
rect 16908 17836 16957 17864
rect 16908 17824 16914 17836
rect 16945 17833 16957 17836
rect 16991 17833 17003 17867
rect 16945 17827 17003 17833
rect 17034 17824 17040 17876
rect 17092 17864 17098 17876
rect 22097 17867 22155 17873
rect 22097 17864 22109 17867
rect 17092 17836 22109 17864
rect 17092 17824 17098 17836
rect 22097 17833 22109 17836
rect 22143 17833 22155 17867
rect 22097 17827 22155 17833
rect 23290 17824 23296 17876
rect 23348 17864 23354 17876
rect 25590 17864 25596 17876
rect 23348 17836 24256 17864
rect 25551 17836 25596 17864
rect 23348 17824 23354 17836
rect 24026 17796 24032 17808
rect 14568 17768 14688 17796
rect 14660 17740 14688 17768
rect 21560 17768 24032 17796
rect 14642 17688 14648 17740
rect 14700 17688 14706 17740
rect 15010 17688 15016 17740
rect 15068 17728 15074 17740
rect 15197 17731 15255 17737
rect 15197 17728 15209 17731
rect 15068 17700 15209 17728
rect 15068 17688 15074 17700
rect 15197 17697 15209 17700
rect 15243 17697 15255 17731
rect 15470 17728 15476 17740
rect 15431 17700 15476 17728
rect 15197 17691 15255 17697
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 18414 17728 18420 17740
rect 18375 17700 18420 17728
rect 18414 17688 18420 17700
rect 18472 17688 18478 17740
rect 18693 17731 18751 17737
rect 18693 17697 18705 17731
rect 18739 17728 18751 17731
rect 19521 17731 19579 17737
rect 19521 17728 19533 17731
rect 18739 17700 19533 17728
rect 18739 17697 18751 17700
rect 18693 17691 18751 17697
rect 19521 17697 19533 17700
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 13173 17663 13231 17669
rect 13173 17629 13185 17663
rect 13219 17660 13231 17663
rect 13262 17660 13268 17672
rect 13219 17632 13268 17660
rect 13219 17629 13231 17632
rect 13173 17623 13231 17629
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17660 18383 17663
rect 19242 17660 19248 17672
rect 18371 17632 19104 17660
rect 19203 17632 19248 17660
rect 18371 17629 18383 17632
rect 18325 17623 18383 17629
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17592 14427 17595
rect 14734 17592 14740 17604
rect 14415 17564 14740 17592
rect 14415 17561 14427 17564
rect 14369 17555 14427 17561
rect 14734 17552 14740 17564
rect 14792 17592 14798 17604
rect 15010 17592 15016 17604
rect 14792 17564 15016 17592
rect 14792 17552 14798 17564
rect 15010 17552 15016 17564
rect 15068 17552 15074 17604
rect 19076 17536 19104 17632
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 21560 17604 21588 17768
rect 21729 17663 21787 17669
rect 21729 17629 21741 17663
rect 21775 17660 21787 17663
rect 21818 17660 21824 17672
rect 21775 17632 21824 17660
rect 21775 17629 21787 17632
rect 21729 17623 21787 17629
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 22741 17663 22799 17669
rect 22741 17629 22753 17663
rect 22787 17660 22799 17663
rect 23198 17660 23204 17672
rect 22787 17632 23204 17660
rect 22787 17629 22799 17632
rect 22741 17623 22799 17629
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 23308 17669 23336 17768
rect 24026 17756 24032 17768
rect 24084 17756 24090 17808
rect 23842 17688 23848 17740
rect 23900 17688 23906 17740
rect 24228 17728 24256 17836
rect 25590 17824 25596 17836
rect 25648 17824 25654 17876
rect 26513 17867 26571 17873
rect 26513 17833 26525 17867
rect 26559 17864 26571 17867
rect 26970 17864 26976 17876
rect 26559 17836 26976 17864
rect 26559 17833 26571 17836
rect 26513 17827 26571 17833
rect 26970 17824 26976 17836
rect 27028 17824 27034 17876
rect 43441 17867 43499 17873
rect 43441 17833 43453 17867
rect 43487 17864 43499 17867
rect 43530 17864 43536 17876
rect 43487 17836 43536 17864
rect 43487 17833 43499 17836
rect 43441 17827 43499 17833
rect 43530 17824 43536 17836
rect 43588 17824 43594 17876
rect 44174 17824 44180 17876
rect 44232 17864 44238 17876
rect 45649 17867 45707 17873
rect 45649 17864 45661 17867
rect 44232 17836 45661 17864
rect 44232 17824 44238 17836
rect 45649 17833 45661 17836
rect 45695 17833 45707 17867
rect 45649 17827 45707 17833
rect 24670 17796 24676 17808
rect 24631 17768 24676 17796
rect 24670 17756 24676 17768
rect 24728 17756 24734 17808
rect 35897 17799 35955 17805
rect 35897 17765 35909 17799
rect 35943 17796 35955 17799
rect 46382 17796 46388 17808
rect 35943 17768 46388 17796
rect 35943 17765 35955 17768
rect 35897 17759 35955 17765
rect 30282 17728 30288 17740
rect 24228 17700 26556 17728
rect 30243 17700 30288 17728
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17662 23535 17663
rect 23658 17662 23664 17672
rect 23523 17634 23664 17662
rect 23523 17629 23535 17634
rect 23477 17623 23535 17629
rect 23658 17620 23664 17634
rect 23716 17620 23722 17672
rect 23860 17660 23888 17688
rect 26528 17672 26556 17700
rect 30282 17688 30288 17700
rect 30340 17688 30346 17740
rect 30561 17731 30619 17737
rect 30561 17697 30573 17731
rect 30607 17728 30619 17731
rect 31110 17728 31116 17740
rect 30607 17700 31116 17728
rect 30607 17697 30619 17700
rect 30561 17691 30619 17697
rect 31110 17688 31116 17700
rect 31168 17728 31174 17740
rect 32217 17731 32275 17737
rect 32217 17728 32229 17731
rect 31168 17700 32229 17728
rect 31168 17688 31174 17700
rect 32217 17697 32229 17700
rect 32263 17697 32275 17731
rect 32217 17691 32275 17697
rect 32401 17731 32459 17737
rect 32401 17697 32413 17731
rect 32447 17728 32459 17731
rect 33134 17728 33140 17740
rect 32447 17700 33140 17728
rect 32447 17697 32459 17700
rect 32401 17691 32459 17697
rect 33134 17688 33140 17700
rect 33192 17688 33198 17740
rect 35526 17728 35532 17740
rect 35176 17700 35532 17728
rect 25498 17660 25504 17672
rect 23860 17632 24532 17660
rect 25459 17632 25504 17660
rect 20530 17552 20536 17604
rect 20588 17552 20594 17604
rect 21542 17592 21548 17604
rect 21503 17564 21548 17592
rect 21542 17552 21548 17564
rect 21600 17552 21606 17604
rect 21910 17592 21916 17604
rect 21871 17564 21916 17592
rect 21910 17552 21916 17564
rect 21968 17552 21974 17604
rect 23569 17595 23627 17601
rect 23569 17561 23581 17595
rect 23615 17561 23627 17595
rect 23569 17555 23627 17561
rect 13265 17527 13323 17533
rect 13265 17493 13277 17527
rect 13311 17524 13323 17527
rect 13446 17524 13452 17536
rect 13311 17496 13452 17524
rect 13311 17493 13323 17496
rect 13265 17487 13323 17493
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 14579 17527 14637 17533
rect 14579 17493 14591 17527
rect 14625 17524 14637 17527
rect 14918 17524 14924 17536
rect 14625 17496 14924 17524
rect 14625 17493 14637 17496
rect 14579 17487 14637 17493
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 19058 17484 19064 17536
rect 19116 17524 19122 17536
rect 20993 17527 21051 17533
rect 20993 17524 21005 17527
rect 19116 17496 21005 17524
rect 19116 17484 19122 17496
rect 20993 17493 21005 17496
rect 21039 17493 21051 17527
rect 20993 17487 21051 17493
rect 21818 17484 21824 17536
rect 21876 17524 21882 17536
rect 22741 17527 22799 17533
rect 21876 17496 21921 17524
rect 21876 17484 21882 17496
rect 22741 17493 22753 17527
rect 22787 17524 22799 17527
rect 23198 17524 23204 17536
rect 22787 17496 23204 17524
rect 22787 17493 22799 17496
rect 22741 17487 22799 17493
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23382 17484 23388 17536
rect 23440 17524 23446 17536
rect 23584 17524 23612 17555
rect 23750 17552 23756 17604
rect 23808 17592 23814 17604
rect 23845 17595 23903 17601
rect 23845 17592 23857 17595
rect 23808 17564 23857 17592
rect 23808 17552 23814 17564
rect 23845 17561 23857 17564
rect 23891 17592 23903 17595
rect 24397 17595 24455 17601
rect 24397 17592 24409 17595
rect 23891 17564 24409 17592
rect 23891 17561 23903 17564
rect 23845 17555 23903 17561
rect 24397 17561 24409 17564
rect 24443 17561 24455 17595
rect 24397 17555 24455 17561
rect 23440 17496 23612 17524
rect 23661 17527 23719 17533
rect 23440 17484 23446 17496
rect 23661 17493 23673 17527
rect 23707 17524 23719 17527
rect 23934 17524 23940 17536
rect 23707 17496 23940 17524
rect 23707 17493 23719 17496
rect 23661 17487 23719 17493
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 24504 17524 24532 17632
rect 25498 17620 25504 17632
rect 25556 17620 25562 17672
rect 25682 17660 25688 17672
rect 25643 17632 25688 17660
rect 25682 17620 25688 17632
rect 25740 17620 25746 17672
rect 26510 17660 26516 17672
rect 26471 17632 26516 17660
rect 26510 17620 26516 17632
rect 26568 17620 26574 17672
rect 30190 17660 30196 17672
rect 30151 17632 30196 17660
rect 30190 17620 30196 17632
rect 30248 17620 30254 17672
rect 35176 17669 35204 17700
rect 35526 17688 35532 17700
rect 35584 17688 35590 17740
rect 35161 17663 35219 17669
rect 35161 17629 35173 17663
rect 35207 17629 35219 17663
rect 35342 17660 35348 17672
rect 35303 17632 35348 17660
rect 35161 17623 35219 17629
rect 35342 17620 35348 17632
rect 35400 17620 35406 17672
rect 35437 17663 35495 17669
rect 35437 17629 35449 17663
rect 35483 17660 35495 17663
rect 35912 17660 35940 17759
rect 46382 17756 46388 17768
rect 46440 17756 46446 17808
rect 45373 17731 45431 17737
rect 45373 17728 45385 17731
rect 44468 17700 45385 17728
rect 35483 17632 35940 17660
rect 35483 17629 35495 17632
rect 35437 17623 35495 17629
rect 34054 17592 34060 17604
rect 34015 17564 34060 17592
rect 34054 17552 34060 17564
rect 34112 17552 34118 17604
rect 34793 17595 34851 17601
rect 34793 17561 34805 17595
rect 34839 17592 34851 17595
rect 35066 17592 35072 17604
rect 34839 17564 35072 17592
rect 34839 17561 34851 17564
rect 34793 17555 34851 17561
rect 35066 17552 35072 17564
rect 35124 17552 35130 17604
rect 24857 17527 24915 17533
rect 24857 17524 24869 17527
rect 24504 17496 24869 17524
rect 24857 17493 24869 17496
rect 24903 17493 24915 17527
rect 24857 17487 24915 17493
rect 26878 17484 26884 17536
rect 26936 17524 26942 17536
rect 35452 17524 35480 17623
rect 42794 17620 42800 17672
rect 42852 17660 42858 17672
rect 43349 17663 43407 17669
rect 43349 17660 43361 17663
rect 42852 17632 43361 17660
rect 42852 17620 42858 17632
rect 43349 17629 43361 17632
rect 43395 17660 43407 17663
rect 43530 17660 43536 17672
rect 43395 17632 43536 17660
rect 43395 17629 43407 17632
rect 43349 17623 43407 17629
rect 43530 17620 43536 17632
rect 43588 17620 43594 17672
rect 44468 17669 44496 17700
rect 45373 17697 45385 17700
rect 45419 17728 45431 17731
rect 45738 17728 45744 17740
rect 45419 17700 45744 17728
rect 45419 17697 45431 17700
rect 45373 17691 45431 17697
rect 45738 17688 45744 17700
rect 45796 17688 45802 17740
rect 46293 17731 46351 17737
rect 46293 17697 46305 17731
rect 46339 17728 46351 17731
rect 46842 17728 46848 17740
rect 46339 17700 46848 17728
rect 46339 17697 46351 17700
rect 46293 17691 46351 17697
rect 46842 17688 46848 17700
rect 46900 17688 46906 17740
rect 44269 17663 44327 17669
rect 44269 17629 44281 17663
rect 44315 17629 44327 17663
rect 44269 17623 44327 17629
rect 44453 17663 44511 17669
rect 44453 17629 44465 17663
rect 44499 17629 44511 17663
rect 44453 17623 44511 17629
rect 44284 17592 44312 17623
rect 44910 17620 44916 17672
rect 44968 17660 44974 17672
rect 45465 17663 45523 17669
rect 45465 17660 45477 17663
rect 44968 17632 45477 17660
rect 44968 17620 44974 17632
rect 45465 17629 45477 17632
rect 45511 17629 45523 17663
rect 45465 17623 45523 17629
rect 46477 17595 46535 17601
rect 44284 17564 45048 17592
rect 45020 17536 45048 17564
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 46934 17592 46940 17604
rect 46523 17564 46940 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 46934 17552 46940 17564
rect 46992 17552 46998 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 44358 17524 44364 17536
rect 26936 17496 35480 17524
rect 44319 17496 44364 17524
rect 26936 17484 26942 17496
rect 44358 17484 44364 17496
rect 44416 17484 44422 17536
rect 45002 17524 45008 17536
rect 44963 17496 45008 17524
rect 45002 17484 45008 17496
rect 45060 17484 45066 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1578 17280 1584 17332
rect 1636 17320 1642 17332
rect 26878 17320 26884 17332
rect 1636 17292 26884 17320
rect 1636 17280 1642 17292
rect 26878 17280 26884 17292
rect 26936 17280 26942 17332
rect 30282 17280 30288 17332
rect 30340 17320 30346 17332
rect 30561 17323 30619 17329
rect 30561 17320 30573 17323
rect 30340 17292 30573 17320
rect 30340 17280 30346 17292
rect 30561 17289 30573 17292
rect 30607 17289 30619 17323
rect 30561 17283 30619 17289
rect 34054 17280 34060 17332
rect 34112 17320 34118 17332
rect 44910 17320 44916 17332
rect 34112 17292 36768 17320
rect 34112 17280 34118 17292
rect 13725 17255 13783 17261
rect 13725 17221 13737 17255
rect 13771 17252 13783 17255
rect 13814 17252 13820 17264
rect 13771 17224 13820 17252
rect 13771 17221 13783 17224
rect 13725 17215 13783 17221
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 15749 17255 15807 17261
rect 15749 17252 15761 17255
rect 14950 17224 15761 17252
rect 15749 17221 15761 17224
rect 15795 17221 15807 17255
rect 15749 17215 15807 17221
rect 20349 17255 20407 17261
rect 20349 17221 20361 17255
rect 20395 17252 20407 17255
rect 20530 17252 20536 17264
rect 20395 17224 20536 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 21818 17212 21824 17264
rect 21876 17252 21882 17264
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 21876 17224 22201 17252
rect 21876 17212 21882 17224
rect 22189 17221 22201 17224
rect 22235 17221 22247 17255
rect 23474 17252 23480 17264
rect 23435 17224 23480 17252
rect 22189 17215 22247 17221
rect 23474 17212 23480 17224
rect 23532 17212 23538 17264
rect 24854 17252 24860 17264
rect 24702 17224 24860 17252
rect 24854 17212 24860 17224
rect 24912 17212 24918 17264
rect 29825 17255 29883 17261
rect 29825 17252 29837 17255
rect 28736 17224 29837 17252
rect 3418 17144 3424 17196
rect 3476 17184 3482 17196
rect 7926 17184 7932 17196
rect 3476 17156 7932 17184
rect 3476 17144 3482 17156
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 13446 17184 13452 17196
rect 13407 17156 13452 17184
rect 11977 17147 12035 17153
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11992 17116 12020 17147
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 15654 17184 15660 17196
rect 15615 17156 15660 17184
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 20257 17187 20315 17193
rect 20257 17153 20269 17187
rect 20303 17184 20315 17187
rect 20622 17184 20628 17196
rect 20303 17156 20628 17184
rect 20303 17153 20315 17156
rect 20257 17147 20315 17153
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22097 17187 22155 17193
rect 22097 17153 22109 17187
rect 22143 17184 22155 17187
rect 22646 17184 22652 17196
rect 22143 17156 22652 17184
rect 22143 17153 22155 17156
rect 22097 17147 22155 17153
rect 11112 17088 14780 17116
rect 11112 17076 11118 17088
rect 14752 17048 14780 17088
rect 15010 17076 15016 17128
rect 15068 17116 15074 17128
rect 15197 17119 15255 17125
rect 15197 17116 15209 17119
rect 15068 17088 15209 17116
rect 15068 17076 15074 17088
rect 15197 17085 15209 17088
rect 15243 17116 15255 17119
rect 16761 17119 16819 17125
rect 16761 17116 16773 17119
rect 15243 17088 16773 17116
rect 15243 17085 15255 17088
rect 15197 17079 15255 17085
rect 16761 17085 16773 17088
rect 16807 17085 16819 17119
rect 16942 17116 16948 17128
rect 16903 17088 16948 17116
rect 16761 17079 16819 17085
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 18601 17119 18659 17125
rect 18601 17085 18613 17119
rect 18647 17116 18659 17119
rect 19150 17116 19156 17128
rect 18647 17088 19156 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 16666 17048 16672 17060
rect 14752 17020 16672 17048
rect 16666 17008 16672 17020
rect 16724 17008 16730 17060
rect 21821 17051 21879 17057
rect 21821 17017 21833 17051
rect 21867 17017 21879 17051
rect 22020 17048 22048 17147
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 23198 17184 23204 17196
rect 23159 17156 23204 17184
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 27982 17144 27988 17196
rect 28040 17184 28046 17196
rect 28077 17187 28135 17193
rect 28077 17184 28089 17187
rect 28040 17156 28089 17184
rect 28040 17144 28046 17156
rect 28077 17153 28089 17156
rect 28123 17153 28135 17187
rect 28258 17184 28264 17196
rect 28219 17156 28264 17184
rect 28077 17147 28135 17153
rect 28258 17144 28264 17156
rect 28316 17144 28322 17196
rect 28534 17144 28540 17196
rect 28592 17184 28598 17196
rect 28736 17193 28764 17224
rect 29825 17221 29837 17224
rect 29871 17221 29883 17255
rect 35066 17252 35072 17264
rect 35027 17224 35072 17252
rect 29825 17215 29883 17221
rect 35066 17212 35072 17224
rect 35124 17212 35130 17264
rect 28721 17187 28779 17193
rect 28721 17184 28733 17187
rect 28592 17156 28733 17184
rect 28592 17144 28598 17156
rect 28721 17153 28733 17156
rect 28767 17153 28779 17187
rect 29641 17187 29699 17193
rect 29641 17184 29653 17187
rect 28721 17147 28779 17153
rect 28828 17156 29653 17184
rect 24026 17076 24032 17128
rect 24084 17116 24090 17128
rect 24949 17119 25007 17125
rect 24949 17116 24961 17119
rect 24084 17088 24961 17116
rect 24084 17076 24090 17088
rect 24949 17085 24961 17088
rect 24995 17085 25007 17119
rect 24949 17079 25007 17085
rect 22094 17048 22100 17060
rect 22020 17020 22100 17048
rect 21821 17011 21879 17017
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 12069 16983 12127 16989
rect 12069 16980 12081 16983
rect 11940 16952 12081 16980
rect 11940 16940 11946 16952
rect 12069 16949 12081 16952
rect 12115 16949 12127 16983
rect 12069 16943 12127 16949
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 21542 16980 21548 16992
rect 14424 16952 21548 16980
rect 14424 16940 14430 16952
rect 21542 16940 21548 16952
rect 21600 16980 21606 16992
rect 21836 16980 21864 17011
rect 22094 17008 22100 17020
rect 22152 17008 22158 17060
rect 27706 17008 27712 17060
rect 27764 17048 27770 17060
rect 28828 17057 28856 17156
rect 29641 17153 29653 17156
rect 29687 17153 29699 17187
rect 29641 17147 29699 17153
rect 30009 17187 30067 17193
rect 30009 17153 30021 17187
rect 30055 17184 30067 17187
rect 30469 17187 30527 17193
rect 30469 17184 30481 17187
rect 30055 17156 30481 17184
rect 30055 17153 30067 17156
rect 30009 17147 30067 17153
rect 30469 17153 30481 17156
rect 30515 17153 30527 17187
rect 30469 17147 30527 17153
rect 30653 17187 30711 17193
rect 30653 17153 30665 17187
rect 30699 17153 30711 17187
rect 30653 17147 30711 17153
rect 28994 17116 29000 17128
rect 28955 17088 29000 17116
rect 28994 17076 29000 17088
rect 29052 17076 29058 17128
rect 29089 17119 29147 17125
rect 29089 17085 29101 17119
rect 29135 17085 29147 17119
rect 29089 17079 29147 17085
rect 28813 17051 28871 17057
rect 28813 17048 28825 17051
rect 27764 17020 28825 17048
rect 27764 17008 27770 17020
rect 28813 17017 28825 17020
rect 28859 17017 28871 17051
rect 29104 17048 29132 17079
rect 29454 17076 29460 17128
rect 29512 17116 29518 17128
rect 30668 17116 30696 17147
rect 36740 17125 36768 17292
rect 43732 17292 44916 17320
rect 43732 17196 43760 17292
rect 44910 17280 44916 17292
rect 44968 17280 44974 17332
rect 45002 17280 45008 17332
rect 45060 17320 45066 17332
rect 47949 17323 48007 17329
rect 47949 17320 47961 17323
rect 45060 17292 47961 17320
rect 45060 17280 45066 17292
rect 47949 17289 47961 17292
rect 47995 17289 48007 17323
rect 47949 17283 48007 17289
rect 44450 17212 44456 17264
rect 44508 17252 44514 17264
rect 45373 17255 45431 17261
rect 44508 17224 45232 17252
rect 44508 17212 44514 17224
rect 44364 17196 44416 17202
rect 43714 17184 43720 17196
rect 43675 17156 43720 17184
rect 43714 17144 43720 17156
rect 43772 17144 43778 17196
rect 45204 17193 45232 17224
rect 45373 17221 45385 17255
rect 45419 17252 45431 17255
rect 46290 17252 46296 17264
rect 45419 17224 46296 17252
rect 45419 17221 45431 17224
rect 45373 17215 45431 17221
rect 46290 17212 46296 17224
rect 46348 17212 46354 17264
rect 47765 17255 47823 17261
rect 47765 17252 47777 17255
rect 46584 17224 47777 17252
rect 45189 17187 45247 17193
rect 45189 17153 45201 17187
rect 45235 17153 45247 17187
rect 45189 17147 45247 17153
rect 44364 17138 44416 17144
rect 29512 17088 30696 17116
rect 34885 17119 34943 17125
rect 29512 17076 29518 17088
rect 34885 17085 34897 17119
rect 34931 17085 34943 17119
rect 34885 17079 34943 17085
rect 36725 17119 36783 17125
rect 36725 17085 36737 17119
rect 36771 17116 36783 17119
rect 41414 17116 41420 17128
rect 36771 17088 41420 17116
rect 36771 17085 36783 17088
rect 36725 17079 36783 17085
rect 30006 17048 30012 17060
rect 29104 17020 30012 17048
rect 28813 17011 28871 17017
rect 30006 17008 30012 17020
rect 30064 17008 30070 17060
rect 30650 17008 30656 17060
rect 30708 17048 30714 17060
rect 34900 17048 34928 17079
rect 41414 17076 41420 17088
rect 41472 17116 41478 17128
rect 41472 17088 44312 17116
rect 41472 17076 41478 17088
rect 42794 17048 42800 17060
rect 30708 17020 42800 17048
rect 30708 17008 30714 17020
rect 42794 17008 42800 17020
rect 42852 17008 42858 17060
rect 44284 17048 44312 17088
rect 45646 17076 45652 17128
rect 45704 17116 45710 17128
rect 46584 17116 46612 17224
rect 47765 17221 47777 17224
rect 47811 17221 47823 17255
rect 47765 17215 47823 17221
rect 46658 17144 46664 17196
rect 46716 17184 46722 17196
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 46716 17156 47593 17184
rect 46716 17144 46722 17156
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 45704 17088 46612 17116
rect 46753 17119 46811 17125
rect 45704 17076 45710 17088
rect 46753 17085 46765 17119
rect 46799 17116 46811 17119
rect 47026 17116 47032 17128
rect 46799 17088 47032 17116
rect 46799 17085 46811 17088
rect 46753 17079 46811 17085
rect 46768 17048 46796 17079
rect 47026 17076 47032 17088
rect 47084 17076 47090 17128
rect 44284 17020 46796 17048
rect 21600 16952 21864 16980
rect 21600 16940 21606 16952
rect 22002 16940 22008 16992
rect 22060 16980 22066 16992
rect 22373 16983 22431 16989
rect 22373 16980 22385 16983
rect 22060 16952 22385 16980
rect 22060 16940 22066 16952
rect 22373 16949 22385 16952
rect 22419 16949 22431 16983
rect 28074 16980 28080 16992
rect 28035 16952 28080 16980
rect 22373 16943 22431 16949
rect 28074 16940 28080 16952
rect 28132 16940 28138 16992
rect 29178 16980 29184 16992
rect 29139 16952 29184 16980
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 14366 16776 14372 16788
rect 11716 16748 14372 16776
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 11716 16649 11744 16748
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 14550 16776 14556 16788
rect 14511 16748 14556 16776
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 17037 16779 17095 16785
rect 17037 16776 17049 16779
rect 17000 16748 17049 16776
rect 17000 16736 17006 16748
rect 17037 16745 17049 16748
rect 17083 16745 17095 16779
rect 17037 16739 17095 16745
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 22336 16748 22477 16776
rect 22336 16736 22342 16748
rect 22465 16745 22477 16748
rect 22511 16745 22523 16779
rect 28534 16776 28540 16788
rect 22465 16739 22523 16745
rect 28092 16748 28540 16776
rect 17218 16708 17224 16720
rect 17052 16680 17224 16708
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16609 11759 16643
rect 11882 16640 11888 16652
rect 11843 16612 11888 16640
rect 11701 16603 11759 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 15010 16640 15016 16652
rect 14568 16612 15016 16640
rect 11054 16582 11060 16594
rect 11015 16554 11060 16582
rect 11054 16542 11060 16554
rect 11112 16542 11118 16594
rect 14568 16581 14596 16612
rect 15010 16600 15016 16612
rect 15068 16600 15074 16652
rect 17052 16640 17080 16680
rect 17218 16668 17224 16680
rect 17276 16708 17282 16720
rect 18598 16708 18604 16720
rect 17276 16680 18604 16708
rect 17276 16668 17282 16680
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 21818 16668 21824 16720
rect 21876 16708 21882 16720
rect 22649 16711 22707 16717
rect 22649 16708 22661 16711
rect 21876 16680 22661 16708
rect 21876 16668 21882 16680
rect 22649 16677 22661 16680
rect 22695 16677 22707 16711
rect 28092 16708 28120 16748
rect 28534 16736 28540 16748
rect 28592 16736 28598 16788
rect 45738 16776 45744 16788
rect 45699 16748 45744 16776
rect 45738 16736 45744 16748
rect 45796 16736 45802 16788
rect 22649 16671 22707 16677
rect 28000 16680 28120 16708
rect 28445 16711 28503 16717
rect 16960 16612 17080 16640
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 14829 16575 14887 16581
rect 14829 16541 14841 16575
rect 14875 16572 14887 16575
rect 14918 16572 14924 16584
rect 14875 16544 14924 16572
rect 14875 16541 14887 16544
rect 14829 16535 14887 16541
rect 14918 16532 14924 16544
rect 14976 16532 14982 16584
rect 16960 16581 16988 16612
rect 18414 16600 18420 16652
rect 18472 16640 18478 16652
rect 22094 16640 22100 16652
rect 18472 16612 21588 16640
rect 18472 16600 18478 16612
rect 16945 16575 17003 16581
rect 16945 16541 16957 16575
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 3510 16464 3516 16516
rect 3568 16504 3574 16516
rect 13541 16507 13599 16513
rect 13541 16504 13553 16507
rect 3568 16476 13553 16504
rect 3568 16464 3574 16476
rect 13541 16473 13553 16476
rect 13587 16473 13599 16507
rect 21560 16504 21588 16612
rect 21652 16612 22100 16640
rect 21652 16581 21680 16612
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 23290 16600 23296 16652
rect 23348 16640 23354 16652
rect 23348 16612 24440 16640
rect 23348 16600 23354 16612
rect 21637 16575 21695 16581
rect 21637 16541 21649 16575
rect 21683 16541 21695 16575
rect 21637 16535 21695 16541
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16572 21879 16575
rect 22002 16572 22008 16584
rect 21867 16544 22008 16572
rect 21867 16541 21879 16544
rect 21821 16535 21879 16541
rect 21836 16504 21864 16535
rect 22002 16532 22008 16544
rect 22060 16532 22066 16584
rect 24412 16581 24440 16612
rect 24397 16575 24455 16581
rect 24397 16541 24409 16575
rect 24443 16541 24455 16575
rect 27154 16572 27160 16584
rect 27115 16544 27160 16572
rect 24397 16535 24455 16541
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 27246 16532 27252 16584
rect 27304 16572 27310 16584
rect 27341 16575 27399 16581
rect 27341 16572 27353 16575
rect 27304 16544 27353 16572
rect 27304 16532 27310 16544
rect 27341 16541 27353 16544
rect 27387 16541 27399 16575
rect 27341 16535 27399 16541
rect 27706 16532 27712 16584
rect 27764 16572 27770 16584
rect 28000 16581 28028 16680
rect 28445 16677 28457 16711
rect 28491 16708 28503 16711
rect 28491 16680 31754 16708
rect 28491 16677 28503 16680
rect 28445 16671 28503 16677
rect 28074 16600 28080 16652
rect 28132 16640 28138 16652
rect 29733 16643 29791 16649
rect 29733 16640 29745 16643
rect 28132 16612 29745 16640
rect 28132 16600 28138 16612
rect 29733 16609 29745 16612
rect 29779 16609 29791 16643
rect 30650 16640 30656 16652
rect 30611 16612 30656 16640
rect 29733 16603 29791 16609
rect 30650 16600 30656 16612
rect 30708 16600 30714 16652
rect 31726 16640 31754 16680
rect 45646 16668 45652 16720
rect 45704 16668 45710 16720
rect 43714 16640 43720 16652
rect 31726 16612 43720 16640
rect 43714 16600 43720 16612
rect 43772 16600 43778 16652
rect 45664 16640 45692 16668
rect 46293 16643 46351 16649
rect 45664 16612 45876 16640
rect 27801 16575 27859 16581
rect 27801 16572 27813 16575
rect 27764 16544 27813 16572
rect 27764 16532 27770 16544
rect 27801 16541 27813 16544
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 27985 16575 28043 16581
rect 27985 16541 27997 16575
rect 28031 16541 28043 16575
rect 29822 16572 29828 16584
rect 27985 16535 28043 16541
rect 28184 16544 28764 16572
rect 29783 16544 29828 16572
rect 21560 16476 21864 16504
rect 22281 16507 22339 16513
rect 13541 16467 13599 16473
rect 22281 16473 22293 16507
rect 22327 16504 22339 16507
rect 22370 16504 22376 16516
rect 22327 16476 22376 16504
rect 22327 16473 22339 16476
rect 22281 16467 22339 16473
rect 22370 16464 22376 16476
rect 22428 16464 22434 16516
rect 22497 16507 22555 16513
rect 22497 16473 22509 16507
rect 22543 16504 22555 16507
rect 23658 16504 23664 16516
rect 22543 16476 23664 16504
rect 22543 16473 22555 16476
rect 22497 16467 22555 16473
rect 23658 16464 23664 16476
rect 23716 16464 23722 16516
rect 28184 16504 28212 16544
rect 28626 16504 28632 16516
rect 27816 16476 28212 16504
rect 28587 16476 28632 16504
rect 27816 16448 27844 16476
rect 28626 16464 28632 16476
rect 28684 16464 28690 16516
rect 28736 16504 28764 16544
rect 29822 16532 29828 16544
rect 29880 16532 29886 16584
rect 35986 16532 35992 16584
rect 36044 16572 36050 16584
rect 36538 16572 36544 16584
rect 36044 16544 36544 16572
rect 36044 16532 36050 16544
rect 36538 16532 36544 16544
rect 36596 16532 36602 16584
rect 45848 16581 45876 16612
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47486 16640 47492 16652
rect 46339 16612 47492 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47486 16600 47492 16612
rect 47544 16600 47550 16652
rect 45649 16575 45707 16581
rect 45649 16541 45661 16575
rect 45695 16541 45707 16575
rect 45649 16535 45707 16541
rect 45833 16575 45891 16581
rect 45833 16541 45845 16575
rect 45879 16541 45891 16575
rect 45833 16535 45891 16541
rect 28997 16507 29055 16513
rect 28997 16504 29009 16507
rect 28736 16476 28856 16504
rect 11149 16439 11207 16445
rect 11149 16405 11161 16439
rect 11195 16436 11207 16439
rect 11698 16436 11704 16448
rect 11195 16408 11704 16436
rect 11195 16405 11207 16408
rect 11149 16399 11207 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 14734 16436 14740 16448
rect 14695 16408 14740 16436
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 21542 16396 21548 16448
rect 21600 16436 21606 16448
rect 21729 16439 21787 16445
rect 21729 16436 21741 16439
rect 21600 16408 21741 16436
rect 21600 16396 21606 16408
rect 21729 16405 21741 16408
rect 21775 16405 21787 16439
rect 21729 16399 21787 16405
rect 23842 16396 23848 16448
rect 23900 16436 23906 16448
rect 24489 16439 24547 16445
rect 24489 16436 24501 16439
rect 23900 16408 24501 16436
rect 23900 16396 23906 16408
rect 24489 16405 24501 16408
rect 24535 16405 24547 16439
rect 24489 16399 24547 16405
rect 27341 16439 27399 16445
rect 27341 16405 27353 16439
rect 27387 16436 27399 16439
rect 27798 16436 27804 16448
rect 27387 16408 27804 16436
rect 27387 16405 27399 16408
rect 27341 16399 27399 16405
rect 27798 16396 27804 16408
rect 27856 16396 27862 16448
rect 27985 16439 28043 16445
rect 27985 16405 27997 16439
rect 28031 16436 28043 16439
rect 28718 16436 28724 16448
rect 28031 16408 28724 16436
rect 28031 16405 28043 16408
rect 27985 16399 28043 16405
rect 28718 16396 28724 16408
rect 28776 16396 28782 16448
rect 28828 16445 28856 16476
rect 28920 16476 29009 16504
rect 28920 16448 28948 16476
rect 28997 16473 29009 16476
rect 29043 16473 29055 16507
rect 28997 16467 29055 16473
rect 28813 16439 28871 16445
rect 28813 16405 28825 16439
rect 28859 16405 28871 16439
rect 28813 16399 28871 16405
rect 28902 16396 28908 16448
rect 28960 16396 28966 16448
rect 45664 16436 45692 16535
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 48130 16504 48136 16516
rect 48091 16476 48136 16504
rect 48130 16464 48136 16476
rect 48188 16464 48194 16516
rect 46566 16436 46572 16448
rect 45664 16408 46572 16436
rect 46566 16396 46572 16408
rect 46624 16396 46630 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 19889 16235 19947 16241
rect 6886 16204 19840 16232
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16096 2099 16099
rect 6886 16096 6914 16204
rect 11698 16164 11704 16176
rect 11659 16136 11704 16164
rect 11698 16124 11704 16136
rect 11756 16124 11762 16176
rect 16868 16136 18368 16164
rect 11514 16096 11520 16108
rect 2087 16068 6914 16096
rect 11475 16068 11520 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 16868 16105 16896 16136
rect 15105 16099 15163 16105
rect 15105 16065 15117 16099
rect 15151 16096 15163 16099
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 15151 16068 16865 16096
rect 15151 16065 15163 16068
rect 15105 16059 15163 16065
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12492 16000 12537 16028
rect 12492 15988 12498 16000
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 17420 16028 17448 16059
rect 15712 16000 17448 16028
rect 18340 16028 18368 16136
rect 18598 16124 18604 16176
rect 18656 16164 18662 16176
rect 19242 16164 19248 16176
rect 18656 16136 19248 16164
rect 18656 16124 18662 16136
rect 19242 16124 19248 16136
rect 19300 16164 19306 16176
rect 19521 16167 19579 16173
rect 19521 16164 19533 16167
rect 19300 16136 19533 16164
rect 19300 16124 19306 16136
rect 19521 16133 19533 16136
rect 19567 16133 19579 16167
rect 19721 16167 19779 16173
rect 19721 16164 19733 16167
rect 19521 16127 19579 16133
rect 19628 16136 19733 16164
rect 18414 16056 18420 16108
rect 18472 16096 18478 16108
rect 18874 16096 18880 16108
rect 18472 16068 18880 16096
rect 18472 16056 18478 16068
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 19058 16096 19064 16108
rect 19019 16068 19064 16096
rect 19058 16056 19064 16068
rect 19116 16096 19122 16108
rect 19628 16096 19656 16136
rect 19721 16133 19733 16136
rect 19767 16133 19779 16167
rect 19812 16164 19840 16204
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 21910 16232 21916 16244
rect 19935 16204 21916 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 22281 16235 22339 16241
rect 22281 16201 22293 16235
rect 22327 16232 22339 16235
rect 22370 16232 22376 16244
rect 22327 16204 22376 16232
rect 22327 16201 22339 16204
rect 22281 16195 22339 16201
rect 22370 16192 22376 16204
rect 22428 16232 22434 16244
rect 25593 16235 25651 16241
rect 25593 16232 25605 16235
rect 22428 16204 25605 16232
rect 22428 16192 22434 16204
rect 20714 16164 20720 16176
rect 19812 16136 20720 16164
rect 19721 16127 19779 16133
rect 20714 16124 20720 16136
rect 20772 16124 20778 16176
rect 22097 16167 22155 16173
rect 22097 16133 22109 16167
rect 22143 16164 22155 16167
rect 22462 16164 22468 16176
rect 22143 16136 22468 16164
rect 22143 16133 22155 16136
rect 22097 16127 22155 16133
rect 22462 16124 22468 16136
rect 22520 16124 22526 16176
rect 19116 16068 19656 16096
rect 20533 16099 20591 16105
rect 19116 16056 19122 16068
rect 20533 16065 20545 16099
rect 20579 16096 20591 16099
rect 20622 16096 20628 16108
rect 20579 16068 20628 16096
rect 20579 16065 20591 16068
rect 20533 16059 20591 16065
rect 20622 16056 20628 16068
rect 20680 16096 20686 16108
rect 22002 16096 22008 16108
rect 20680 16068 22008 16096
rect 20680 16056 20686 16068
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16065 22431 16099
rect 22940 16096 22968 16204
rect 25593 16201 25605 16204
rect 25639 16201 25651 16235
rect 25593 16195 25651 16201
rect 27249 16235 27307 16241
rect 27249 16201 27261 16235
rect 27295 16232 27307 16235
rect 27982 16232 27988 16244
rect 27295 16204 27988 16232
rect 27295 16201 27307 16204
rect 27249 16195 27307 16201
rect 27982 16192 27988 16204
rect 28040 16192 28046 16244
rect 28258 16192 28264 16244
rect 28316 16232 28322 16244
rect 28537 16235 28595 16241
rect 28537 16232 28549 16235
rect 28316 16204 28549 16232
rect 28316 16192 28322 16204
rect 28537 16201 28549 16204
rect 28583 16201 28595 16235
rect 28537 16195 28595 16201
rect 29457 16235 29515 16241
rect 29457 16201 29469 16235
rect 29503 16232 29515 16235
rect 29822 16232 29828 16244
rect 29503 16204 29828 16232
rect 29503 16201 29515 16204
rect 29457 16195 29515 16201
rect 29822 16192 29828 16204
rect 29880 16192 29886 16244
rect 36538 16192 36544 16244
rect 36596 16232 36602 16244
rect 46934 16232 46940 16244
rect 36596 16204 44772 16232
rect 46895 16204 46940 16232
rect 36596 16192 36602 16204
rect 24762 16124 24768 16176
rect 24820 16124 24826 16176
rect 28000 16164 28028 16192
rect 28902 16164 28908 16176
rect 28000 16136 28908 16164
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 43901 16167 43959 16173
rect 43901 16133 43913 16167
rect 43947 16164 43959 16167
rect 44637 16167 44695 16173
rect 44637 16164 44649 16167
rect 43947 16136 44649 16164
rect 43947 16133 43959 16136
rect 43901 16127 43959 16133
rect 44637 16133 44649 16136
rect 44683 16133 44695 16167
rect 44744 16164 44772 16204
rect 46934 16192 46940 16204
rect 46992 16192 46998 16244
rect 47670 16232 47676 16244
rect 47631 16204 47676 16232
rect 47670 16192 47676 16204
rect 47728 16192 47734 16244
rect 44744 16136 47624 16164
rect 44637 16127 44695 16133
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 22940 16068 23029 16096
rect 22373 16059 22431 16065
rect 23017 16065 23029 16068
rect 23063 16065 23075 16099
rect 23842 16096 23848 16108
rect 23803 16068 23848 16096
rect 23017 16059 23075 16065
rect 19978 16028 19984 16040
rect 18340 16000 19984 16028
rect 15712 15988 15718 16000
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 22388 16028 22416 16059
rect 23842 16056 23848 16068
rect 23900 16056 23906 16108
rect 27154 16096 27160 16108
rect 27067 16068 27160 16096
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27246 16056 27252 16108
rect 27304 16096 27310 16108
rect 27341 16099 27399 16105
rect 27341 16096 27353 16099
rect 27304 16068 27353 16096
rect 27304 16056 27310 16068
rect 27341 16065 27353 16068
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 27798 16056 27804 16108
rect 27856 16096 27862 16108
rect 28445 16099 28503 16105
rect 28445 16096 28457 16099
rect 27856 16068 28457 16096
rect 27856 16056 27862 16068
rect 28445 16065 28457 16068
rect 28491 16065 28503 16099
rect 28445 16059 28503 16065
rect 28626 16056 28632 16108
rect 28684 16096 28690 16108
rect 29178 16096 29184 16108
rect 28684 16068 29184 16096
rect 28684 16056 28690 16068
rect 29178 16056 29184 16068
rect 29236 16096 29242 16108
rect 29273 16099 29331 16105
rect 29273 16096 29285 16099
rect 29236 16068 29285 16096
rect 29236 16056 29242 16068
rect 29273 16065 29285 16068
rect 29319 16065 29331 16099
rect 29273 16059 29331 16065
rect 43809 16099 43867 16105
rect 43809 16065 43821 16099
rect 43855 16065 43867 16099
rect 44450 16096 44456 16108
rect 44411 16068 44456 16096
rect 43809 16059 43867 16065
rect 23109 16031 23167 16037
rect 23109 16028 23121 16031
rect 22388 16000 23121 16028
rect 23109 15997 23121 16000
rect 23155 16028 23167 16031
rect 23750 16028 23756 16040
rect 23155 16000 23756 16028
rect 23155 15997 23167 16000
rect 23109 15991 23167 15997
rect 23750 15988 23756 16000
rect 23808 15988 23814 16040
rect 24121 16031 24179 16037
rect 24121 16028 24133 16031
rect 23952 16000 24133 16028
rect 19150 15920 19156 15972
rect 19208 15960 19214 15972
rect 19208 15932 20760 15960
rect 19208 15920 19214 15932
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 15197 15895 15255 15901
rect 15197 15892 15209 15895
rect 14608 15864 15209 15892
rect 14608 15852 14614 15864
rect 15197 15861 15209 15864
rect 15243 15861 15255 15895
rect 16850 15892 16856 15904
rect 16811 15864 16856 15892
rect 15197 15855 15255 15861
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 17497 15895 17555 15901
rect 17497 15861 17509 15895
rect 17543 15892 17555 15895
rect 17586 15892 17592 15904
rect 17543 15864 17592 15892
rect 17543 15861 17555 15864
rect 17497 15855 17555 15861
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 18969 15895 19027 15901
rect 18969 15861 18981 15895
rect 19015 15892 19027 15895
rect 19334 15892 19340 15904
rect 19015 15864 19340 15892
rect 19015 15861 19027 15864
rect 18969 15855 19027 15861
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 19705 15895 19763 15901
rect 19705 15892 19717 15895
rect 19484 15864 19717 15892
rect 19484 15852 19490 15864
rect 19705 15861 19717 15864
rect 19751 15861 19763 15895
rect 20622 15892 20628 15904
rect 20583 15864 20628 15892
rect 19705 15855 19763 15861
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 20732 15892 20760 15932
rect 22094 15920 22100 15972
rect 22152 15960 22158 15972
rect 23385 15963 23443 15969
rect 22152 15932 22197 15960
rect 22152 15920 22158 15932
rect 23385 15929 23397 15963
rect 23431 15960 23443 15963
rect 23952 15960 23980 16000
rect 24121 15997 24133 16000
rect 24167 15997 24179 16031
rect 24121 15991 24179 15997
rect 24578 15988 24584 16040
rect 24636 16028 24642 16040
rect 27172 16028 27200 16056
rect 24636 16000 27200 16028
rect 24636 15988 24642 16000
rect 28718 15988 28724 16040
rect 28776 16028 28782 16040
rect 29089 16031 29147 16037
rect 29089 16028 29101 16031
rect 28776 16000 29101 16028
rect 28776 15988 28782 16000
rect 29089 15997 29101 16000
rect 29135 16028 29147 16031
rect 29454 16028 29460 16040
rect 29135 16000 29460 16028
rect 29135 15997 29147 16000
rect 29089 15991 29147 15997
rect 29454 15988 29460 16000
rect 29512 15988 29518 16040
rect 43824 16028 43852 16059
rect 44450 16056 44456 16068
rect 44508 16056 44514 16108
rect 46845 16099 46903 16105
rect 46845 16065 46857 16099
rect 46891 16096 46903 16099
rect 47118 16096 47124 16108
rect 46891 16068 47124 16096
rect 46891 16065 46903 16068
rect 46845 16059 46903 16065
rect 47118 16056 47124 16068
rect 47176 16096 47182 16108
rect 47394 16096 47400 16108
rect 47176 16068 47400 16096
rect 47176 16056 47182 16068
rect 47394 16056 47400 16068
rect 47452 16056 47458 16108
rect 47596 16105 47624 16136
rect 47581 16099 47639 16105
rect 47581 16065 47593 16099
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 45554 16028 45560 16040
rect 43824 16000 45560 16028
rect 45554 15988 45560 16000
rect 45612 15988 45618 16040
rect 46106 16028 46112 16040
rect 46067 16000 46112 16028
rect 46106 15988 46112 16000
rect 46164 15988 46170 16040
rect 23431 15932 23980 15960
rect 45572 15960 45600 15988
rect 47118 15960 47124 15972
rect 45572 15932 47124 15960
rect 23431 15929 23443 15932
rect 23385 15923 23443 15929
rect 47118 15920 47124 15932
rect 47176 15920 47182 15972
rect 25498 15892 25504 15904
rect 20732 15864 25504 15892
rect 25498 15852 25504 15864
rect 25556 15852 25562 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 24578 15688 24584 15700
rect 6886 15660 24584 15688
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 6886 15552 6914 15660
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 25498 15648 25504 15700
rect 25556 15688 25562 15700
rect 45554 15688 45560 15700
rect 25556 15660 45560 15688
rect 25556 15648 25562 15660
rect 45554 15648 45560 15660
rect 45612 15648 45618 15700
rect 47486 15648 47492 15700
rect 47544 15688 47550 15700
rect 47673 15691 47731 15697
rect 47673 15688 47685 15691
rect 47544 15660 47685 15688
rect 47544 15648 47550 15660
rect 47673 15657 47685 15660
rect 47719 15657 47731 15691
rect 47673 15651 47731 15657
rect 18598 15620 18604 15632
rect 18559 15592 18604 15620
rect 18598 15580 18604 15592
rect 18656 15580 18662 15632
rect 14550 15552 14556 15564
rect 5500 15524 6914 15552
rect 14511 15524 14556 15552
rect 5500 15512 5506 15524
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 16850 15552 16856 15564
rect 16811 15524 16856 15552
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 19334 15552 19340 15564
rect 19295 15524 19340 15552
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 21542 15552 21548 15564
rect 21503 15524 21548 15552
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 2041 15447 2099 15453
rect 19352 15456 19441 15484
rect 19352 15428 19380 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19978 15444 19984 15496
rect 20036 15484 20042 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20036 15456 20545 15484
rect 20036 15444 20042 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15484 20867 15487
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 20855 15456 21281 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 24670 15484 24676 15496
rect 24631 15456 24676 15484
rect 21269 15447 21327 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 43530 15484 43536 15496
rect 43491 15456 43536 15484
rect 43530 15444 43536 15456
rect 43588 15444 43594 15496
rect 14826 15416 14832 15428
rect 14787 15388 14832 15416
rect 14826 15376 14832 15388
rect 14884 15376 14890 15428
rect 15562 15376 15568 15428
rect 15620 15376 15626 15428
rect 17126 15416 17132 15428
rect 17087 15388 17132 15416
rect 17126 15376 17132 15388
rect 17184 15376 17190 15428
rect 17586 15376 17592 15428
rect 17644 15376 17650 15428
rect 19334 15376 19340 15428
rect 19392 15376 19398 15428
rect 22278 15376 22284 15428
rect 22336 15376 22342 15428
rect 16298 15348 16304 15360
rect 16259 15320 16304 15348
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 19484 15320 19809 15348
rect 19484 15308 19490 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 19797 15311 19855 15317
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 23017 15351 23075 15357
rect 23017 15348 23029 15351
rect 22520 15320 23029 15348
rect 22520 15308 22526 15320
rect 23017 15317 23029 15320
rect 23063 15317 23075 15351
rect 23017 15311 23075 15317
rect 43625 15351 43683 15357
rect 43625 15317 43637 15351
rect 43671 15348 43683 15351
rect 43806 15348 43812 15360
rect 43671 15320 43812 15348
rect 43671 15317 43683 15320
rect 43625 15311 43683 15317
rect 43806 15308 43812 15320
rect 43864 15308 43870 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 15562 15144 15568 15156
rect 15523 15116 15568 15144
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 17126 15104 17132 15156
rect 17184 15144 17190 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 17184 15116 17325 15144
rect 17184 15104 17190 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 17313 15107 17371 15113
rect 17880 15116 18797 15144
rect 14734 15076 14740 15088
rect 14292 15048 14740 15076
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 14292 15017 14320 15048
rect 14734 15036 14740 15048
rect 14792 15076 14798 15088
rect 16298 15076 16304 15088
rect 14792 15048 16304 15076
rect 14792 15036 14798 15048
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 15008 15531 15011
rect 15654 15008 15660 15020
rect 15519 14980 15660 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17773 15011 17831 15017
rect 17773 14977 17785 15011
rect 17819 15008 17831 15011
rect 17880 15008 17908 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 22278 15104 22284 15156
rect 22336 15144 22342 15156
rect 22373 15147 22431 15153
rect 22373 15144 22385 15147
rect 22336 15116 22385 15144
rect 22336 15104 22342 15116
rect 22373 15113 22385 15116
rect 22419 15113 22431 15147
rect 22373 15107 22431 15113
rect 18414 15076 18420 15088
rect 18375 15048 18420 15076
rect 18414 15036 18420 15048
rect 18472 15036 18478 15088
rect 18633 15079 18691 15085
rect 18633 15045 18645 15079
rect 18679 15076 18691 15079
rect 18874 15076 18880 15088
rect 18679 15048 18880 15076
rect 18679 15045 18691 15048
rect 18633 15039 18691 15045
rect 18874 15036 18880 15048
rect 18932 15036 18938 15088
rect 19426 15036 19432 15088
rect 19484 15076 19490 15088
rect 19521 15079 19579 15085
rect 19521 15076 19533 15079
rect 19484 15048 19533 15076
rect 19484 15036 19490 15048
rect 19521 15045 19533 15048
rect 19567 15045 19579 15079
rect 43806 15076 43812 15088
rect 43767 15048 43812 15076
rect 19521 15039 19579 15045
rect 43806 15036 43812 15048
rect 43864 15036 43870 15088
rect 17819 14980 17908 15008
rect 17957 15011 18015 15017
rect 17819 14977 17831 14980
rect 17773 14971 17831 14977
rect 17957 14977 17969 15011
rect 18003 15008 18015 15011
rect 18506 15008 18512 15020
rect 18003 14980 18512 15008
rect 18003 14977 18015 14980
rect 17957 14971 18015 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14940 14703 14943
rect 14826 14940 14832 14952
rect 14691 14912 14832 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 14384 14872 14412 14903
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 14918 14872 14924 14884
rect 14384 14844 14924 14872
rect 14918 14832 14924 14844
rect 14976 14872 14982 14884
rect 17512 14872 17540 14971
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 20622 14968 20628 15020
rect 20680 14968 20686 15020
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 22060 14980 22293 15008
rect 22060 14968 22066 14980
rect 22281 14977 22293 14980
rect 22327 15008 22339 15011
rect 24670 15008 24676 15020
rect 22327 14980 24676 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 24670 14968 24676 14980
rect 24728 14968 24734 15020
rect 42794 14968 42800 15020
rect 42852 15008 42858 15020
rect 43625 15011 43683 15017
rect 43625 15008 43637 15011
rect 42852 14980 43637 15008
rect 42852 14968 42858 14980
rect 43625 14977 43637 14980
rect 43671 14977 43683 15011
rect 43625 14971 43683 14977
rect 46842 14968 46848 15020
rect 46900 15008 46906 15020
rect 47765 15011 47823 15017
rect 47765 15008 47777 15011
rect 46900 14980 47777 15008
rect 46900 14968 46906 14980
rect 47765 14977 47777 14980
rect 47811 14977 47823 15011
rect 47765 14971 47823 14977
rect 18598 14900 18604 14952
rect 18656 14940 18662 14952
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 18656 14912 19257 14940
rect 18656 14900 18662 14912
rect 19245 14909 19257 14912
rect 19291 14909 19303 14943
rect 45278 14940 45284 14952
rect 45239 14912 45284 14940
rect 19245 14903 19303 14909
rect 45278 14900 45284 14912
rect 45336 14900 45342 14952
rect 14976 14844 17540 14872
rect 14976 14832 14982 14844
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 18472 14844 19380 14872
rect 18472 14832 18478 14844
rect 19352 14816 19380 14844
rect 18601 14807 18659 14813
rect 18601 14773 18613 14807
rect 18647 14804 18659 14807
rect 19058 14804 19064 14816
rect 18647 14776 19064 14804
rect 18647 14773 18659 14776
rect 18601 14767 18659 14773
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 20993 14807 21051 14813
rect 20993 14804 21005 14807
rect 19392 14776 21005 14804
rect 19392 14764 19398 14776
rect 20993 14773 21005 14776
rect 21039 14773 21051 14807
rect 20993 14767 21051 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 18598 14600 18604 14612
rect 18559 14572 18604 14600
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 19978 14532 19984 14544
rect 18708 14504 19984 14532
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2682 14396 2688 14408
rect 2179 14368 2688 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 16666 14396 16672 14408
rect 2740 14368 6914 14396
rect 16579 14368 16672 14396
rect 2740 14356 2746 14368
rect 6886 14328 6914 14368
rect 16666 14356 16672 14368
rect 16724 14396 16730 14408
rect 17678 14396 17684 14408
rect 16724 14368 17684 14396
rect 16724 14356 16730 14368
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 18601 14399 18659 14405
rect 18601 14365 18613 14399
rect 18647 14396 18659 14399
rect 18708 14396 18736 14504
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 19242 14464 19248 14476
rect 19203 14436 19248 14464
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 20714 14464 20720 14476
rect 20675 14436 20720 14464
rect 20714 14424 20720 14436
rect 20772 14424 20778 14476
rect 21821 14467 21879 14473
rect 21821 14433 21833 14467
rect 21867 14464 21879 14467
rect 22462 14464 22468 14476
rect 21867 14436 22468 14464
rect 21867 14433 21879 14436
rect 21821 14427 21879 14433
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 23382 14464 23388 14476
rect 23343 14436 23388 14464
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 18647 14368 18736 14396
rect 18647 14365 18659 14368
rect 18601 14359 18659 14365
rect 17586 14328 17592 14340
rect 6886 14300 17592 14328
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 16761 14263 16819 14269
rect 16761 14229 16773 14263
rect 16807 14260 16819 14263
rect 16850 14260 16856 14272
rect 16807 14232 16856 14260
rect 16807 14229 16819 14232
rect 16761 14223 16819 14229
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 17788 14260 17816 14359
rect 47118 14356 47124 14408
rect 47176 14396 47182 14408
rect 47213 14399 47271 14405
rect 47213 14396 47225 14399
rect 47176 14368 47225 14396
rect 47176 14356 47182 14368
rect 47213 14365 47225 14368
rect 47259 14365 47271 14399
rect 47213 14359 47271 14365
rect 17865 14331 17923 14337
rect 17865 14297 17877 14331
rect 17911 14328 17923 14331
rect 19429 14331 19487 14337
rect 19429 14328 19441 14331
rect 17911 14300 19441 14328
rect 17911 14297 17923 14300
rect 17865 14291 17923 14297
rect 19429 14297 19441 14300
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 22005 14331 22063 14337
rect 22005 14297 22017 14331
rect 22051 14328 22063 14331
rect 22094 14328 22100 14340
rect 22051 14300 22100 14328
rect 22051 14297 22063 14300
rect 22005 14291 22063 14297
rect 22094 14288 22100 14300
rect 22152 14288 22158 14340
rect 21634 14260 21640 14272
rect 17788 14232 21640 14260
rect 21634 14220 21640 14232
rect 21692 14220 21698 14272
rect 47302 14260 47308 14272
rect 47263 14232 47308 14260
rect 47302 14220 47308 14232
rect 47360 14220 47366 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 17586 14016 17592 14068
rect 17644 14056 17650 14068
rect 20622 14056 20628 14068
rect 17644 14028 20628 14056
rect 17644 14016 17650 14028
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 22152 14028 22197 14056
rect 22152 14016 22158 14028
rect 16850 13988 16856 14000
rect 16811 13960 16856 13988
rect 16850 13948 16856 13960
rect 16908 13948 16914 14000
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16356 13892 16681 13920
rect 16356 13880 16362 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 19058 13880 19064 13932
rect 19116 13920 19122 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19116 13892 19441 13920
rect 19116 13880 19122 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21692 13892 22017 13920
rect 21692 13880 21698 13892
rect 22005 13889 22017 13892
rect 22051 13920 22063 13923
rect 30466 13920 30472 13932
rect 22051 13892 30472 13920
rect 22051 13889 22063 13892
rect 22005 13883 22063 13889
rect 30466 13880 30472 13892
rect 30524 13880 30530 13932
rect 18506 13852 18512 13864
rect 18467 13824 18512 13852
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 19610 13852 19616 13864
rect 19571 13824 19616 13852
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 21358 13852 21364 13864
rect 21315 13824 21364 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 15746 13784 15752 13796
rect 3476 13756 15752 13784
rect 3476 13744 3482 13756
rect 15746 13744 15752 13756
rect 15804 13744 15810 13796
rect 16298 13744 16304 13796
rect 16356 13784 16362 13796
rect 18414 13784 18420 13796
rect 16356 13756 18420 13784
rect 16356 13744 16362 13756
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 47762 13716 47768 13728
rect 47723 13688 47768 13716
rect 47762 13676 47768 13688
rect 47820 13676 47826 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 19337 13515 19395 13521
rect 14884 13484 16804 13512
rect 14884 13472 14890 13484
rect 16776 13385 16804 13484
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19610 13512 19616 13524
rect 19383 13484 19616 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 46293 13379 46351 13385
rect 46293 13345 46305 13379
rect 46339 13376 46351 13379
rect 47762 13376 47768 13388
rect 46339 13348 47768 13376
rect 46339 13345 46351 13348
rect 46293 13339 46351 13345
rect 47762 13336 47768 13348
rect 47820 13336 47826 13388
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 15657 13271 15715 13277
rect 15672 13172 15700 13271
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 17736 13280 19257 13308
rect 17736 13268 17742 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 15749 13243 15807 13249
rect 15749 13209 15761 13243
rect 15795 13240 15807 13243
rect 16485 13243 16543 13249
rect 16485 13240 16497 13243
rect 15795 13212 16497 13240
rect 15795 13209 15807 13212
rect 15749 13203 15807 13209
rect 16485 13209 16497 13212
rect 16531 13209 16543 13243
rect 16485 13203 16543 13209
rect 46477 13243 46535 13249
rect 46477 13209 46489 13243
rect 46523 13240 46535 13243
rect 47302 13240 47308 13252
rect 46523 13212 47308 13240
rect 46523 13209 46535 13212
rect 46477 13203 46535 13209
rect 47302 13200 47308 13212
rect 47360 13200 47366 13252
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 17218 13172 17224 13184
rect 15672 13144 17224 13172
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 22370 12900 22376 12912
rect 21836 12872 22376 12900
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 21836 12841 21864 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 22002 12764 22008 12776
rect 21963 12736 22008 12764
rect 22002 12724 22008 12736
rect 22060 12724 22066 12776
rect 22281 12767 22339 12773
rect 22281 12733 22293 12767
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 3602 12656 3608 12708
rect 3660 12696 3666 12708
rect 22296 12696 22324 12727
rect 3660 12668 22324 12696
rect 3660 12656 3666 12668
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 32030 12628 32036 12640
rect 1627 12600 32036 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 32030 12588 32036 12600
rect 32088 12588 32094 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 21729 12427 21787 12433
rect 21729 12393 21741 12427
rect 21775 12424 21787 12427
rect 22002 12424 22008 12436
rect 21775 12396 22008 12424
rect 21775 12393 21787 12396
rect 21729 12387 21787 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 21637 12223 21695 12229
rect 21637 12220 21649 12223
rect 17276 12192 21649 12220
rect 17276 12180 17282 12192
rect 21637 12189 21649 12192
rect 21683 12189 21695 12223
rect 21637 12183 21695 12189
rect 45922 12180 45928 12232
rect 45980 12220 45986 12232
rect 46753 12223 46811 12229
rect 46753 12220 46765 12223
rect 45980 12192 46765 12220
rect 45980 12180 45986 12192
rect 46753 12189 46765 12192
rect 46799 12189 46811 12223
rect 46753 12183 46811 12189
rect 46474 12044 46480 12096
rect 46532 12084 46538 12096
rect 46845 12087 46903 12093
rect 46845 12084 46857 12087
rect 46532 12056 46857 12084
rect 46532 12044 46538 12056
rect 46845 12053 46857 12056
rect 46891 12053 46903 12087
rect 46845 12047 46903 12053
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 46474 11200 46480 11212
rect 46435 11172 46480 11200
rect 46474 11160 46480 11172
rect 46532 11160 46538 11212
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 12434 10996 12440 11008
rect 3016 10968 12440 10996
rect 3016 10956 3022 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 47394 10616 47400 10668
rect 47452 10656 47458 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 47452 10628 47593 10656
rect 47452 10616 47458 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 47029 10455 47087 10461
rect 47029 10452 47041 10455
rect 46348 10424 47041 10452
rect 46348 10412 46354 10424
rect 47029 10421 47041 10424
rect 47075 10421 47087 10455
rect 47670 10452 47676 10464
rect 47631 10424 47676 10452
rect 47029 10415 47087 10421
rect 47670 10412 47676 10424
rect 47728 10412 47734 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 46477 10115 46535 10121
rect 46477 10081 46489 10115
rect 46523 10112 46535 10115
rect 47670 10112 47676 10124
rect 46523 10084 47676 10112
rect 46523 10081 46535 10084
rect 46477 10075 46535 10081
rect 47670 10072 47676 10084
rect 47728 10072 47734 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 47854 9568 47860 9580
rect 47815 9540 47860 9568
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 47946 9392 47952 9444
rect 48004 9432 48010 9444
rect 48041 9435 48099 9441
rect 48041 9432 48053 9435
rect 48004 9404 48053 9432
rect 48004 9392 48010 9404
rect 48041 9401 48053 9404
rect 48087 9401 48099 9435
rect 48041 9395 48099 9401
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47762 8888 47768 8900
rect 47723 8860 47768 8888
rect 47762 8848 47768 8860
rect 47820 8848 47826 8900
rect 29914 8780 29920 8832
rect 29972 8820 29978 8832
rect 47857 8823 47915 8829
rect 47857 8820 47869 8823
rect 29972 8792 47869 8820
rect 29972 8780 29978 8792
rect 47857 8789 47869 8792
rect 47903 8789 47915 8823
rect 47857 8783 47915 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 46842 8440 46848 8492
rect 46900 8480 46906 8492
rect 48133 8483 48191 8489
rect 48133 8480 48145 8483
rect 46900 8452 48145 8480
rect 46900 8440 46906 8452
rect 48133 8449 48145 8452
rect 48179 8449 48191 8483
rect 48133 8443 48191 8449
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 46842 8276 46848 8288
rect 18564 8248 46848 8276
rect 18564 8236 18570 8248
rect 46842 8236 46848 8248
rect 46900 8236 46906 8288
rect 47118 8236 47124 8288
rect 47176 8276 47182 8288
rect 47949 8279 48007 8285
rect 47949 8276 47961 8279
rect 47176 8248 47961 8276
rect 47176 8236 47182 8248
rect 47949 8245 47961 8248
rect 47995 8245 48007 8279
rect 47949 8239 48007 8245
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 20714 8072 20720 8084
rect 3568 8044 20720 8072
rect 3568 8032 3574 8044
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 46768 7976 47440 8004
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 20162 7936 20168 7948
rect 19392 7908 20168 7936
rect 19392 7896 19398 7908
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 45557 7939 45615 7945
rect 45557 7905 45569 7939
rect 45603 7936 45615 7939
rect 45646 7936 45652 7948
rect 45603 7908 45652 7936
rect 45603 7905 45615 7908
rect 45557 7899 45615 7905
rect 45646 7896 45652 7908
rect 45704 7896 45710 7948
rect 20162 7760 20168 7812
rect 20220 7800 20226 7812
rect 20438 7800 20444 7812
rect 20220 7772 20444 7800
rect 20220 7760 20226 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 45649 7803 45707 7809
rect 45649 7769 45661 7803
rect 45695 7800 45707 7803
rect 46198 7800 46204 7812
rect 45695 7772 46204 7800
rect 45695 7769 45707 7772
rect 45649 7763 45707 7769
rect 46198 7760 46204 7772
rect 46256 7760 46262 7812
rect 46566 7800 46572 7812
rect 46479 7772 46572 7800
rect 46566 7760 46572 7772
rect 46624 7800 46630 7812
rect 46768 7800 46796 7976
rect 47118 7936 47124 7948
rect 47079 7908 47124 7936
rect 47118 7896 47124 7908
rect 47176 7896 47182 7948
rect 47412 7945 47440 7976
rect 47397 7939 47455 7945
rect 47397 7905 47409 7939
rect 47443 7905 47455 7939
rect 47397 7899 47455 7905
rect 46624 7772 46796 7800
rect 47213 7803 47271 7809
rect 46624 7760 46630 7772
rect 47213 7769 47225 7803
rect 47259 7800 47271 7803
rect 47578 7800 47584 7812
rect 47259 7772 47584 7800
rect 47259 7769 47271 7772
rect 47213 7763 47271 7769
rect 47578 7760 47584 7772
rect 47636 7760 47642 7812
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 47578 7528 47584 7540
rect 47539 7500 47584 7528
rect 47578 7488 47584 7500
rect 47636 7488 47642 7540
rect 46198 7352 46204 7404
rect 46256 7392 46262 7404
rect 46293 7395 46351 7401
rect 46293 7392 46305 7395
rect 46256 7364 46305 7392
rect 46256 7352 46262 7364
rect 46293 7361 46305 7364
rect 46339 7361 46351 7395
rect 47765 7395 47823 7401
rect 47765 7392 47777 7395
rect 46293 7355 46351 7361
rect 46768 7364 47777 7392
rect 46768 7333 46796 7364
rect 47765 7361 47777 7364
rect 47811 7361 47823 7395
rect 47765 7355 47823 7361
rect 46753 7327 46811 7333
rect 46753 7293 46765 7327
rect 46799 7293 46811 7327
rect 46753 7287 46811 7293
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 2096 7228 45554 7256
rect 2096 7216 2102 7228
rect 45526 7188 45554 7228
rect 46017 7191 46075 7197
rect 46017 7188 46029 7191
rect 45526 7160 46029 7188
rect 46017 7157 46029 7160
rect 46063 7188 46075 7191
rect 46385 7191 46443 7197
rect 46385 7188 46397 7191
rect 46063 7160 46397 7188
rect 46063 7157 46075 7160
rect 46017 7151 46075 7157
rect 46385 7157 46397 7160
rect 46431 7157 46443 7191
rect 46385 7151 46443 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 23382 6848 23388 6860
rect 3384 6820 23388 6848
rect 3384 6808 3390 6820
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 38657 6851 38715 6857
rect 38657 6817 38669 6851
rect 38703 6848 38715 6851
rect 39390 6848 39396 6860
rect 38703 6820 39396 6848
rect 38703 6817 38715 6820
rect 38657 6811 38715 6817
rect 39390 6808 39396 6820
rect 39448 6808 39454 6860
rect 47302 6848 47308 6860
rect 47263 6820 47308 6848
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 47210 6740 47216 6792
rect 47268 6780 47274 6792
rect 47581 6783 47639 6789
rect 47581 6780 47593 6783
rect 47268 6752 47593 6780
rect 47268 6740 47274 6752
rect 47581 6749 47593 6752
rect 47627 6749 47639 6783
rect 47581 6743 47639 6749
rect 37645 6715 37703 6721
rect 37645 6681 37657 6715
rect 37691 6681 37703 6715
rect 37645 6675 37703 6681
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 37277 6647 37335 6653
rect 37277 6644 37289 6647
rect 6696 6616 37289 6644
rect 6696 6604 6702 6616
rect 37277 6613 37289 6616
rect 37323 6644 37335 6647
rect 37660 6644 37688 6675
rect 37734 6672 37740 6724
rect 37792 6712 37798 6724
rect 37792 6684 37837 6712
rect 37792 6672 37798 6684
rect 37323 6616 37688 6644
rect 37323 6613 37335 6616
rect 37277 6607 37335 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 37553 6443 37611 6449
rect 37553 6409 37565 6443
rect 37599 6440 37611 6443
rect 37734 6440 37740 6452
rect 37599 6412 37740 6440
rect 37599 6409 37611 6412
rect 37553 6403 37611 6409
rect 37734 6400 37740 6412
rect 37792 6400 37798 6452
rect 43990 6400 43996 6452
rect 44048 6440 44054 6452
rect 48041 6443 48099 6449
rect 48041 6440 48053 6443
rect 44048 6412 48053 6440
rect 44048 6400 44054 6412
rect 48041 6409 48053 6412
rect 48087 6409 48099 6443
rect 48041 6403 48099 6409
rect 38470 6372 38476 6384
rect 38431 6344 38476 6372
rect 38470 6332 38476 6344
rect 38528 6332 38534 6384
rect 39390 6372 39396 6384
rect 39351 6344 39396 6372
rect 39390 6332 39396 6344
rect 39448 6332 39454 6384
rect 37734 6304 37740 6316
rect 37695 6276 37740 6304
rect 37734 6264 37740 6276
rect 37792 6264 37798 6316
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 38378 6236 38384 6248
rect 38339 6208 38384 6236
rect 38378 6196 38384 6208
rect 38436 6236 38442 6248
rect 39206 6236 39212 6248
rect 38436 6208 39212 6236
rect 38436 6196 38442 6208
rect 39206 6196 39212 6208
rect 39264 6196 39270 6248
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 37734 5352 37740 5364
rect 37695 5324 37740 5352
rect 37734 5312 37740 5324
rect 37792 5312 37798 5364
rect 37277 5219 37335 5225
rect 37277 5185 37289 5219
rect 37323 5216 37335 5219
rect 38470 5216 38476 5228
rect 37323 5188 38476 5216
rect 37323 5185 37335 5188
rect 37277 5179 37335 5185
rect 38470 5176 38476 5188
rect 38528 5176 38534 5228
rect 39666 5216 39672 5228
rect 39627 5188 39672 5216
rect 39666 5176 39672 5188
rect 39724 5176 39730 5228
rect 47857 5219 47915 5225
rect 47857 5185 47869 5219
rect 47903 5216 47915 5219
rect 47946 5216 47952 5228
rect 47903 5188 47952 5216
rect 47903 5185 47915 5188
rect 47857 5179 47915 5185
rect 47946 5176 47952 5188
rect 48004 5176 48010 5228
rect 26602 5040 26608 5092
rect 26660 5080 26666 5092
rect 48041 5083 48099 5089
rect 48041 5080 48053 5083
rect 26660 5052 48053 5080
rect 26660 5040 26666 5052
rect 48041 5049 48053 5052
rect 48087 5049 48099 5083
rect 48041 5043 48099 5049
rect 37366 5012 37372 5024
rect 37327 4984 37372 5012
rect 37366 4972 37372 4984
rect 37424 4972 37430 5024
rect 39114 4972 39120 5024
rect 39172 5012 39178 5024
rect 39761 5015 39819 5021
rect 39761 5012 39773 5015
rect 39172 4984 39773 5012
rect 39172 4972 39178 4984
rect 39761 4981 39773 4984
rect 39807 4981 39819 5015
rect 39761 4975 39819 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 20070 4700 20076 4752
rect 20128 4740 20134 4752
rect 26234 4740 26240 4752
rect 20128 4712 26240 4740
rect 20128 4700 20134 4712
rect 26234 4700 26240 4712
rect 26292 4700 26298 4752
rect 46290 4700 46296 4752
rect 46348 4740 46354 4752
rect 46348 4712 47624 4740
rect 46348 4700 46354 4712
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 41877 4675 41935 4681
rect 41877 4672 41889 4675
rect 4028 4644 41889 4672
rect 4028 4632 4034 4644
rect 41877 4641 41889 4644
rect 41923 4672 41935 4675
rect 42337 4675 42395 4681
rect 42337 4672 42349 4675
rect 41923 4644 42349 4672
rect 41923 4641 41935 4644
rect 41877 4635 41935 4641
rect 42337 4641 42349 4644
rect 42383 4641 42395 4675
rect 43254 4672 43260 4684
rect 43215 4644 43260 4672
rect 42337 4635 42395 4641
rect 43254 4632 43260 4644
rect 43312 4632 43318 4684
rect 47486 4672 47492 4684
rect 46676 4644 47492 4672
rect 14458 4604 14464 4616
rect 14419 4576 14464 4604
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4604 15255 4607
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15243 4576 15761 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4604 15899 4607
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 15887 4576 16405 4604
rect 15887 4573 15899 4576
rect 15841 4567 15899 4573
rect 16393 4573 16405 4576
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4604 16543 4607
rect 17037 4607 17095 4613
rect 17037 4604 17049 4607
rect 16531 4576 17049 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 17037 4573 17049 4576
rect 17083 4573 17095 4607
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 17037 4567 17095 4573
rect 15120 4536 15148 4567
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4604 21051 4607
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 21039 4576 21557 4604
rect 21039 4573 21051 4576
rect 20993 4567 21051 4573
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 39114 4604 39120 4616
rect 39075 4576 39120 4604
rect 21545 4567 21603 4573
rect 39114 4564 39120 4576
rect 39172 4564 39178 4616
rect 39853 4607 39911 4613
rect 39853 4573 39865 4607
rect 39899 4604 39911 4607
rect 40126 4604 40132 4616
rect 39899 4576 40132 4604
rect 39899 4573 39911 4576
rect 39853 4567 39911 4573
rect 40126 4564 40132 4576
rect 40184 4564 40190 4616
rect 40862 4604 40868 4616
rect 40823 4576 40868 4604
rect 40862 4564 40868 4576
rect 40920 4564 40926 4616
rect 46676 4613 46704 4644
rect 47486 4632 47492 4644
rect 47544 4632 47550 4684
rect 47596 4681 47624 4712
rect 47581 4675 47639 4681
rect 47581 4641 47593 4675
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 46661 4607 46719 4613
rect 46661 4573 46673 4607
rect 46707 4573 46719 4607
rect 46661 4567 46719 4573
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47305 4607 47363 4613
rect 47305 4604 47317 4607
rect 46900 4576 47317 4604
rect 46900 4564 46906 4576
rect 47305 4573 47317 4576
rect 47351 4573 47363 4607
rect 47305 4567 47363 4573
rect 15654 4536 15660 4548
rect 15120 4508 15660 4536
rect 15654 4496 15660 4508
rect 15712 4496 15718 4548
rect 26145 4539 26203 4545
rect 26145 4536 26157 4539
rect 26068 4508 26157 4536
rect 14553 4471 14611 4477
rect 14553 4437 14565 4471
rect 14599 4468 14611 4471
rect 15838 4468 15844 4480
rect 14599 4440 15844 4468
rect 14599 4437 14611 4440
rect 14553 4431 14611 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 16666 4428 16672 4480
rect 16724 4468 16730 4480
rect 17129 4471 17187 4477
rect 17129 4468 17141 4471
rect 16724 4440 17141 4468
rect 16724 4428 16730 4440
rect 17129 4437 17141 4440
rect 17175 4437 17187 4471
rect 17129 4431 17187 4437
rect 21637 4471 21695 4477
rect 21637 4437 21649 4471
rect 21683 4468 21695 4471
rect 23382 4468 23388 4480
rect 21683 4440 23388 4468
rect 21683 4437 21695 4440
rect 21637 4431 21695 4437
rect 23382 4428 23388 4440
rect 23440 4428 23446 4480
rect 24854 4428 24860 4480
rect 24912 4468 24918 4480
rect 26068 4468 26096 4508
rect 26145 4505 26157 4508
rect 26191 4505 26203 4539
rect 26145 4499 26203 4505
rect 26234 4496 26240 4548
rect 26292 4536 26298 4548
rect 26970 4536 26976 4548
rect 26292 4508 26976 4536
rect 26292 4496 26298 4508
rect 26970 4496 26976 4508
rect 27028 4496 27034 4548
rect 27157 4539 27215 4545
rect 27157 4505 27169 4539
rect 27203 4536 27215 4539
rect 27706 4536 27712 4548
rect 27203 4508 27712 4536
rect 27203 4505 27215 4508
rect 27157 4499 27215 4505
rect 27706 4496 27712 4508
rect 27764 4496 27770 4548
rect 39942 4496 39948 4548
rect 40000 4536 40006 4548
rect 40037 4539 40095 4545
rect 40037 4536 40049 4539
rect 40000 4508 40049 4536
rect 40000 4496 40006 4508
rect 40037 4505 40049 4508
rect 40083 4505 40095 4539
rect 40037 4499 40095 4505
rect 42429 4539 42487 4545
rect 42429 4505 42441 4539
rect 42475 4536 42487 4539
rect 44082 4536 44088 4548
rect 42475 4508 44088 4536
rect 42475 4505 42487 4508
rect 42429 4499 42487 4505
rect 44082 4496 44088 4508
rect 44140 4496 44146 4548
rect 38378 4468 38384 4480
rect 24912 4440 38384 4468
rect 24912 4428 24918 4440
rect 38378 4428 38384 4440
rect 38436 4428 38442 4480
rect 38654 4428 38660 4480
rect 38712 4468 38718 4480
rect 39209 4471 39267 4477
rect 39209 4468 39221 4471
rect 38712 4440 39221 4468
rect 38712 4428 38718 4440
rect 39209 4437 39221 4440
rect 39255 4437 39267 4471
rect 40218 4468 40224 4480
rect 40179 4440 40224 4468
rect 39209 4431 39267 4437
rect 40218 4428 40224 4440
rect 40276 4428 40282 4480
rect 40681 4471 40739 4477
rect 40681 4437 40693 4471
rect 40727 4468 40739 4471
rect 41046 4468 41052 4480
rect 40727 4440 41052 4468
rect 40727 4437 40739 4440
rect 40681 4431 40739 4437
rect 41046 4428 41052 4440
rect 41104 4428 41110 4480
rect 46474 4428 46480 4480
rect 46532 4468 46538 4480
rect 46753 4471 46811 4477
rect 46753 4468 46765 4471
rect 46532 4440 46765 4468
rect 46532 4428 46538 4440
rect 46753 4437 46765 4440
rect 46799 4437 46811 4471
rect 46753 4431 46811 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 14458 4224 14464 4276
rect 14516 4264 14522 4276
rect 14553 4267 14611 4273
rect 14553 4264 14565 4267
rect 14516 4236 14565 4264
rect 14516 4224 14522 4236
rect 14553 4233 14565 4236
rect 14599 4233 14611 4267
rect 14553 4227 14611 4233
rect 20898 4224 20904 4276
rect 20956 4264 20962 4276
rect 21177 4267 21235 4273
rect 21177 4264 21189 4267
rect 20956 4236 21189 4264
rect 20956 4224 20962 4236
rect 21177 4233 21189 4236
rect 21223 4233 21235 4267
rect 21177 4227 21235 4233
rect 39482 4224 39488 4276
rect 39540 4264 39546 4276
rect 46845 4267 46903 4273
rect 46845 4264 46857 4267
rect 39540 4236 46857 4264
rect 39540 4224 39546 4236
rect 46845 4233 46857 4236
rect 46891 4233 46903 4267
rect 46845 4227 46903 4233
rect 40218 4196 40224 4208
rect 21928 4168 22140 4196
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 7190 4060 7196 4072
rect 7151 4032 7196 4060
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4060 7435 4063
rect 8110 4060 8116 4072
rect 7423 4032 8116 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 10612 4060 10640 4091
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 13412 4100 13553 4128
rect 13412 4088 13418 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 13872 4100 14473 4128
rect 13872 4088 13878 4100
rect 14461 4097 14473 4100
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4128 17003 4131
rect 17494 4128 17500 4140
rect 16991 4100 17500 4128
rect 16991 4097 17003 4100
rect 16945 4091 17003 4097
rect 15746 4060 15752 4072
rect 8260 4032 8305 4060
rect 10612 4032 15752 4060
rect 8260 4020 8266 4032
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 15856 4060 15884 4091
rect 17494 4088 17500 4100
rect 17552 4088 17558 4140
rect 17957 4131 18015 4137
rect 17957 4097 17969 4131
rect 18003 4128 18015 4131
rect 18230 4128 18236 4140
rect 18003 4100 18236 4128
rect 18003 4097 18015 4100
rect 17957 4091 18015 4097
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 19484 4100 19533 4128
rect 19484 4088 19490 4100
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 20438 4128 20444 4140
rect 20399 4100 20444 4128
rect 19521 4091 19579 4097
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 21085 4131 21143 4137
rect 21085 4128 21097 4131
rect 20864 4100 21097 4128
rect 20864 4088 20870 4100
rect 21085 4097 21097 4100
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 21174 4088 21180 4140
rect 21232 4128 21238 4140
rect 21928 4128 21956 4168
rect 21232 4100 21956 4128
rect 22005 4131 22063 4137
rect 21232 4088 21238 4100
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 17218 4060 17224 4072
rect 15856 4032 17224 4060
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 17310 4020 17316 4072
rect 17368 4060 17374 4072
rect 20162 4060 20168 4072
rect 17368 4032 20168 4060
rect 17368 4020 17374 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 22020 4060 22048 4091
rect 20680 4032 22048 4060
rect 22112 4060 22140 4168
rect 39408 4168 40224 4196
rect 22278 4088 22284 4140
rect 22336 4128 22342 4140
rect 28718 4128 28724 4140
rect 22336 4100 28724 4128
rect 22336 4088 22342 4100
rect 28718 4088 28724 4100
rect 28776 4088 28782 4140
rect 38381 4131 38439 4137
rect 38381 4097 38393 4131
rect 38427 4128 38439 4131
rect 38654 4128 38660 4140
rect 38427 4100 38660 4128
rect 38427 4097 38439 4100
rect 38381 4091 38439 4097
rect 38654 4088 38660 4100
rect 38712 4088 38718 4140
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4128 39267 4131
rect 39408 4128 39436 4168
rect 40218 4156 40224 4168
rect 40276 4156 40282 4208
rect 42886 4196 42892 4208
rect 42847 4168 42892 4196
rect 42886 4156 42892 4168
rect 42944 4156 42950 4208
rect 43254 4156 43260 4208
rect 43312 4196 43318 4208
rect 43809 4199 43867 4205
rect 43809 4196 43821 4199
rect 43312 4168 43821 4196
rect 43312 4156 43318 4168
rect 43809 4165 43821 4168
rect 43855 4165 43867 4199
rect 43809 4159 43867 4165
rect 46382 4156 46388 4208
rect 46440 4196 46446 4208
rect 46569 4199 46627 4205
rect 46569 4196 46581 4199
rect 46440 4168 46581 4196
rect 46440 4156 46446 4168
rect 46569 4165 46581 4168
rect 46615 4165 46627 4199
rect 46569 4159 46627 4165
rect 46658 4156 46664 4208
rect 46716 4196 46722 4208
rect 47765 4199 47823 4205
rect 47765 4196 47777 4199
rect 46716 4168 47777 4196
rect 46716 4156 46722 4168
rect 47765 4165 47777 4168
rect 47811 4165 47823 4199
rect 47765 4159 47823 4165
rect 39669 4131 39727 4137
rect 39669 4128 39681 4131
rect 39255 4100 39436 4128
rect 39500 4100 39681 4128
rect 39255 4097 39267 4100
rect 39209 4091 39267 4097
rect 32214 4060 32220 4072
rect 22112 4032 32220 4060
rect 20680 4020 20686 4032
rect 32214 4020 32220 4032
rect 32272 4020 32278 4072
rect 38473 4063 38531 4069
rect 38473 4029 38485 4063
rect 38519 4060 38531 4063
rect 39500 4060 39528 4100
rect 39669 4097 39681 4100
rect 39715 4097 39727 4131
rect 44450 4128 44456 4140
rect 44411 4100 44456 4128
rect 39669 4091 39727 4097
rect 44450 4088 44456 4100
rect 44508 4088 44514 4140
rect 38519 4032 39528 4060
rect 38519 4029 38531 4032
rect 38473 4023 38531 4029
rect 39574 4020 39580 4072
rect 39632 4060 39638 4072
rect 39853 4063 39911 4069
rect 39853 4060 39865 4063
rect 39632 4032 39865 4060
rect 39632 4020 39638 4032
rect 39853 4029 39865 4032
rect 39899 4029 39911 4063
rect 41414 4060 41420 4072
rect 41375 4032 41420 4060
rect 39853 4023 39911 4029
rect 41414 4020 41420 4032
rect 41472 4020 41478 4072
rect 41506 4020 41512 4072
rect 41564 4060 41570 4072
rect 42797 4063 42855 4069
rect 42797 4060 42809 4063
rect 41564 4032 42809 4060
rect 41564 4020 41570 4032
rect 42797 4029 42809 4032
rect 42843 4060 42855 4063
rect 45646 4060 45652 4072
rect 42843 4032 45652 4060
rect 42843 4029 42855 4032
rect 42797 4023 42855 4029
rect 45646 4020 45652 4032
rect 45704 4020 45710 4072
rect 21726 3992 21732 4004
rect 6886 3964 21732 3992
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1636 3896 2145 3924
rect 1636 3884 1642 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2866 3924 2872 3936
rect 2827 3896 2872 3924
rect 2133 3887 2191 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 6886 3924 6914 3964
rect 21726 3952 21732 3964
rect 21784 3952 21790 4004
rect 21910 3952 21916 4004
rect 21968 3992 21974 4004
rect 22833 3995 22891 4001
rect 22833 3992 22845 3995
rect 21968 3964 22845 3992
rect 21968 3952 21974 3964
rect 22833 3961 22845 3964
rect 22879 3961 22891 3995
rect 39482 3992 39488 4004
rect 22833 3955 22891 3961
rect 26206 3964 39488 3992
rect 10686 3924 10692 3936
rect 3844 3896 6914 3924
rect 10647 3896 10692 3924
rect 3844 3884 3850 3896
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 13633 3927 13691 3933
rect 13633 3893 13645 3927
rect 13679 3924 13691 3927
rect 13722 3924 13728 3936
rect 13679 3896 13728 3924
rect 13679 3893 13691 3896
rect 13633 3887 13691 3893
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15160 3896 15301 3924
rect 15160 3884 15166 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15930 3924 15936 3936
rect 15891 3896 15936 3924
rect 15289 3887 15347 3893
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 17037 3927 17095 3933
rect 17037 3893 17049 3927
rect 17083 3924 17095 3927
rect 17954 3924 17960 3936
rect 17083 3896 17960 3924
rect 17083 3893 17095 3896
rect 17037 3887 17095 3893
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 19242 3924 19248 3936
rect 18095 3896 19248 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3924 19671 3927
rect 20070 3924 20076 3936
rect 19659 3896 20076 3924
rect 19659 3893 19671 3896
rect 19613 3887 19671 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20533 3927 20591 3933
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 20714 3924 20720 3936
rect 20579 3896 20720 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 22094 3924 22100 3936
rect 22055 3896 22100 3924
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 26206 3924 26234 3964
rect 39482 3952 39488 3964
rect 39540 3952 39546 4004
rect 22244 3896 26234 3924
rect 22244 3884 22250 3896
rect 29454 3884 29460 3936
rect 29512 3924 29518 3936
rect 36538 3924 36544 3936
rect 29512 3896 36544 3924
rect 29512 3884 29518 3896
rect 36538 3884 36544 3896
rect 36596 3884 36602 3936
rect 39025 3927 39083 3933
rect 39025 3893 39037 3927
rect 39071 3924 39083 3927
rect 39574 3924 39580 3936
rect 39071 3896 39580 3924
rect 39071 3893 39083 3896
rect 39025 3887 39083 3893
rect 39574 3884 39580 3896
rect 39632 3884 39638 3936
rect 44082 3884 44088 3936
rect 44140 3924 44146 3936
rect 44269 3927 44327 3933
rect 44269 3924 44281 3927
rect 44140 3896 44281 3924
rect 44140 3884 44146 3896
rect 44269 3893 44281 3896
rect 44315 3893 44327 3927
rect 44269 3887 44327 3893
rect 46017 3927 46075 3933
rect 46017 3893 46029 3927
rect 46063 3924 46075 3927
rect 46290 3924 46296 3936
rect 46063 3896 46296 3924
rect 46063 3893 46075 3896
rect 46017 3887 46075 3893
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 47854 3924 47860 3936
rect 47815 3896 47860 3924
rect 47854 3884 47860 3896
rect 47912 3884 47918 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 8110 3720 8116 3732
rect 8071 3692 8116 3720
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 17494 3720 17500 3732
rect 10520 3692 16252 3720
rect 17455 3692 17500 3720
rect 10410 3652 10416 3664
rect 8036 3624 10416 3652
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 1820 3556 3985 3584
rect 1820 3544 1826 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 3973 3547 4031 3553
rect 2682 3516 2688 3528
rect 2643 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 8036 3525 8064 3624
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 10520 3584 10548 3692
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 13044 3624 16068 3652
rect 13044 3612 13050 3624
rect 10686 3584 10692 3596
rect 9876 3556 10548 3584
rect 10647 3556 10692 3584
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6604 3488 6745 3516
rect 6604 3476 6610 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1360 3420 1869 3448
rect 1360 3408 1366 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 1857 3411 1915 3417
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 7282 3448 7288 3460
rect 2271 3420 7288 3448
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 7392 3448 7420 3479
rect 9122 3476 9128 3528
rect 9180 3516 9186 3528
rect 9876 3525 9904 3556
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 15102 3584 15108 3596
rect 13280 3556 14412 3584
rect 15063 3556 15108 3584
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9180 3488 9321 3516
rect 9180 3476 9186 3488
rect 9309 3485 9321 3488
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9861 3519 9919 3525
rect 9861 3485 9873 3519
rect 9907 3485 9919 3519
rect 10502 3516 10508 3528
rect 10463 3488 10508 3516
rect 9861 3479 9919 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 13170 3448 13176 3460
rect 7392 3420 13176 3448
rect 13170 3408 13176 3420
rect 13228 3408 13234 3460
rect 2774 3380 2780 3392
rect 2735 3352 2780 3380
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 6788 3352 7481 3380
rect 6788 3340 6794 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9953 3383 10011 3389
rect 9953 3380 9965 3383
rect 9364 3352 9965 3380
rect 9364 3340 9370 3352
rect 9953 3349 9965 3352
rect 9999 3349 10011 3383
rect 9953 3343 10011 3349
rect 10410 3340 10416 3392
rect 10468 3380 10474 3392
rect 13280 3380 13308 3556
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 13372 3448 13400 3479
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13596 3488 14289 3516
rect 13596 3476 13602 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 13998 3448 14004 3460
rect 13372 3420 14004 3448
rect 13998 3408 14004 3420
rect 14056 3408 14062 3460
rect 14384 3448 14412 3556
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15930 3584 15936 3596
rect 15335 3556 15936 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16040 3593 16068 3624
rect 16025 3587 16083 3593
rect 16025 3553 16037 3587
rect 16071 3553 16083 3587
rect 16224 3584 16252 3692
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 19334 3720 19340 3732
rect 18380 3692 19340 3720
rect 18380 3680 18386 3692
rect 19334 3680 19340 3692
rect 19392 3720 19398 3732
rect 21726 3720 21732 3732
rect 19392 3692 21312 3720
rect 21687 3692 21732 3720
rect 19392 3680 19398 3692
rect 16298 3612 16304 3664
rect 16356 3652 16362 3664
rect 21174 3652 21180 3664
rect 16356 3624 21180 3652
rect 16356 3612 16362 3624
rect 21174 3612 21180 3624
rect 21232 3612 21238 3664
rect 19978 3584 19984 3596
rect 16224 3556 19984 3584
rect 16025 3547 16083 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 21284 3584 21312 3692
rect 21726 3680 21732 3692
rect 21784 3720 21790 3732
rect 24854 3720 24860 3732
rect 21784 3692 24860 3720
rect 21784 3680 21790 3692
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 39209 3723 39267 3729
rect 39209 3689 39221 3723
rect 39255 3720 39267 3723
rect 39666 3720 39672 3732
rect 39255 3692 39672 3720
rect 39255 3689 39267 3692
rect 39209 3683 39267 3689
rect 39666 3680 39672 3692
rect 39724 3680 39730 3732
rect 40126 3720 40132 3732
rect 40087 3692 40132 3720
rect 40126 3680 40132 3692
rect 40184 3680 40190 3732
rect 40405 3723 40463 3729
rect 40405 3689 40417 3723
rect 40451 3720 40463 3723
rect 40862 3720 40868 3732
rect 40451 3692 40868 3720
rect 40451 3689 40463 3692
rect 40405 3683 40463 3689
rect 40862 3680 40868 3692
rect 40920 3680 40926 3732
rect 21358 3612 21364 3664
rect 21416 3652 21422 3664
rect 30926 3652 30932 3664
rect 21416 3624 30932 3652
rect 21416 3612 21422 3624
rect 30926 3612 30932 3624
rect 30984 3612 30990 3664
rect 32950 3612 32956 3664
rect 33008 3652 33014 3664
rect 33873 3655 33931 3661
rect 33873 3652 33885 3655
rect 33008 3624 33885 3652
rect 33008 3612 33014 3624
rect 33873 3621 33885 3624
rect 33919 3621 33931 3655
rect 33873 3615 33931 3621
rect 36538 3612 36544 3664
rect 36596 3652 36602 3664
rect 47854 3652 47860 3664
rect 36596 3624 47860 3652
rect 36596 3612 36602 3624
rect 47854 3612 47860 3624
rect 47912 3612 47918 3664
rect 23569 3587 23627 3593
rect 23569 3584 23581 3587
rect 21284 3556 22416 3584
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17405 3519 17463 3525
rect 17405 3516 17417 3519
rect 16816 3488 17417 3516
rect 16816 3476 16822 3488
rect 17405 3485 17417 3488
rect 17451 3485 17463 3519
rect 17405 3479 17463 3485
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 18012 3488 18061 3516
rect 18012 3476 18018 3488
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 19242 3516 19248 3528
rect 19203 3488 19248 3516
rect 18049 3479 18107 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19889 3519 19947 3525
rect 19889 3516 19901 3519
rect 19392 3488 19901 3516
rect 19392 3476 19398 3488
rect 19889 3485 19901 3488
rect 19935 3485 19947 3519
rect 19889 3479 19947 3485
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20220 3488 20545 3516
rect 20220 3476 20226 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 22005 3519 22063 3525
rect 22005 3485 22017 3519
rect 22051 3516 22063 3519
rect 22186 3516 22192 3528
rect 22051 3488 22192 3516
rect 22051 3485 22063 3488
rect 22005 3479 22063 3485
rect 22186 3476 22192 3488
rect 22244 3476 22250 3528
rect 16942 3448 16948 3460
rect 14384 3420 16948 3448
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 22278 3448 22284 3460
rect 17052 3420 22284 3448
rect 10468 3352 13308 3380
rect 10468 3340 10474 3352
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 13449 3383 13507 3389
rect 13449 3380 13461 3383
rect 13412 3352 13461 3380
rect 13412 3340 13418 3352
rect 13449 3349 13461 3352
rect 13495 3349 13507 3383
rect 13449 3343 13507 3349
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 17052 3380 17080 3420
rect 22278 3408 22284 3420
rect 22336 3408 22342 3460
rect 22388 3448 22416 3556
rect 22848 3556 23581 3584
rect 22848 3525 22876 3556
rect 23569 3553 23581 3556
rect 23615 3553 23627 3587
rect 23569 3547 23627 3553
rect 23658 3544 23664 3596
rect 23716 3584 23722 3596
rect 26145 3587 26203 3593
rect 26145 3584 26157 3587
rect 23716 3556 26157 3584
rect 23716 3544 23722 3556
rect 26145 3553 26157 3556
rect 26191 3553 26203 3587
rect 26145 3547 26203 3553
rect 27157 3587 27215 3593
rect 27157 3553 27169 3587
rect 27203 3584 27215 3587
rect 27706 3584 27712 3596
rect 27203 3556 27712 3584
rect 27203 3553 27215 3556
rect 27157 3547 27215 3553
rect 27706 3544 27712 3556
rect 27764 3544 27770 3596
rect 32766 3544 32772 3596
rect 32824 3584 32830 3596
rect 36446 3584 36452 3596
rect 32824 3556 36452 3584
rect 32824 3544 32830 3556
rect 36446 3544 36452 3556
rect 36504 3544 36510 3596
rect 41046 3584 41052 3596
rect 41007 3556 41052 3584
rect 41046 3544 41052 3556
rect 41104 3544 41110 3596
rect 41414 3584 41420 3596
rect 41375 3556 41420 3584
rect 41414 3544 41420 3556
rect 41472 3544 41478 3596
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23382 3476 23388 3528
rect 23440 3516 23446 3528
rect 23477 3519 23535 3525
rect 23477 3516 23489 3519
rect 23440 3488 23489 3516
rect 23440 3476 23446 3488
rect 23477 3485 23489 3488
rect 23523 3485 23535 3519
rect 24765 3519 24823 3525
rect 24765 3516 24777 3519
rect 23477 3479 23535 3485
rect 23584 3488 24777 3516
rect 23584 3448 23612 3488
rect 24765 3485 24777 3488
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 25593 3519 25651 3525
rect 25593 3485 25605 3519
rect 25639 3485 25651 3519
rect 25593 3479 25651 3485
rect 33045 3519 33103 3525
rect 33045 3485 33057 3519
rect 33091 3516 33103 3519
rect 39114 3516 39120 3528
rect 33091 3488 34008 3516
rect 39075 3488 39120 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 22388 3420 23612 3448
rect 24578 3408 24584 3460
rect 24636 3448 24642 3460
rect 25608 3448 25636 3479
rect 24636 3420 25636 3448
rect 24636 3408 24642 3420
rect 26234 3408 26240 3460
rect 26292 3448 26298 3460
rect 33980 3448 34008 3488
rect 39114 3476 39120 3488
rect 39172 3476 39178 3528
rect 39853 3519 39911 3525
rect 39853 3485 39865 3519
rect 39899 3516 39911 3519
rect 39942 3516 39948 3528
rect 39899 3488 39948 3516
rect 39899 3485 39911 3488
rect 39853 3479 39911 3485
rect 39942 3476 39948 3488
rect 40000 3476 40006 3528
rect 40221 3519 40279 3525
rect 40221 3485 40233 3519
rect 40267 3516 40279 3519
rect 40586 3516 40592 3528
rect 40267 3488 40592 3516
rect 40267 3485 40279 3488
rect 40221 3479 40279 3485
rect 40586 3476 40592 3488
rect 40644 3476 40650 3528
rect 40862 3516 40868 3528
rect 40823 3488 40868 3516
rect 40862 3476 40868 3488
rect 40920 3476 40926 3528
rect 43165 3519 43223 3525
rect 43165 3516 43177 3519
rect 42260 3488 43177 3516
rect 35710 3448 35716 3460
rect 26292 3420 26337 3448
rect 33980 3420 35716 3448
rect 26292 3408 26298 3420
rect 35710 3408 35716 3420
rect 35768 3448 35774 3460
rect 42260 3448 42288 3488
rect 43165 3485 43177 3488
rect 43211 3485 43223 3519
rect 43165 3479 43223 3485
rect 43993 3519 44051 3525
rect 43993 3485 44005 3519
rect 44039 3485 44051 3519
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 43993 3479 44051 3485
rect 35768 3420 42288 3448
rect 35768 3408 35774 3420
rect 42794 3408 42800 3460
rect 42852 3448 42858 3460
rect 44008 3448 44036 3479
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 42852 3420 44036 3448
rect 45664 3448 45692 3479
rect 47394 3448 47400 3460
rect 45664 3420 47400 3448
rect 42852 3408 42858 3420
rect 47394 3408 47400 3420
rect 47452 3408 47458 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 13688 3352 17080 3380
rect 13688 3340 13694 3352
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 18141 3383 18199 3389
rect 18141 3380 18153 3383
rect 17644 3352 18153 3380
rect 17644 3340 17650 3352
rect 18141 3349 18153 3352
rect 18187 3349 18199 3383
rect 18141 3343 18199 3349
rect 18782 3340 18788 3392
rect 18840 3380 18846 3392
rect 19337 3383 19395 3389
rect 19337 3380 19349 3383
rect 18840 3352 19349 3380
rect 18840 3340 18846 3352
rect 19337 3349 19349 3352
rect 19383 3349 19395 3383
rect 19978 3380 19984 3392
rect 19939 3352 19984 3380
rect 19337 3343 19395 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 20254 3340 20260 3392
rect 20312 3380 20318 3392
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 20312 3352 20637 3380
rect 20312 3340 20318 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 20625 3343 20683 3349
rect 24762 3340 24768 3392
rect 24820 3380 24826 3392
rect 24857 3383 24915 3389
rect 24857 3380 24869 3383
rect 24820 3352 24869 3380
rect 24820 3340 24826 3352
rect 24857 3349 24869 3352
rect 24903 3349 24915 3383
rect 33134 3380 33140 3392
rect 33095 3352 33140 3380
rect 24857 3343 24915 3349
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 34422 3340 34428 3392
rect 34480 3380 34486 3392
rect 42426 3380 42432 3392
rect 34480 3352 42432 3380
rect 34480 3340 34486 3352
rect 42426 3340 42432 3352
rect 42484 3340 42490 3392
rect 42978 3340 42984 3392
rect 43036 3380 43042 3392
rect 43257 3383 43315 3389
rect 43257 3380 43269 3383
rect 43036 3352 43269 3380
rect 43036 3340 43042 3352
rect 43257 3349 43269 3352
rect 43303 3349 43315 3383
rect 43257 3343 43315 3349
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 16758 3176 16764 3188
rect 3936 3148 16620 3176
rect 16719 3148 16764 3176
rect 3936 3136 3942 3148
rect 1949 3111 2007 3117
rect 1949 3077 1961 3111
rect 1995 3108 2007 3111
rect 2774 3108 2780 3120
rect 1995 3080 2780 3108
rect 1995 3077 2007 3080
rect 1949 3071 2007 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 6730 3108 6736 3120
rect 6691 3080 6736 3108
rect 6730 3068 6736 3080
rect 6788 3068 6794 3120
rect 7282 3068 7288 3120
rect 7340 3108 7346 3120
rect 9306 3108 9312 3120
rect 7340 3080 8432 3108
rect 9267 3080 9312 3108
rect 7340 3068 7346 3080
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 7009 2975 7067 2981
rect 7009 2972 7021 2975
rect 6512 2944 7021 2972
rect 6512 2932 6518 2944
rect 7009 2941 7021 2944
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 8404 2904 8432 3080
rect 9306 3068 9312 3080
rect 9364 3068 9370 3120
rect 10520 3080 13400 3108
rect 9122 3040 9128 3052
rect 9083 3012 9128 3040
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 9088 2944 9597 2972
rect 9088 2932 9094 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 10520 2904 10548 3080
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 12400 2944 12633 2972
rect 12400 2932 12406 2944
rect 12621 2941 12633 2944
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 7800 2876 8340 2904
rect 8404 2876 10548 2904
rect 12728 2904 12756 3003
rect 13372 2972 13400 3080
rect 13446 3068 13452 3120
rect 13504 3108 13510 3120
rect 13504 3080 15608 3108
rect 13504 3068 13510 3080
rect 13538 3040 13544 3052
rect 13499 3012 13544 3040
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13446 2972 13452 2984
rect 13372 2944 13452 2972
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 14182 2972 14188 2984
rect 13780 2944 13825 2972
rect 14143 2944 14188 2972
rect 13780 2932 13786 2944
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 15580 2972 15608 3080
rect 15654 3068 15660 3120
rect 15712 3108 15718 3120
rect 15933 3111 15991 3117
rect 15933 3108 15945 3111
rect 15712 3080 15945 3108
rect 15712 3068 15718 3080
rect 15933 3077 15945 3080
rect 15979 3077 15991 3111
rect 16592 3108 16620 3148
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 18230 3176 18236 3188
rect 16868 3148 17724 3176
rect 18191 3148 18236 3176
rect 16868 3108 16896 3148
rect 17586 3108 17592 3120
rect 16592 3080 16896 3108
rect 17420 3080 17592 3108
rect 15933 3071 15991 3077
rect 15838 3040 15844 3052
rect 15799 3012 15844 3040
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17420 3049 17448 3080
rect 17586 3068 17592 3080
rect 17644 3068 17650 3120
rect 17696 3108 17724 3148
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18877 3179 18935 3185
rect 18877 3145 18889 3179
rect 18923 3176 18935 3179
rect 19334 3176 19340 3188
rect 18923 3148 19340 3176
rect 18923 3145 18935 3148
rect 18877 3139 18935 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 19521 3179 19579 3185
rect 19521 3176 19533 3179
rect 19484 3148 19533 3176
rect 19484 3136 19490 3148
rect 19521 3145 19533 3148
rect 19567 3145 19579 3179
rect 20162 3176 20168 3188
rect 20123 3148 20168 3176
rect 19521 3139 19579 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 20806 3176 20812 3188
rect 20767 3148 20812 3176
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 32766 3176 32772 3188
rect 20956 3148 32772 3176
rect 20956 3136 20962 3148
rect 32766 3136 32772 3148
rect 32824 3136 32830 3188
rect 32968 3148 35572 3176
rect 32968 3108 32996 3148
rect 33134 3108 33140 3120
rect 17696 3080 32996 3108
rect 33095 3080 33140 3108
rect 33134 3068 33140 3080
rect 33192 3068 33198 3120
rect 35544 3108 35572 3148
rect 39114 3136 39120 3188
rect 39172 3176 39178 3188
rect 39853 3179 39911 3185
rect 39853 3176 39865 3179
rect 39172 3148 39865 3176
rect 39172 3136 39178 3148
rect 39853 3145 39865 3148
rect 39899 3145 39911 3179
rect 39853 3139 39911 3145
rect 40862 3136 40868 3188
rect 40920 3176 40926 3188
rect 41049 3179 41107 3185
rect 41049 3176 41061 3179
rect 40920 3148 41061 3176
rect 40920 3136 40926 3148
rect 41049 3145 41061 3148
rect 41095 3145 41107 3179
rect 45094 3176 45100 3188
rect 41049 3139 41107 3145
rect 41386 3148 45100 3176
rect 41386 3108 41414 3148
rect 45094 3136 45100 3148
rect 45152 3136 45158 3188
rect 47670 3136 47676 3188
rect 47728 3176 47734 3188
rect 47857 3179 47915 3185
rect 47857 3176 47869 3179
rect 47728 3148 47869 3176
rect 47728 3136 47734 3148
rect 47857 3145 47869 3148
rect 47903 3145 47915 3179
rect 47857 3139 47915 3145
rect 42978 3108 42984 3120
rect 35544 3080 41414 3108
rect 42939 3080 42984 3108
rect 42978 3068 42984 3080
rect 43036 3068 43042 3120
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 17543 3012 18153 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 18141 3009 18153 3012
rect 18187 3009 18199 3043
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18141 3003 18199 3009
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 19978 3040 19984 3052
rect 19475 3012 19984 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 20070 3000 20076 3052
rect 20128 3040 20134 3052
rect 20714 3040 20720 3052
rect 20128 3012 20173 3040
rect 20675 3012 20720 3040
rect 20128 3000 20134 3012
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 21910 3040 21916 3052
rect 21871 3012 21916 3040
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 24578 3040 24584 3052
rect 24539 3012 24584 3040
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 26970 3040 26976 3052
rect 26931 3012 26976 3040
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 27062 3000 27068 3052
rect 27120 3040 27126 3052
rect 27985 3043 28043 3049
rect 27985 3040 27997 3043
rect 27120 3012 27997 3040
rect 27120 3000 27126 3012
rect 27985 3009 27997 3012
rect 28031 3009 28043 3043
rect 27985 3003 28043 3009
rect 28169 3043 28227 3049
rect 28169 3009 28181 3043
rect 28215 3040 28227 3043
rect 29362 3040 29368 3052
rect 28215 3012 29368 3040
rect 28215 3009 28227 3012
rect 28169 3003 28227 3009
rect 29362 3000 29368 3012
rect 29420 3000 29426 3052
rect 32950 3040 32956 3052
rect 32911 3012 32956 3040
rect 32950 3000 32956 3012
rect 33008 3000 33014 3052
rect 39114 3000 39120 3052
rect 39172 3040 39178 3052
rect 39393 3043 39451 3049
rect 39393 3040 39405 3043
rect 39172 3012 39405 3040
rect 39172 3000 39178 3012
rect 39393 3009 39405 3012
rect 39439 3040 39451 3043
rect 39942 3040 39948 3052
rect 39439 3012 39948 3040
rect 39439 3009 39451 3012
rect 39393 3003 39451 3009
rect 39942 3000 39948 3012
rect 40000 3000 40006 3052
rect 41506 3040 41512 3052
rect 40512 3012 41512 3040
rect 18322 2972 18328 2984
rect 15580 2944 18328 2972
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 21266 2972 21272 2984
rect 19392 2944 21272 2972
rect 19392 2932 19398 2944
rect 21266 2932 21272 2944
rect 21324 2932 21330 2984
rect 22094 2972 22100 2984
rect 22055 2944 22100 2972
rect 22094 2932 22100 2944
rect 22152 2932 22158 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 24762 2972 24768 2984
rect 24723 2944 24768 2972
rect 24762 2932 24768 2944
rect 24820 2932 24826 2984
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 26418 2932 26424 2984
rect 26476 2972 26482 2984
rect 27433 2975 27491 2981
rect 27433 2972 27445 2975
rect 26476 2944 27445 2972
rect 26476 2932 26482 2944
rect 27433 2941 27445 2944
rect 27479 2941 27491 2975
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 27433 2935 27491 2941
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 39206 2972 39212 2984
rect 39167 2944 39212 2972
rect 39206 2932 39212 2944
rect 39264 2972 39270 2984
rect 40405 2975 40463 2981
rect 40405 2972 40417 2975
rect 39264 2944 40417 2972
rect 39264 2932 39270 2944
rect 40405 2941 40417 2944
rect 40451 2972 40463 2975
rect 40512 2972 40540 3012
rect 41506 3000 41512 3012
rect 41564 3000 41570 3052
rect 42794 3040 42800 3052
rect 42755 3012 42800 3040
rect 42794 3000 42800 3012
rect 42852 3000 42858 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3040 47823 3043
rect 48314 3040 48320 3052
rect 47811 3012 48320 3040
rect 47811 3009 47823 3012
rect 47765 3003 47823 3009
rect 48314 3000 48320 3012
rect 48372 3000 48378 3052
rect 40451 2944 40540 2972
rect 40451 2941 40463 2944
rect 40405 2935 40463 2941
rect 40586 2932 40592 2984
rect 40644 2972 40650 2984
rect 41690 2972 41696 2984
rect 40644 2944 41696 2972
rect 40644 2932 40650 2944
rect 41690 2932 41696 2944
rect 41748 2932 41754 2984
rect 43162 2932 43168 2984
rect 43220 2972 43226 2984
rect 43257 2975 43315 2981
rect 43257 2972 43269 2975
rect 43220 2944 43269 2972
rect 43220 2932 43226 2944
rect 43257 2941 43269 2944
rect 43303 2941 43315 2975
rect 43257 2935 43315 2941
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 41414 2904 41420 2916
rect 12728 2876 41420 2904
rect 7800 2864 7806 2876
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 8202 2836 8208 2848
rect 7156 2808 8208 2836
rect 7156 2796 7162 2808
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8312 2836 8340 2876
rect 41414 2864 41420 2876
rect 41472 2864 41478 2916
rect 12986 2836 12992 2848
rect 8312 2808 12992 2836
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 14090 2836 14096 2848
rect 13127 2808 14096 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 20898 2836 20904 2848
rect 15804 2808 20904 2836
rect 15804 2796 15810 2808
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 27249 2839 27307 2845
rect 27249 2805 27261 2839
rect 27295 2836 27307 2839
rect 33134 2836 33140 2848
rect 27295 2808 33140 2836
rect 27295 2805 27307 2808
rect 27249 2799 27307 2805
rect 33134 2796 33140 2808
rect 33192 2796 33198 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 2866 2592 2872 2644
rect 2924 2592 2930 2644
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 4614 2632 4620 2644
rect 4571 2604 4620 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7248 2604 7481 2632
rect 7248 2592 7254 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 7469 2595 7527 2601
rect 10502 2592 10508 2644
rect 10560 2632 10566 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10560 2604 10793 2632
rect 10560 2592 10566 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 10781 2595 10839 2601
rect 13449 2635 13507 2641
rect 13449 2601 13461 2635
rect 13495 2632 13507 2635
rect 13814 2632 13820 2644
rect 13495 2604 13820 2632
rect 13495 2601 13507 2604
rect 13449 2595 13507 2601
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 14056 2604 14197 2632
rect 14056 2592 14062 2604
rect 14185 2601 14197 2604
rect 14231 2601 14243 2635
rect 14185 2595 14243 2601
rect 19889 2635 19947 2641
rect 19889 2601 19901 2635
rect 19935 2632 19947 2635
rect 20438 2632 20444 2644
rect 19935 2604 20444 2632
rect 19935 2601 19947 2604
rect 19889 2595 19947 2601
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 20530 2592 20536 2644
rect 20588 2632 20594 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20588 2604 20913 2632
rect 20588 2592 20594 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 20901 2595 20959 2601
rect 22186 2592 22192 2644
rect 22244 2632 22250 2644
rect 22373 2635 22431 2641
rect 22373 2632 22385 2635
rect 22244 2604 22385 2632
rect 22244 2592 22250 2604
rect 22373 2601 22385 2604
rect 22419 2601 22431 2635
rect 22373 2595 22431 2601
rect 23385 2635 23443 2641
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 23658 2632 23664 2644
rect 23431 2604 23664 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 24949 2635 25007 2641
rect 24949 2601 24961 2635
rect 24995 2632 25007 2635
rect 25038 2632 25044 2644
rect 24995 2604 25044 2632
rect 24995 2601 25007 2604
rect 24949 2595 25007 2601
rect 25038 2592 25044 2604
rect 25096 2592 25102 2644
rect 26234 2592 26240 2644
rect 26292 2632 26298 2644
rect 28629 2635 28687 2641
rect 26292 2604 26337 2632
rect 26292 2592 26298 2604
rect 28629 2601 28641 2635
rect 28675 2632 28687 2635
rect 28810 2632 28816 2644
rect 28675 2604 28816 2632
rect 28675 2601 28687 2604
rect 28629 2595 28687 2601
rect 28810 2592 28816 2604
rect 28868 2592 28874 2644
rect 33134 2592 33140 2644
rect 33192 2632 33198 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 33192 2604 35541 2632
rect 33192 2592 33198 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 36354 2632 36360 2644
rect 36315 2604 36360 2632
rect 35529 2595 35587 2601
rect 36354 2592 36360 2604
rect 36412 2592 36418 2644
rect 39114 2632 39120 2644
rect 39075 2604 39120 2632
rect 39114 2592 39120 2604
rect 39172 2592 39178 2644
rect 41690 2632 41696 2644
rect 41651 2604 41696 2632
rect 41690 2592 41696 2604
rect 41748 2592 41754 2644
rect 42518 2632 42524 2644
rect 42479 2604 42524 2632
rect 42518 2592 42524 2604
rect 42576 2592 42582 2644
rect 42889 2635 42947 2641
rect 42889 2601 42901 2635
rect 42935 2632 42947 2635
rect 44450 2632 44456 2644
rect 42935 2604 44456 2632
rect 42935 2601 42947 2604
rect 42889 2595 42947 2601
rect 44450 2592 44456 2604
rect 44508 2592 44514 2644
rect 2884 2564 2912 2592
rect 1412 2536 2912 2564
rect 15841 2567 15899 2573
rect 1412 2505 1440 2536
rect 15841 2533 15853 2567
rect 15887 2564 15899 2567
rect 37366 2564 37372 2576
rect 15887 2536 37372 2564
rect 15887 2533 15899 2536
rect 15841 2527 15899 2533
rect 37366 2524 37372 2536
rect 37424 2524 37430 2576
rect 41233 2567 41291 2573
rect 41233 2533 41245 2567
rect 41279 2564 41291 2567
rect 43070 2564 43076 2576
rect 41279 2536 43076 2564
rect 41279 2533 41291 2536
rect 41233 2527 41291 2533
rect 43070 2524 43076 2536
rect 43128 2524 43134 2576
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2866 2496 2872 2508
rect 2827 2468 2872 2496
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2496 9735 2499
rect 27246 2496 27252 2508
rect 9723 2468 27108 2496
rect 27207 2468 27252 2496
rect 9723 2465 9735 2468
rect 9677 2459 9735 2465
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 5445 2391 5503 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 19797 2431 19855 2437
rect 19797 2397 19809 2431
rect 19843 2428 19855 2431
rect 20254 2428 20260 2440
rect 19843 2400 20260 2428
rect 19843 2397 19855 2400
rect 19797 2391 19855 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23256 2400 23581 2428
rect 23256 2388 23262 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 26418 2428 26424 2440
rect 26379 2400 26424 2428
rect 23569 2391 23627 2397
rect 26418 2388 26424 2400
rect 26476 2388 26482 2440
rect 26510 2388 26516 2440
rect 26568 2428 26574 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26568 2400 26985 2428
rect 26568 2388 26574 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 27080 2428 27108 2468
rect 27246 2456 27252 2468
rect 27304 2456 27310 2508
rect 34238 2456 34244 2508
rect 34296 2496 34302 2508
rect 38381 2499 38439 2505
rect 38381 2496 38393 2499
rect 34296 2468 38393 2496
rect 34296 2456 34302 2468
rect 38381 2465 38393 2468
rect 38427 2465 38439 2499
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 38381 2459 38439 2465
rect 38488 2468 40509 2496
rect 27890 2428 27896 2440
rect 27080 2400 27896 2428
rect 26973 2391 27031 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 38488 2428 38516 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 42886 2496 42892 2508
rect 40497 2459 40555 2465
rect 42444 2468 42892 2496
rect 35713 2391 35771 2397
rect 35866 2400 38516 2428
rect 39301 2431 39359 2437
rect 4249 2363 4307 2369
rect 4249 2329 4261 2363
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 4264 2292 4292 2323
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8444 2332 9413 2360
rect 8444 2320 8450 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 15528 2332 15669 2360
rect 15528 2320 15534 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 21910 2320 21916 2372
rect 21968 2360 21974 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21968 2332 22293 2360
rect 21968 2320 21974 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22281 2323 22339 2329
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24544 2332 24869 2360
rect 24544 2320 24550 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 32398 2320 32404 2372
rect 32456 2360 32462 2372
rect 35866 2360 35894 2400
rect 39301 2397 39313 2431
rect 39347 2428 39359 2431
rect 39942 2428 39948 2440
rect 39347 2400 39948 2428
rect 39347 2397 39359 2400
rect 39301 2391 39359 2397
rect 39942 2388 39948 2400
rect 40000 2388 40006 2440
rect 41230 2388 41236 2440
rect 41288 2428 41294 2440
rect 42444 2437 42472 2468
rect 42886 2456 42892 2468
rect 42944 2496 42950 2508
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 42944 2468 46489 2496
rect 42944 2456 42950 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 46477 2459 46535 2465
rect 46750 2456 46756 2508
rect 46808 2496 46814 2508
rect 47857 2499 47915 2505
rect 47857 2496 47869 2499
rect 46808 2468 47869 2496
rect 46808 2456 46814 2468
rect 47857 2465 47869 2468
rect 47903 2465 47915 2499
rect 47857 2459 47915 2465
rect 41877 2431 41935 2437
rect 41877 2428 41889 2431
rect 41288 2400 41889 2428
rect 41288 2388 41294 2400
rect 41877 2397 41889 2400
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 42429 2431 42487 2437
rect 42429 2397 42441 2431
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 46201 2431 46259 2437
rect 46201 2397 46213 2431
rect 46247 2428 46259 2431
rect 47026 2428 47032 2440
rect 46247 2400 47032 2428
rect 46247 2397 46259 2400
rect 46201 2391 46259 2397
rect 32456 2332 35894 2360
rect 32456 2320 32462 2332
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 38197 2363 38255 2369
rect 38197 2360 38209 2363
rect 38068 2332 38209 2360
rect 38068 2320 38074 2332
rect 38197 2329 38209 2332
rect 38243 2329 38255 2363
rect 38197 2323 38255 2329
rect 39390 2320 39396 2372
rect 39448 2360 39454 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39448 2332 40325 2360
rect 39448 2320 39454 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41049 2363 41107 2369
rect 41049 2360 41061 2363
rect 40644 2332 41061 2360
rect 40644 2320 40650 2332
rect 41049 2329 41061 2332
rect 41095 2329 41107 2363
rect 43916 2360 43944 2391
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 47673 2431 47731 2437
rect 47673 2397 47685 2431
rect 47719 2428 47731 2431
rect 48038 2428 48044 2440
rect 47719 2400 48044 2428
rect 47719 2397 47731 2400
rect 47673 2391 47731 2397
rect 48038 2388 48044 2400
rect 48096 2388 48102 2440
rect 41049 2323 41107 2329
rect 41156 2332 43944 2360
rect 45373 2363 45431 2369
rect 2648 2264 4292 2292
rect 5261 2295 5319 2301
rect 2648 2252 2654 2264
rect 5261 2261 5273 2295
rect 5307 2292 5319 2295
rect 12342 2292 12348 2304
rect 5307 2264 12348 2292
rect 5307 2261 5319 2264
rect 5261 2255 5319 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 25222 2292 25228 2304
rect 16899 2264 25228 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 25222 2252 25228 2264
rect 25280 2252 25286 2304
rect 29730 2292 29736 2304
rect 29691 2264 29736 2292
rect 29730 2252 29736 2264
rect 29788 2252 29794 2304
rect 38470 2252 38476 2304
rect 38528 2292 38534 2304
rect 41156 2292 41184 2332
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46750 2360 46756 2372
rect 45419 2332 46756 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46750 2320 46756 2332
rect 46808 2320 46814 2372
rect 38528 2264 41184 2292
rect 38528 2252 38534 2264
rect 41782 2252 41788 2304
rect 41840 2292 41846 2304
rect 45465 2295 45523 2301
rect 45465 2292 45477 2295
rect 41840 2264 45477 2292
rect 41840 2252 41846 2264
rect 45465 2261 45477 2264
rect 45511 2261 45523 2295
rect 45465 2255 45523 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 29730 1980 29736 2032
rect 29788 2020 29794 2032
rect 42518 2020 42524 2032
rect 29788 1992 42524 2020
rect 29788 1980 29794 1992
rect 42518 1980 42524 1992
rect 42576 1980 42582 2032
rect 32858 1912 32864 1964
rect 32916 1952 32922 1964
rect 41782 1952 41788 1964
rect 32916 1924 41788 1952
rect 32916 1912 32922 1924
rect 41782 1912 41788 1924
rect 41840 1912 41846 1964
<< via1 >>
rect 44824 47404 44876 47456
rect 45468 47404 45520 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 22284 47132 22336 47184
rect 30196 47132 30248 47184
rect 40132 47132 40184 47184
rect 48044 47132 48096 47184
rect 30748 47107 30800 47116
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 43168 47107 43220 47116
rect 43168 47073 43177 47107
rect 43177 47073 43211 47107
rect 43211 47073 43220 47107
rect 43168 47064 43220 47073
rect 48320 47064 48372 47116
rect 1952 46996 2004 47048
rect 3240 46996 3292 47048
rect 4712 47039 4764 47048
rect 4712 47005 4721 47039
rect 4721 47005 4755 47039
rect 4755 47005 4764 47039
rect 4712 46996 4764 47005
rect 5816 46996 5868 47048
rect 7288 47039 7340 47048
rect 7288 47005 7297 47039
rect 7297 47005 7331 47039
rect 7331 47005 7340 47039
rect 7288 46996 7340 47005
rect 9036 46996 9088 47048
rect 11612 46996 11664 47048
rect 12256 46996 12308 47048
rect 12624 47039 12676 47048
rect 12624 47005 12633 47039
rect 12633 47005 12667 47039
rect 12667 47005 12676 47039
rect 12624 46996 12676 47005
rect 13820 46996 13872 47048
rect 16488 46996 16540 47048
rect 20720 47039 20772 47048
rect 20720 47005 20729 47039
rect 20729 47005 20763 47039
rect 20763 47005 20772 47039
rect 20720 46996 20772 47005
rect 4068 46971 4120 46980
rect 2596 46860 2648 46912
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 4988 46971 5040 46980
rect 4988 46937 4997 46971
rect 4997 46937 5031 46971
rect 5031 46937 5040 46971
rect 4988 46928 5040 46937
rect 6644 46971 6696 46980
rect 6644 46937 6653 46971
rect 6653 46937 6687 46971
rect 6687 46937 6696 46971
rect 6644 46928 6696 46937
rect 9496 46928 9548 46980
rect 11796 46928 11848 46980
rect 2872 46903 2924 46912
rect 2872 46869 2881 46903
rect 2881 46869 2915 46903
rect 2915 46869 2924 46903
rect 7472 46903 7524 46912
rect 2872 46860 2924 46869
rect 7472 46869 7481 46903
rect 7481 46869 7515 46903
rect 7515 46869 7524 46903
rect 7472 46860 7524 46869
rect 12900 46860 12952 46912
rect 15568 46928 15620 46980
rect 20076 46971 20128 46980
rect 14648 46903 14700 46912
rect 14648 46869 14657 46903
rect 14657 46869 14691 46903
rect 14691 46869 14700 46903
rect 14648 46860 14700 46869
rect 18696 46860 18748 46912
rect 20076 46937 20085 46971
rect 20085 46937 20119 46971
rect 20119 46937 20128 46971
rect 20076 46928 20128 46937
rect 19984 46860 20036 46912
rect 28448 46996 28500 47048
rect 29644 46996 29696 47048
rect 31576 46996 31628 47048
rect 38108 46996 38160 47048
rect 40224 46996 40276 47048
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 28356 46928 28408 46980
rect 42800 46971 42852 46980
rect 21824 46903 21876 46912
rect 21824 46869 21833 46903
rect 21833 46869 21867 46903
rect 21867 46869 21876 46903
rect 21824 46860 21876 46869
rect 39304 46860 39356 46912
rect 42800 46937 42809 46971
rect 42809 46937 42843 46971
rect 42843 46937 42852 46971
rect 42800 46928 42852 46937
rect 45100 46928 45152 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1860 46631 1912 46640
rect 1860 46597 1869 46631
rect 1869 46597 1903 46631
rect 1903 46597 1912 46631
rect 1860 46588 1912 46597
rect 3884 46588 3936 46640
rect 32036 46588 32088 46640
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 47952 46563 48004 46572
rect 47952 46529 47961 46563
rect 47961 46529 47995 46563
rect 47995 46529 48004 46563
rect 47952 46520 48004 46529
rect 3976 46495 4028 46504
rect 3976 46461 3985 46495
rect 3985 46461 4019 46495
rect 4019 46461 4028 46495
rect 3976 46452 4028 46461
rect 5172 46452 5224 46504
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 14280 46452 14332 46461
rect 19616 46495 19668 46504
rect 19616 46461 19625 46495
rect 19625 46461 19659 46495
rect 19659 46461 19668 46495
rect 19616 46452 19668 46461
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 27620 46452 27672 46504
rect 2044 46427 2096 46436
rect 2044 46393 2053 46427
rect 2053 46393 2087 46427
rect 2087 46393 2096 46427
rect 2044 46384 2096 46393
rect 25780 46384 25832 46436
rect 32312 46452 32364 46504
rect 38292 46495 38344 46504
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 45192 46495 45244 46504
rect 42524 46384 42576 46436
rect 45192 46461 45201 46495
rect 45201 46461 45235 46495
rect 45235 46461 45244 46495
rect 45192 46452 45244 46461
rect 45560 46452 45612 46504
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 1400 46316 1452 46368
rect 10416 46316 10468 46368
rect 25228 46316 25280 46368
rect 41328 46316 41380 46368
rect 41420 46316 41472 46368
rect 47216 46316 47268 46368
rect 47308 46316 47360 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3976 46112 4028 46164
rect 5172 46155 5224 46164
rect 5172 46121 5181 46155
rect 5181 46121 5215 46155
rect 5215 46121 5224 46155
rect 5172 46112 5224 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 19616 46112 19668 46164
rect 27620 46155 27672 46164
rect 1400 46019 1452 46028
rect 1400 45985 1409 46019
rect 1409 45985 1443 46019
rect 1443 45985 1452 46019
rect 1400 45976 1452 45985
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 10416 46019 10468 46028
rect 10416 45985 10425 46019
rect 10425 45985 10459 46019
rect 10459 45985 10468 46019
rect 10416 45976 10468 45985
rect 10968 45976 11020 46028
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 18420 45908 18472 45960
rect 18604 45908 18656 45960
rect 20720 46044 20772 46096
rect 26240 46019 26292 46028
rect 26240 45985 26249 46019
rect 26249 45985 26283 46019
rect 26283 45985 26292 46019
rect 26240 45976 26292 45985
rect 21640 45908 21692 45960
rect 25228 45951 25280 45960
rect 25228 45917 25237 45951
rect 25237 45917 25271 45951
rect 25271 45917 25280 45951
rect 25228 45908 25280 45917
rect 2228 45840 2280 45892
rect 10600 45883 10652 45892
rect 10600 45849 10609 45883
rect 10609 45849 10643 45883
rect 10643 45849 10652 45883
rect 10600 45840 10652 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 25504 45840 25556 45892
rect 27620 46121 27629 46155
rect 27629 46121 27663 46155
rect 27663 46121 27672 46155
rect 27620 46112 27672 46121
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 42432 46112 42484 46164
rect 41420 46044 41472 46096
rect 41328 46019 41380 46028
rect 41328 45985 41337 46019
rect 41337 45985 41371 46019
rect 41371 45985 41380 46019
rect 41328 45976 41380 45985
rect 41880 46019 41932 46028
rect 41880 45985 41889 46019
rect 41889 45985 41923 46019
rect 41923 45985 41932 46019
rect 41880 45976 41932 45985
rect 46480 45976 46532 46028
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 38200 45951 38252 45960
rect 38200 45917 38209 45951
rect 38209 45917 38243 45951
rect 38243 45917 38252 45951
rect 38200 45908 38252 45917
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 41512 45883 41564 45892
rect 25136 45772 25188 45824
rect 26240 45772 26292 45824
rect 41512 45849 41521 45883
rect 41521 45849 41555 45883
rect 41555 45849 41564 45883
rect 41512 45840 41564 45849
rect 44180 45883 44232 45892
rect 44180 45849 44189 45883
rect 44189 45849 44223 45883
rect 44223 45849 44232 45883
rect 44180 45840 44232 45849
rect 47676 45840 47728 45892
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 2228 45611 2280 45620
rect 2228 45577 2237 45611
rect 2237 45577 2271 45611
rect 2271 45577 2280 45611
rect 2228 45568 2280 45577
rect 10600 45611 10652 45620
rect 10600 45577 10609 45611
rect 10609 45577 10643 45611
rect 10643 45577 10652 45611
rect 10600 45568 10652 45577
rect 25412 45568 25464 45620
rect 38200 45568 38252 45620
rect 41512 45568 41564 45620
rect 42616 45568 42668 45620
rect 45744 45568 45796 45620
rect 46572 45543 46624 45552
rect 46572 45509 46581 45543
rect 46581 45509 46615 45543
rect 46615 45509 46624 45543
rect 46572 45500 46624 45509
rect 47676 45543 47728 45552
rect 47676 45509 47685 45543
rect 47685 45509 47719 45543
rect 47719 45509 47728 45543
rect 47676 45500 47728 45509
rect 2320 45432 2372 45484
rect 18512 45432 18564 45484
rect 26056 45475 26108 45484
rect 26056 45441 26065 45475
rect 26065 45441 26099 45475
rect 26099 45441 26108 45475
rect 26056 45432 26108 45441
rect 41328 45475 41380 45484
rect 41328 45441 41337 45475
rect 41337 45441 41371 45475
rect 41371 45441 41380 45475
rect 41328 45432 41380 45441
rect 42432 45475 42484 45484
rect 42432 45441 42441 45475
rect 42441 45441 42475 45475
rect 42475 45441 42484 45475
rect 42432 45432 42484 45441
rect 42892 45432 42944 45484
rect 47216 45432 47268 45484
rect 47492 45432 47544 45484
rect 44456 45364 44508 45416
rect 45376 45407 45428 45416
rect 45376 45373 45385 45407
rect 45385 45373 45419 45407
rect 45419 45373 45428 45407
rect 45376 45364 45428 45373
rect 43260 45228 43312 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 42800 45024 42852 45076
rect 45928 44888 45980 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 38660 44863 38712 44872
rect 38660 44829 38669 44863
rect 38669 44829 38703 44863
rect 38703 44829 38712 44863
rect 38660 44820 38712 44829
rect 42892 44820 42944 44872
rect 45468 44863 45520 44872
rect 38752 44727 38804 44736
rect 38752 44693 38761 44727
rect 38761 44693 38795 44727
rect 38795 44693 38804 44727
rect 38752 44684 38804 44693
rect 45468 44829 45477 44863
rect 45477 44829 45511 44863
rect 45511 44829 45520 44863
rect 45468 44820 45520 44829
rect 46296 44863 46348 44872
rect 46296 44829 46305 44863
rect 46305 44829 46339 44863
rect 46339 44829 46348 44863
rect 46296 44820 46348 44829
rect 45652 44795 45704 44804
rect 45652 44761 45661 44795
rect 45661 44761 45695 44795
rect 45695 44761 45704 44795
rect 45652 44752 45704 44761
rect 47676 44752 47728 44804
rect 47584 44684 47636 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 45560 44480 45612 44532
rect 47676 44523 47728 44532
rect 47676 44489 47685 44523
rect 47685 44489 47719 44523
rect 47719 44489 47728 44523
rect 47676 44480 47728 44489
rect 38752 44455 38804 44464
rect 38752 44421 38761 44455
rect 38761 44421 38795 44455
rect 38795 44421 38804 44455
rect 38752 44412 38804 44421
rect 44456 44387 44508 44396
rect 44456 44353 44465 44387
rect 44465 44353 44499 44387
rect 44499 44353 44508 44387
rect 44456 44344 44508 44353
rect 46296 44412 46348 44464
rect 45744 44344 45796 44396
rect 46204 44387 46256 44396
rect 46204 44353 46213 44387
rect 46213 44353 46247 44387
rect 46247 44353 46256 44387
rect 46204 44344 46256 44353
rect 38568 44319 38620 44328
rect 38568 44285 38577 44319
rect 38577 44285 38611 44319
rect 38611 44285 38620 44319
rect 38568 44276 38620 44285
rect 40040 44319 40092 44328
rect 40040 44285 40049 44319
rect 40049 44285 40083 44319
rect 40083 44285 40092 44319
rect 40040 44276 40092 44285
rect 41328 44276 41380 44328
rect 45100 44208 45152 44260
rect 46940 44183 46992 44192
rect 46940 44149 46949 44183
rect 46949 44149 46983 44183
rect 46983 44149 46992 44183
rect 46940 44140 46992 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 45192 43936 45244 43988
rect 45928 43800 45980 43852
rect 46940 43800 46992 43852
rect 48228 43800 48280 43852
rect 26424 43732 26476 43784
rect 38568 43596 38620 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 45284 43256 45336 43308
rect 46480 43256 46532 43308
rect 1492 43188 1544 43240
rect 47768 43095 47820 43104
rect 47768 43061 47777 43095
rect 47777 43061 47811 43095
rect 47811 43061 47820 43095
rect 47768 43052 47820 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47768 42712 47820 42764
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 47584 42211 47636 42220
rect 47584 42177 47593 42211
rect 47593 42177 47627 42211
rect 47627 42177 47636 42211
rect 47584 42168 47636 42177
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47676 41624 47728 41676
rect 48136 41599 48188 41608
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46480 41216 46532 41268
rect 14096 41080 14148 41132
rect 42432 41080 42484 41132
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 39672 40876 39724 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 1952 40375 2004 40384
rect 1952 40341 1961 40375
rect 1961 40341 1995 40375
rect 1995 40341 2004 40375
rect 1952 40332 2004 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 20168 39516 20220 39568
rect 38660 39516 38712 39568
rect 22652 39448 22704 39500
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 22468 39423 22520 39432
rect 22468 39389 22477 39423
rect 22477 39389 22511 39423
rect 22511 39389 22520 39423
rect 22468 39380 22520 39389
rect 25504 39380 25556 39432
rect 23480 39244 23532 39296
rect 25320 39287 25372 39296
rect 25320 39253 25329 39287
rect 25329 39253 25363 39287
rect 25363 39253 25372 39287
rect 25320 39244 25372 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 25320 39040 25372 39092
rect 20168 38972 20220 39024
rect 20444 38972 20496 39024
rect 21824 38972 21876 39024
rect 19432 38947 19484 38956
rect 19432 38913 19441 38947
rect 19441 38913 19475 38947
rect 19475 38913 19484 38947
rect 19432 38904 19484 38913
rect 22652 38972 22704 39024
rect 22836 38972 22888 39024
rect 22100 38879 22152 38888
rect 22100 38845 22109 38879
rect 22109 38845 22143 38879
rect 22143 38845 22152 38879
rect 22376 38879 22428 38888
rect 22100 38836 22152 38845
rect 22376 38845 22385 38879
rect 22385 38845 22419 38879
rect 22419 38845 22428 38879
rect 22376 38836 22428 38845
rect 25504 38904 25556 38956
rect 47676 38947 47728 38956
rect 47676 38913 47685 38947
rect 47685 38913 47719 38947
rect 47719 38913 47728 38947
rect 47676 38904 47728 38913
rect 24400 38836 24452 38888
rect 47860 38879 47912 38888
rect 47860 38845 47869 38879
rect 47869 38845 47903 38879
rect 47903 38845 47912 38879
rect 47860 38836 47912 38845
rect 20536 38700 20588 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 22376 38496 22428 38548
rect 20168 38428 20220 38480
rect 41328 38496 41380 38548
rect 12624 38360 12676 38412
rect 19432 38335 19484 38344
rect 19432 38301 19441 38335
rect 19441 38301 19475 38335
rect 19475 38301 19484 38335
rect 19432 38292 19484 38301
rect 18512 38267 18564 38276
rect 18512 38233 18521 38267
rect 18521 38233 18555 38267
rect 18555 38233 18564 38267
rect 18512 38224 18564 38233
rect 20168 38224 20220 38276
rect 21364 38267 21416 38276
rect 21364 38233 21373 38267
rect 21373 38233 21407 38267
rect 21407 38233 21416 38267
rect 21364 38224 21416 38233
rect 22100 38360 22152 38412
rect 26976 38360 27028 38412
rect 23480 38292 23532 38344
rect 25964 38292 26016 38344
rect 29184 38292 29236 38344
rect 46940 38292 46992 38344
rect 24584 38224 24636 38276
rect 25412 38224 25464 38276
rect 23664 38199 23716 38208
rect 23664 38165 23673 38199
rect 23673 38165 23707 38199
rect 23707 38165 23716 38199
rect 23664 38156 23716 38165
rect 24492 38156 24544 38208
rect 26148 38199 26200 38208
rect 26148 38165 26157 38199
rect 26157 38165 26191 38199
rect 26191 38165 26200 38199
rect 26148 38156 26200 38165
rect 27988 38199 28040 38208
rect 27988 38165 27997 38199
rect 27997 38165 28031 38199
rect 28031 38165 28040 38199
rect 27988 38156 28040 38165
rect 28264 38156 28316 38208
rect 38200 38156 38252 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 19432 37952 19484 38004
rect 22836 37952 22888 38004
rect 24584 37995 24636 38004
rect 24584 37961 24593 37995
rect 24593 37961 24627 37995
rect 24627 37961 24636 37995
rect 24584 37952 24636 37961
rect 25412 37952 25464 38004
rect 23664 37884 23716 37936
rect 19064 37816 19116 37868
rect 19432 37859 19484 37868
rect 19432 37825 19441 37859
rect 19441 37825 19475 37859
rect 19475 37825 19484 37859
rect 19432 37816 19484 37825
rect 19616 37816 19668 37868
rect 19432 37680 19484 37732
rect 24400 37859 24452 37868
rect 24400 37825 24409 37859
rect 24409 37825 24443 37859
rect 24443 37825 24452 37859
rect 27988 37884 28040 37936
rect 24400 37816 24452 37825
rect 24860 37816 24912 37868
rect 25964 37816 26016 37868
rect 26976 37859 27028 37868
rect 26976 37825 26985 37859
rect 26985 37825 27019 37859
rect 27019 37825 27028 37859
rect 26976 37816 27028 37825
rect 29184 37859 29236 37868
rect 29184 37825 29193 37859
rect 29193 37825 29227 37859
rect 29227 37825 29236 37859
rect 29184 37816 29236 37825
rect 31024 37816 31076 37868
rect 47492 37816 47544 37868
rect 24492 37791 24544 37800
rect 24492 37757 24501 37791
rect 24501 37757 24535 37791
rect 24535 37757 24544 37791
rect 24492 37748 24544 37757
rect 27252 37791 27304 37800
rect 27252 37757 27261 37791
rect 27261 37757 27295 37791
rect 27295 37757 27304 37791
rect 27252 37748 27304 37757
rect 24952 37680 25004 37732
rect 21364 37612 21416 37664
rect 28264 37612 28316 37664
rect 28724 37655 28776 37664
rect 28724 37621 28733 37655
rect 28733 37621 28767 37655
rect 28767 37621 28776 37655
rect 28724 37612 28776 37621
rect 29276 37655 29328 37664
rect 29276 37621 29285 37655
rect 29285 37621 29319 37655
rect 29319 37621 29328 37655
rect 29276 37612 29328 37621
rect 47676 37655 47728 37664
rect 47676 37621 47685 37655
rect 47685 37621 47719 37655
rect 47719 37621 47728 37655
rect 47676 37612 47728 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19616 37451 19668 37460
rect 19616 37417 19625 37451
rect 19625 37417 19659 37451
rect 19659 37417 19668 37451
rect 19616 37408 19668 37417
rect 19984 37408 20036 37460
rect 26148 37408 26200 37460
rect 24400 37340 24452 37392
rect 25780 37340 25832 37392
rect 26976 37272 27028 37324
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 1768 37204 1820 37256
rect 14188 37204 14240 37256
rect 14648 37204 14700 37256
rect 20260 37204 20312 37256
rect 25504 37247 25556 37256
rect 25504 37213 25513 37247
rect 25513 37213 25547 37247
rect 25547 37213 25556 37247
rect 25504 37204 25556 37213
rect 25596 37204 25648 37256
rect 26792 37247 26844 37256
rect 26792 37213 26801 37247
rect 26801 37213 26835 37247
rect 26835 37213 26844 37247
rect 26792 37204 26844 37213
rect 31024 37204 31076 37256
rect 25872 37136 25924 37188
rect 21916 37111 21968 37120
rect 21916 37077 21925 37111
rect 21925 37077 21959 37111
rect 21959 37077 21968 37111
rect 21916 37068 21968 37077
rect 24860 37068 24912 37120
rect 25412 37068 25464 37120
rect 29276 37136 29328 37188
rect 28356 37068 28408 37120
rect 30840 37111 30892 37120
rect 30840 37077 30849 37111
rect 30849 37077 30883 37111
rect 30883 37077 30892 37111
rect 30840 37068 30892 37077
rect 47676 37136 47728 37188
rect 46940 37068 46992 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 24952 36907 25004 36916
rect 24952 36873 24961 36907
rect 24961 36873 24995 36907
rect 24995 36873 25004 36907
rect 24952 36864 25004 36873
rect 11796 36796 11848 36848
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 25228 36796 25280 36848
rect 24676 36771 24728 36780
rect 24676 36737 24685 36771
rect 24685 36737 24719 36771
rect 24719 36737 24728 36771
rect 24676 36728 24728 36737
rect 25688 36864 25740 36916
rect 25780 36864 25832 36916
rect 27252 36864 27304 36916
rect 27988 36864 28040 36916
rect 28724 36864 28776 36916
rect 26240 36796 26292 36848
rect 30840 36796 30892 36848
rect 26148 36728 26200 36780
rect 27252 36771 27304 36780
rect 27252 36737 27261 36771
rect 27261 36737 27295 36771
rect 27295 36737 27304 36771
rect 27252 36728 27304 36737
rect 27528 36771 27580 36780
rect 27528 36737 27537 36771
rect 27537 36737 27571 36771
rect 27571 36737 27580 36771
rect 27528 36728 27580 36737
rect 25688 36703 25740 36712
rect 25688 36669 25697 36703
rect 25697 36669 25731 36703
rect 25731 36669 25740 36703
rect 25688 36660 25740 36669
rect 25964 36660 26016 36712
rect 24860 36592 24912 36644
rect 21180 36524 21232 36576
rect 22376 36524 22428 36576
rect 27712 36592 27764 36644
rect 27896 36524 27948 36576
rect 29000 36660 29052 36712
rect 29828 36703 29880 36712
rect 29828 36669 29837 36703
rect 29837 36669 29871 36703
rect 29871 36669 29880 36703
rect 29828 36660 29880 36669
rect 31116 36524 31168 36576
rect 31300 36567 31352 36576
rect 31300 36533 31309 36567
rect 31309 36533 31343 36567
rect 31343 36533 31352 36567
rect 31300 36524 31352 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 9496 36320 9548 36372
rect 26424 36363 26476 36372
rect 19156 36184 19208 36236
rect 22192 36184 22244 36236
rect 23388 36227 23440 36236
rect 23388 36193 23397 36227
rect 23397 36193 23431 36227
rect 23431 36193 23440 36227
rect 23388 36184 23440 36193
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 19340 36116 19392 36168
rect 19984 36116 20036 36168
rect 24676 36252 24728 36304
rect 24860 36252 24912 36304
rect 19432 36048 19484 36100
rect 21180 36091 21232 36100
rect 21180 36057 21189 36091
rect 21189 36057 21223 36091
rect 21223 36057 21232 36091
rect 21180 36048 21232 36057
rect 21916 36048 21968 36100
rect 19984 36023 20036 36032
rect 19984 35989 19993 36023
rect 19993 35989 20027 36023
rect 20027 35989 20036 36023
rect 19984 35980 20036 35989
rect 22928 36048 22980 36100
rect 25964 36252 26016 36304
rect 25228 36184 25280 36236
rect 26424 36329 26433 36363
rect 26433 36329 26467 36363
rect 26467 36329 26476 36363
rect 26424 36320 26476 36329
rect 26792 36320 26844 36372
rect 27712 36320 27764 36372
rect 28080 36252 28132 36304
rect 29828 36320 29880 36372
rect 25412 36159 25464 36168
rect 25412 36125 25421 36159
rect 25421 36125 25455 36159
rect 25455 36125 25464 36159
rect 25412 36116 25464 36125
rect 25504 36048 25556 36100
rect 25688 36048 25740 36100
rect 26240 36159 26292 36168
rect 26240 36125 26249 36159
rect 26249 36125 26283 36159
rect 26283 36125 26292 36159
rect 26240 36116 26292 36125
rect 26884 36048 26936 36100
rect 23572 35980 23624 36032
rect 25872 35980 25924 36032
rect 27988 36116 28040 36168
rect 28540 36048 28592 36100
rect 29828 36159 29880 36168
rect 29828 36125 29837 36159
rect 29837 36125 29871 36159
rect 29871 36125 29880 36159
rect 31300 36184 31352 36236
rect 29828 36116 29880 36125
rect 30840 36116 30892 36168
rect 31024 36116 31076 36168
rect 27436 35980 27488 36032
rect 33140 35980 33192 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 28540 35819 28592 35828
rect 28540 35785 28549 35819
rect 28549 35785 28583 35819
rect 28583 35785 28592 35819
rect 28540 35776 28592 35785
rect 29828 35776 29880 35828
rect 30932 35776 30984 35828
rect 19984 35708 20036 35760
rect 21548 35708 21600 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 21824 35683 21876 35692
rect 21824 35649 21833 35683
rect 21833 35649 21867 35683
rect 21867 35649 21876 35683
rect 21824 35640 21876 35649
rect 26976 35708 27028 35760
rect 28172 35751 28224 35760
rect 22284 35640 22336 35692
rect 22376 35683 22428 35692
rect 22376 35649 22385 35683
rect 22385 35649 22419 35683
rect 22419 35649 22428 35683
rect 22376 35640 22428 35649
rect 22836 35640 22888 35692
rect 18604 35572 18656 35624
rect 19156 35615 19208 35624
rect 19156 35581 19165 35615
rect 19165 35581 19199 35615
rect 19199 35581 19208 35615
rect 19156 35572 19208 35581
rect 22652 35572 22704 35624
rect 23572 35640 23624 35692
rect 21640 35504 21692 35556
rect 24768 35572 24820 35624
rect 25596 35640 25648 35692
rect 27436 35683 27488 35692
rect 27436 35649 27445 35683
rect 27445 35649 27479 35683
rect 27479 35649 27488 35683
rect 27436 35640 27488 35649
rect 28172 35717 28181 35751
rect 28181 35717 28215 35751
rect 28215 35717 28224 35751
rect 28172 35708 28224 35717
rect 31300 35708 31352 35760
rect 33140 35708 33192 35760
rect 28356 35640 28408 35692
rect 29460 35640 29512 35692
rect 30380 35683 30432 35692
rect 30380 35649 30389 35683
rect 30389 35649 30423 35683
rect 30423 35649 30432 35683
rect 30380 35640 30432 35649
rect 30840 35683 30892 35692
rect 30840 35649 30849 35683
rect 30849 35649 30883 35683
rect 30883 35649 30892 35683
rect 30840 35640 30892 35649
rect 48136 35683 48188 35692
rect 48136 35649 48145 35683
rect 48145 35649 48179 35683
rect 48179 35649 48188 35683
rect 48136 35640 48188 35649
rect 25688 35572 25740 35624
rect 2228 35436 2280 35488
rect 24676 35479 24728 35488
rect 24676 35445 24685 35479
rect 24685 35445 24719 35479
rect 24719 35445 24728 35479
rect 24676 35436 24728 35445
rect 25872 35504 25924 35556
rect 27160 35572 27212 35624
rect 29092 35572 29144 35624
rect 32128 35615 32180 35624
rect 32128 35581 32137 35615
rect 32137 35581 32171 35615
rect 32171 35581 32180 35615
rect 32128 35572 32180 35581
rect 32496 35572 32548 35624
rect 28264 35504 28316 35556
rect 25780 35436 25832 35488
rect 31024 35436 31076 35488
rect 32036 35436 32088 35488
rect 47124 35436 47176 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 21640 35275 21692 35284
rect 21640 35241 21649 35275
rect 21649 35241 21683 35275
rect 21683 35241 21692 35275
rect 21640 35232 21692 35241
rect 21824 35275 21876 35284
rect 21824 35241 21833 35275
rect 21833 35241 21867 35275
rect 21867 35241 21876 35275
rect 21824 35232 21876 35241
rect 22560 35232 22612 35284
rect 23388 35232 23440 35284
rect 24584 35232 24636 35284
rect 24768 35275 24820 35284
rect 24768 35241 24777 35275
rect 24777 35241 24811 35275
rect 24811 35241 24820 35275
rect 24768 35232 24820 35241
rect 27252 35232 27304 35284
rect 28080 35275 28132 35284
rect 28080 35241 28089 35275
rect 28089 35241 28123 35275
rect 28123 35241 28132 35275
rect 28080 35232 28132 35241
rect 28540 35275 28592 35284
rect 28540 35241 28549 35275
rect 28549 35241 28583 35275
rect 28583 35241 28592 35275
rect 28540 35232 28592 35241
rect 28908 35232 28960 35284
rect 31852 35232 31904 35284
rect 32496 35275 32548 35284
rect 32496 35241 32505 35275
rect 32505 35241 32539 35275
rect 32539 35241 32548 35275
rect 32496 35232 32548 35241
rect 25504 35164 25556 35216
rect 23480 35096 23532 35148
rect 28724 35164 28776 35216
rect 31944 35164 31996 35216
rect 20352 35028 20404 35080
rect 22100 35028 22152 35080
rect 22652 35071 22704 35080
rect 22652 35037 22661 35071
rect 22661 35037 22695 35071
rect 22695 35037 22704 35071
rect 22652 35028 22704 35037
rect 26332 35028 26384 35080
rect 27160 35071 27212 35080
rect 27160 35037 27169 35071
rect 27169 35037 27203 35071
rect 27203 35037 27212 35071
rect 27160 35028 27212 35037
rect 27804 35096 27856 35148
rect 32036 35139 32088 35148
rect 27896 35028 27948 35080
rect 28264 35071 28316 35080
rect 28264 35037 28273 35071
rect 28273 35037 28307 35071
rect 28307 35037 28316 35071
rect 28264 35028 28316 35037
rect 28356 35071 28408 35080
rect 28356 35037 28365 35071
rect 28365 35037 28399 35071
rect 28399 35037 28408 35071
rect 28632 35071 28684 35080
rect 28356 35028 28408 35037
rect 28632 35037 28641 35071
rect 28641 35037 28675 35071
rect 28675 35037 28684 35071
rect 28632 35028 28684 35037
rect 29092 35028 29144 35080
rect 30104 35071 30156 35080
rect 23572 34960 23624 35012
rect 24584 35003 24636 35012
rect 24584 34969 24593 35003
rect 24593 34969 24627 35003
rect 24627 34969 24636 35003
rect 24584 34960 24636 34969
rect 27344 35003 27396 35012
rect 27344 34969 27354 35003
rect 27354 34969 27388 35003
rect 27388 34969 27396 35003
rect 27344 34960 27396 34969
rect 27436 35003 27488 35012
rect 27436 34969 27471 35003
rect 27471 34969 27488 35003
rect 30104 35037 30113 35071
rect 30113 35037 30147 35071
rect 30147 35037 30156 35071
rect 30104 35028 30156 35037
rect 30932 35071 30984 35080
rect 30932 35037 30941 35071
rect 30941 35037 30975 35071
rect 30975 35037 30984 35071
rect 30932 35028 30984 35037
rect 31024 35071 31076 35080
rect 31024 35037 31033 35071
rect 31033 35037 31067 35071
rect 31067 35037 31076 35071
rect 31024 35028 31076 35037
rect 27436 34960 27488 34969
rect 30564 34960 30616 35012
rect 22468 34892 22520 34944
rect 27712 34892 27764 34944
rect 31668 35028 31720 35080
rect 32036 35105 32045 35139
rect 32045 35105 32079 35139
rect 32079 35105 32088 35139
rect 32036 35096 32088 35105
rect 32864 35096 32916 35148
rect 31852 35028 31904 35080
rect 32312 35071 32364 35080
rect 32312 35037 32321 35071
rect 32321 35037 32355 35071
rect 32355 35037 32364 35071
rect 32312 35028 32364 35037
rect 48228 35028 48280 35080
rect 47860 34892 47912 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 20260 34688 20312 34740
rect 20536 34688 20588 34740
rect 19616 34620 19668 34672
rect 26976 34688 27028 34740
rect 28908 34731 28960 34740
rect 28908 34697 28917 34731
rect 28917 34697 28951 34731
rect 28951 34697 28960 34731
rect 28908 34688 28960 34697
rect 30840 34688 30892 34740
rect 31208 34688 31260 34740
rect 26332 34620 26384 34672
rect 28172 34620 28224 34672
rect 18604 34527 18656 34536
rect 18604 34493 18613 34527
rect 18613 34493 18647 34527
rect 18647 34493 18656 34527
rect 18604 34484 18656 34493
rect 21088 34484 21140 34536
rect 22928 34595 22980 34604
rect 22928 34561 22937 34595
rect 22937 34561 22971 34595
rect 22971 34561 22980 34595
rect 22928 34552 22980 34561
rect 24584 34595 24636 34604
rect 24584 34561 24593 34595
rect 24593 34561 24627 34595
rect 24627 34561 24636 34595
rect 24584 34552 24636 34561
rect 27436 34552 27488 34604
rect 30288 34620 30340 34672
rect 30472 34620 30524 34672
rect 28816 34552 28868 34604
rect 22560 34484 22612 34536
rect 25136 34484 25188 34536
rect 27160 34484 27212 34536
rect 27712 34484 27764 34536
rect 27528 34416 27580 34468
rect 28080 34484 28132 34536
rect 29368 34484 29420 34536
rect 30104 34552 30156 34604
rect 30840 34552 30892 34604
rect 47768 34595 47820 34604
rect 47768 34561 47777 34595
rect 47777 34561 47811 34595
rect 47811 34561 47820 34595
rect 47768 34552 47820 34561
rect 20260 34348 20312 34400
rect 22560 34348 22612 34400
rect 23204 34348 23256 34400
rect 28816 34416 28868 34468
rect 30472 34416 30524 34468
rect 31024 34484 31076 34536
rect 30656 34416 30708 34468
rect 30380 34391 30432 34400
rect 30380 34357 30389 34391
rect 30389 34357 30423 34391
rect 30423 34357 30432 34391
rect 30380 34348 30432 34357
rect 30564 34348 30616 34400
rect 47216 34348 47268 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19616 34187 19668 34196
rect 19616 34153 19625 34187
rect 19625 34153 19659 34187
rect 19659 34153 19668 34187
rect 19616 34144 19668 34153
rect 20260 34144 20312 34196
rect 22100 34144 22152 34196
rect 23848 34144 23900 34196
rect 25228 34144 25280 34196
rect 28816 34144 28868 34196
rect 30104 34144 30156 34196
rect 30656 34076 30708 34128
rect 1952 34008 2004 34060
rect 20536 33940 20588 33992
rect 20996 33983 21048 33992
rect 20996 33949 21005 33983
rect 21005 33949 21039 33983
rect 21039 33949 21048 33983
rect 20996 33940 21048 33949
rect 21088 33983 21140 33992
rect 21088 33949 21097 33983
rect 21097 33949 21131 33983
rect 21131 33949 21140 33983
rect 21088 33940 21140 33949
rect 22008 33983 22060 33992
rect 22008 33949 22017 33983
rect 22017 33949 22051 33983
rect 22051 33949 22060 33983
rect 22008 33940 22060 33949
rect 22192 34008 22244 34060
rect 23296 34008 23348 34060
rect 22560 33940 22612 33992
rect 22744 33940 22796 33992
rect 23020 33983 23072 33992
rect 23020 33949 23029 33983
rect 23029 33949 23063 33983
rect 23063 33949 23072 33983
rect 23020 33940 23072 33949
rect 28632 34008 28684 34060
rect 31392 34008 31444 34060
rect 47124 34051 47176 34060
rect 47124 34017 47133 34051
rect 47133 34017 47167 34051
rect 47167 34017 47176 34051
rect 47124 34008 47176 34017
rect 47676 34051 47728 34060
rect 47676 34017 47685 34051
rect 47685 34017 47719 34051
rect 47719 34017 47728 34051
rect 47676 34008 47728 34017
rect 29552 33940 29604 33992
rect 30012 33983 30064 33992
rect 30012 33949 30021 33983
rect 30021 33949 30055 33983
rect 30055 33949 30064 33983
rect 30012 33940 30064 33949
rect 24676 33915 24728 33924
rect 24676 33881 24685 33915
rect 24685 33881 24719 33915
rect 24719 33881 24728 33915
rect 24676 33872 24728 33881
rect 25136 33872 25188 33924
rect 27252 33915 27304 33924
rect 27252 33881 27261 33915
rect 27261 33881 27295 33915
rect 27295 33881 27304 33915
rect 27252 33872 27304 33881
rect 28264 33872 28316 33924
rect 28908 33872 28960 33924
rect 30840 33940 30892 33992
rect 47216 33915 47268 33924
rect 47216 33881 47225 33915
rect 47225 33881 47259 33915
rect 47259 33881 47268 33915
rect 47216 33872 47268 33881
rect 23572 33804 23624 33856
rect 25320 33804 25372 33856
rect 27344 33847 27396 33856
rect 27344 33813 27353 33847
rect 27353 33813 27387 33847
rect 27387 33813 27396 33847
rect 27344 33804 27396 33813
rect 28724 33804 28776 33856
rect 29276 33804 29328 33856
rect 30564 33804 30616 33856
rect 31300 33804 31352 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 23296 33643 23348 33652
rect 23296 33609 23305 33643
rect 23305 33609 23339 33643
rect 23339 33609 23348 33643
rect 23296 33600 23348 33609
rect 47768 33600 47820 33652
rect 25044 33532 25096 33584
rect 29276 33575 29328 33584
rect 29276 33541 29285 33575
rect 29285 33541 29319 33575
rect 29319 33541 29328 33575
rect 29276 33532 29328 33541
rect 1584 33507 1636 33516
rect 1584 33473 1593 33507
rect 1593 33473 1627 33507
rect 1627 33473 1636 33507
rect 1584 33464 1636 33473
rect 2228 33507 2280 33516
rect 2228 33473 2237 33507
rect 2237 33473 2271 33507
rect 2271 33473 2280 33507
rect 2228 33464 2280 33473
rect 20536 33464 20588 33516
rect 22008 33507 22060 33516
rect 22008 33473 22017 33507
rect 22017 33473 22051 33507
rect 22051 33473 22060 33507
rect 22008 33464 22060 33473
rect 24124 33507 24176 33516
rect 24124 33473 24153 33507
rect 24153 33473 24176 33507
rect 25228 33507 25280 33516
rect 24124 33464 24176 33473
rect 3792 33396 3844 33448
rect 4620 33396 4672 33448
rect 23664 33396 23716 33448
rect 23940 33439 23992 33448
rect 23940 33405 23949 33439
rect 23949 33405 23983 33439
rect 23983 33405 23992 33439
rect 23940 33396 23992 33405
rect 25228 33473 25237 33507
rect 25237 33473 25271 33507
rect 25271 33473 25280 33507
rect 25228 33464 25280 33473
rect 25320 33507 25372 33516
rect 25320 33473 25329 33507
rect 25329 33473 25363 33507
rect 25363 33473 25372 33507
rect 25320 33464 25372 33473
rect 24400 33371 24452 33380
rect 24400 33337 24409 33371
rect 24409 33337 24443 33371
rect 24443 33337 24452 33371
rect 24400 33328 24452 33337
rect 24492 33328 24544 33380
rect 27344 33464 27396 33516
rect 30380 33464 30432 33516
rect 46848 33507 46900 33516
rect 46848 33473 46857 33507
rect 46857 33473 46891 33507
rect 46891 33473 46900 33507
rect 46848 33464 46900 33473
rect 47308 33464 47360 33516
rect 29000 33439 29052 33448
rect 29000 33405 29009 33439
rect 29009 33405 29043 33439
rect 29043 33405 29052 33439
rect 29000 33396 29052 33405
rect 29276 33396 29328 33448
rect 30012 33396 30064 33448
rect 2780 33260 2832 33312
rect 19984 33260 20036 33312
rect 21824 33303 21876 33312
rect 21824 33269 21833 33303
rect 21833 33269 21867 33303
rect 21867 33269 21876 33303
rect 21824 33260 21876 33269
rect 22192 33303 22244 33312
rect 22192 33269 22201 33303
rect 22201 33269 22235 33303
rect 22235 33269 22244 33303
rect 22192 33260 22244 33269
rect 22560 33260 22612 33312
rect 24952 33260 25004 33312
rect 44180 33328 44232 33380
rect 30656 33260 30708 33312
rect 46940 33303 46992 33312
rect 46940 33269 46949 33303
rect 46949 33269 46983 33303
rect 46983 33269 46992 33303
rect 46940 33260 46992 33269
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2780 33099 2832 33108
rect 2780 33065 2789 33099
rect 2789 33065 2823 33099
rect 2823 33065 2832 33099
rect 2780 33056 2832 33065
rect 3792 33099 3844 33108
rect 3792 33065 3801 33099
rect 3801 33065 3835 33099
rect 3835 33065 3844 33099
rect 3792 33056 3844 33065
rect 22008 33056 22060 33108
rect 22192 33056 22244 33108
rect 24400 33056 24452 33108
rect 27988 33056 28040 33108
rect 28356 33056 28408 33108
rect 29000 33056 29052 33108
rect 32128 33056 32180 33108
rect 1400 32963 1452 32972
rect 1400 32929 1409 32963
rect 1409 32929 1443 32963
rect 1443 32929 1452 32963
rect 1400 32920 1452 32929
rect 2688 32895 2740 32904
rect 2688 32861 2697 32895
rect 2697 32861 2731 32895
rect 2731 32861 2740 32895
rect 2688 32852 2740 32861
rect 21824 32920 21876 32972
rect 18144 32852 18196 32904
rect 18604 32852 18656 32904
rect 25228 32988 25280 33040
rect 22284 32920 22336 32972
rect 24676 32920 24728 32972
rect 19984 32784 20036 32836
rect 22560 32852 22612 32904
rect 22928 32895 22980 32904
rect 22928 32861 22937 32895
rect 22937 32861 22971 32895
rect 22971 32861 22980 32895
rect 22928 32852 22980 32861
rect 23940 32852 23992 32904
rect 24952 32920 25004 32972
rect 29276 32988 29328 33040
rect 29552 33031 29604 33040
rect 29552 32997 29561 33031
rect 29561 32997 29595 33031
rect 29595 32997 29604 33031
rect 29552 32988 29604 32997
rect 27252 32920 27304 32972
rect 28172 32895 28224 32904
rect 23664 32784 23716 32836
rect 28172 32861 28181 32895
rect 28181 32861 28215 32895
rect 28215 32861 28224 32895
rect 28172 32852 28224 32861
rect 27988 32784 28040 32836
rect 19432 32716 19484 32768
rect 20260 32716 20312 32768
rect 21272 32716 21324 32768
rect 27160 32716 27212 32768
rect 27436 32759 27488 32768
rect 27436 32725 27445 32759
rect 27445 32725 27479 32759
rect 27479 32725 27488 32759
rect 28816 32852 28868 32904
rect 30656 32988 30708 33040
rect 31392 33031 31444 33040
rect 31392 32997 31401 33031
rect 31401 32997 31435 33031
rect 31435 32997 31444 33031
rect 31392 32988 31444 32997
rect 32036 32988 32088 33040
rect 46204 33056 46256 33108
rect 46480 33056 46532 33108
rect 31300 32895 31352 32904
rect 28724 32784 28776 32836
rect 31300 32861 31309 32895
rect 31309 32861 31343 32895
rect 31343 32861 31352 32895
rect 31300 32852 31352 32861
rect 31392 32852 31444 32904
rect 31576 32852 31628 32904
rect 32588 32895 32640 32904
rect 32588 32861 32597 32895
rect 32597 32861 32631 32895
rect 32631 32861 32640 32895
rect 32588 32852 32640 32861
rect 46296 32852 46348 32904
rect 30656 32827 30708 32836
rect 30656 32793 30665 32827
rect 30665 32793 30699 32827
rect 30699 32793 30708 32827
rect 30656 32784 30708 32793
rect 30748 32784 30800 32836
rect 32036 32784 32088 32836
rect 32404 32784 32456 32836
rect 27436 32716 27488 32725
rect 31024 32716 31076 32768
rect 32496 32759 32548 32768
rect 32496 32725 32505 32759
rect 32505 32725 32539 32759
rect 32539 32725 32548 32759
rect 32496 32716 32548 32725
rect 46848 32716 46900 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 19984 32512 20036 32564
rect 20536 32512 20588 32564
rect 22928 32512 22980 32564
rect 23480 32512 23532 32564
rect 25044 32555 25096 32564
rect 25044 32521 25053 32555
rect 25053 32521 25087 32555
rect 25087 32521 25096 32555
rect 25044 32512 25096 32521
rect 30380 32512 30432 32564
rect 30472 32512 30524 32564
rect 31024 32512 31076 32564
rect 31576 32555 31628 32564
rect 19432 32444 19484 32496
rect 20260 32444 20312 32496
rect 30748 32444 30800 32496
rect 30932 32444 30984 32496
rect 31576 32521 31585 32555
rect 31585 32521 31619 32555
rect 31619 32521 31628 32555
rect 31576 32512 31628 32521
rect 46940 32512 46992 32564
rect 32404 32487 32456 32496
rect 32404 32453 32413 32487
rect 32413 32453 32447 32487
rect 32447 32453 32456 32487
rect 32404 32444 32456 32453
rect 33416 32444 33468 32496
rect 18144 32419 18196 32428
rect 18144 32385 18153 32419
rect 18153 32385 18187 32419
rect 18187 32385 18196 32419
rect 18144 32376 18196 32385
rect 21916 32376 21968 32428
rect 1676 32308 1728 32360
rect 2228 32308 2280 32360
rect 2780 32351 2832 32360
rect 2780 32317 2789 32351
rect 2789 32317 2823 32351
rect 2823 32317 2832 32351
rect 2780 32308 2832 32317
rect 20536 32308 20588 32360
rect 21272 32351 21324 32360
rect 21272 32317 21281 32351
rect 21281 32317 21315 32351
rect 21315 32317 21324 32351
rect 21272 32308 21324 32317
rect 23204 32351 23256 32360
rect 23204 32317 23213 32351
rect 23213 32317 23247 32351
rect 23247 32317 23256 32351
rect 23204 32308 23256 32317
rect 23388 32419 23440 32428
rect 23388 32385 23397 32419
rect 23397 32385 23431 32419
rect 23431 32385 23440 32419
rect 23388 32376 23440 32385
rect 24124 32376 24176 32428
rect 24860 32376 24912 32428
rect 27068 32376 27120 32428
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 28172 32376 28224 32428
rect 29092 32376 29144 32428
rect 25228 32308 25280 32360
rect 29368 32308 29420 32360
rect 21088 32215 21140 32224
rect 21088 32181 21097 32215
rect 21097 32181 21131 32215
rect 21131 32181 21140 32215
rect 21088 32172 21140 32181
rect 27620 32240 27672 32292
rect 28264 32240 28316 32292
rect 24400 32215 24452 32224
rect 24400 32181 24409 32215
rect 24409 32181 24443 32215
rect 24443 32181 24452 32215
rect 24400 32172 24452 32181
rect 26332 32172 26384 32224
rect 27160 32172 27212 32224
rect 29920 32172 29972 32224
rect 31116 32376 31168 32428
rect 31484 32376 31536 32428
rect 32128 32419 32180 32428
rect 32128 32385 32137 32419
rect 32137 32385 32171 32419
rect 32171 32385 32180 32419
rect 32128 32376 32180 32385
rect 46480 32376 46532 32428
rect 32772 32172 32824 32224
rect 46480 32172 46532 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1676 32011 1728 32020
rect 1676 31977 1685 32011
rect 1685 31977 1719 32011
rect 1719 31977 1728 32011
rect 1676 31968 1728 31977
rect 2228 32011 2280 32020
rect 2228 31977 2237 32011
rect 2237 31977 2271 32011
rect 2271 31977 2280 32011
rect 2228 31968 2280 31977
rect 19432 32011 19484 32020
rect 19432 31977 19441 32011
rect 19441 31977 19475 32011
rect 19475 31977 19484 32011
rect 19432 31968 19484 31977
rect 21916 32011 21968 32020
rect 21916 31977 21925 32011
rect 21925 31977 21959 32011
rect 21959 31977 21968 32011
rect 21916 31968 21968 31977
rect 24768 32011 24820 32020
rect 24768 31977 24777 32011
rect 24777 31977 24811 32011
rect 24811 31977 24820 32011
rect 24768 31968 24820 31977
rect 25228 32011 25280 32020
rect 25228 31977 25237 32011
rect 25237 31977 25271 32011
rect 25271 31977 25280 32011
rect 25228 31968 25280 31977
rect 23940 31900 23992 31952
rect 2688 31832 2740 31884
rect 4620 31875 4672 31884
rect 4620 31841 4629 31875
rect 4629 31841 4663 31875
rect 4663 31841 4672 31875
rect 4620 31832 4672 31841
rect 5448 31832 5500 31884
rect 21272 31832 21324 31884
rect 2320 31764 2372 31816
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 18144 31764 18196 31816
rect 18512 31764 18564 31816
rect 19984 31764 20036 31816
rect 21088 31764 21140 31816
rect 24400 31832 24452 31884
rect 24860 31875 24912 31884
rect 24860 31841 24869 31875
rect 24869 31841 24903 31875
rect 24903 31841 24912 31875
rect 24860 31832 24912 31841
rect 29000 31968 29052 32020
rect 32588 31968 32640 32020
rect 33416 31968 33468 32020
rect 48044 31968 48096 32020
rect 26332 31875 26384 31884
rect 26332 31841 26341 31875
rect 26341 31841 26375 31875
rect 26375 31841 26384 31875
rect 26332 31832 26384 31841
rect 27344 31832 27396 31884
rect 27528 31832 27580 31884
rect 27988 31832 28040 31884
rect 46296 31875 46348 31884
rect 23388 31764 23440 31816
rect 24124 31764 24176 31816
rect 22100 31696 22152 31748
rect 23296 31696 23348 31748
rect 28264 31807 28316 31816
rect 28264 31773 28273 31807
rect 28273 31773 28307 31807
rect 28307 31773 28316 31807
rect 29920 31807 29972 31816
rect 28264 31764 28316 31773
rect 29920 31773 29929 31807
rect 29929 31773 29963 31807
rect 29963 31773 29972 31807
rect 29920 31764 29972 31773
rect 30012 31764 30064 31816
rect 31484 31764 31536 31816
rect 46296 31841 46305 31875
rect 46305 31841 46339 31875
rect 46339 31841 46348 31875
rect 46296 31832 46348 31841
rect 46480 31875 46532 31884
rect 46480 31841 46489 31875
rect 46489 31841 46523 31875
rect 46523 31841 46532 31875
rect 46480 31832 46532 31841
rect 48136 31875 48188 31884
rect 48136 31841 48145 31875
rect 48145 31841 48179 31875
rect 48179 31841 48188 31875
rect 48136 31832 48188 31841
rect 32588 31764 32640 31816
rect 32772 31764 32824 31816
rect 34612 31764 34664 31816
rect 18512 31628 18564 31680
rect 23204 31628 23256 31680
rect 27344 31628 27396 31680
rect 28724 31628 28776 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 24584 31424 24636 31476
rect 27068 31424 27120 31476
rect 18512 31399 18564 31408
rect 18512 31365 18521 31399
rect 18521 31365 18555 31399
rect 18555 31365 18564 31399
rect 18512 31356 18564 31365
rect 18144 31288 18196 31340
rect 21916 31288 21968 31340
rect 20260 31220 20312 31272
rect 22100 31263 22152 31272
rect 22100 31229 22109 31263
rect 22109 31229 22143 31263
rect 22143 31229 22152 31263
rect 22100 31220 22152 31229
rect 23112 31288 23164 31340
rect 24860 31356 24912 31408
rect 23940 31331 23992 31340
rect 23940 31297 23949 31331
rect 23949 31297 23983 31331
rect 23983 31297 23992 31331
rect 23940 31288 23992 31297
rect 24124 31288 24176 31340
rect 24584 31331 24636 31340
rect 24584 31297 24593 31331
rect 24593 31297 24627 31331
rect 24627 31297 24636 31331
rect 24584 31288 24636 31297
rect 26148 31356 26200 31408
rect 26700 31288 26752 31340
rect 27160 31288 27212 31340
rect 27344 31331 27396 31340
rect 27344 31297 27353 31331
rect 27353 31297 27387 31331
rect 27387 31297 27396 31331
rect 27344 31288 27396 31297
rect 27620 31288 27672 31340
rect 31484 31220 31536 31272
rect 21824 31084 21876 31136
rect 23296 31152 23348 31204
rect 23480 31084 23532 31136
rect 26240 31127 26292 31136
rect 26240 31093 26249 31127
rect 26249 31093 26283 31127
rect 26283 31093 26292 31127
rect 26240 31084 26292 31093
rect 27068 31084 27120 31136
rect 30564 31152 30616 31204
rect 31024 31127 31076 31136
rect 31024 31093 31048 31127
rect 31048 31093 31076 31127
rect 31024 31084 31076 31093
rect 31116 31127 31168 31136
rect 31116 31093 31125 31127
rect 31125 31093 31159 31127
rect 31159 31093 31168 31127
rect 31116 31084 31168 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 20536 30880 20588 30932
rect 23940 30880 23992 30932
rect 25320 30880 25372 30932
rect 26148 30880 26200 30932
rect 27436 30880 27488 30932
rect 31760 30880 31812 30932
rect 32496 30880 32548 30932
rect 29092 30812 29144 30864
rect 21088 30744 21140 30796
rect 23480 30787 23532 30796
rect 21180 30676 21232 30728
rect 21824 30719 21876 30728
rect 21824 30685 21833 30719
rect 21833 30685 21867 30719
rect 21867 30685 21876 30719
rect 21824 30676 21876 30685
rect 21916 30719 21968 30728
rect 21916 30685 21926 30719
rect 21926 30685 21960 30719
rect 21960 30685 21968 30719
rect 21916 30676 21968 30685
rect 23204 30719 23256 30728
rect 22008 30608 22060 30660
rect 20812 30540 20864 30592
rect 20904 30540 20956 30592
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 23480 30753 23489 30787
rect 23489 30753 23523 30787
rect 23523 30753 23532 30787
rect 23480 30744 23532 30753
rect 24768 30744 24820 30796
rect 27068 30787 27120 30796
rect 23848 30676 23900 30728
rect 27068 30753 27077 30787
rect 27077 30753 27111 30787
rect 27111 30753 27120 30787
rect 27068 30744 27120 30753
rect 29000 30744 29052 30796
rect 31024 30812 31076 30864
rect 30840 30744 30892 30796
rect 26056 30676 26108 30728
rect 27528 30676 27580 30728
rect 27712 30676 27764 30728
rect 28080 30676 28132 30728
rect 28264 30676 28316 30728
rect 28632 30676 28684 30728
rect 31944 30744 31996 30796
rect 32588 30744 32640 30796
rect 33048 30744 33100 30796
rect 47676 30787 47728 30796
rect 47676 30753 47685 30787
rect 47685 30753 47719 30787
rect 47719 30753 47728 30787
rect 47676 30744 47728 30753
rect 48044 30744 48096 30796
rect 32036 30719 32088 30728
rect 25596 30608 25648 30660
rect 29828 30651 29880 30660
rect 29828 30617 29837 30651
rect 29837 30617 29871 30651
rect 29871 30617 29880 30651
rect 29828 30608 29880 30617
rect 23756 30583 23808 30592
rect 23756 30549 23765 30583
rect 23765 30549 23799 30583
rect 23799 30549 23808 30583
rect 23756 30540 23808 30549
rect 25228 30540 25280 30592
rect 31116 30608 31168 30660
rect 31576 30608 31628 30660
rect 32036 30685 32045 30719
rect 32045 30685 32079 30719
rect 32079 30685 32088 30719
rect 32036 30676 32088 30685
rect 33692 30676 33744 30728
rect 32680 30608 32732 30660
rect 33876 30583 33928 30592
rect 33876 30549 33885 30583
rect 33885 30549 33919 30583
rect 33919 30549 33928 30583
rect 33876 30540 33928 30549
rect 34520 30608 34572 30660
rect 35992 30608 36044 30660
rect 46112 30608 46164 30660
rect 47308 30608 47360 30660
rect 47952 30608 48004 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4620 30336 4672 30388
rect 20904 30336 20956 30388
rect 14096 30200 14148 30252
rect 17316 30200 17368 30252
rect 19340 30200 19392 30252
rect 20628 30200 20680 30252
rect 23664 30268 23716 30320
rect 20812 30243 20864 30252
rect 20812 30209 20821 30243
rect 20821 30209 20855 30243
rect 20855 30209 20864 30243
rect 20812 30200 20864 30209
rect 21180 30200 21232 30252
rect 17408 30175 17460 30184
rect 17408 30141 17417 30175
rect 17417 30141 17451 30175
rect 17451 30141 17460 30175
rect 17408 30132 17460 30141
rect 17592 30175 17644 30184
rect 17592 30141 17601 30175
rect 17601 30141 17635 30175
rect 17635 30141 17644 30175
rect 17592 30132 17644 30141
rect 20996 30132 21048 30184
rect 23204 30132 23256 30184
rect 24952 30268 25004 30320
rect 25136 30268 25188 30320
rect 29828 30336 29880 30388
rect 29276 30311 29328 30320
rect 25228 30243 25280 30252
rect 25228 30209 25237 30243
rect 25237 30209 25271 30243
rect 25271 30209 25280 30243
rect 25228 30200 25280 30209
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 29276 30277 29285 30311
rect 29285 30277 29319 30311
rect 29319 30277 29328 30311
rect 29276 30268 29328 30277
rect 30472 30268 30524 30320
rect 27068 30243 27120 30252
rect 27068 30209 27077 30243
rect 27077 30209 27111 30243
rect 27111 30209 27120 30243
rect 27068 30200 27120 30209
rect 28172 30243 28224 30252
rect 28172 30209 28181 30243
rect 28181 30209 28215 30243
rect 28215 30209 28224 30243
rect 28172 30200 28224 30209
rect 28724 30200 28776 30252
rect 29092 30202 29144 30254
rect 29184 30243 29236 30252
rect 29184 30209 29193 30243
rect 29193 30209 29227 30243
rect 29227 30209 29236 30243
rect 29184 30200 29236 30209
rect 29460 30200 29512 30252
rect 30932 30200 30984 30252
rect 31392 30200 31444 30252
rect 32036 30200 32088 30252
rect 32772 30200 32824 30252
rect 33416 30243 33468 30252
rect 33416 30209 33425 30243
rect 33425 30209 33459 30243
rect 33459 30209 33468 30243
rect 33416 30200 33468 30209
rect 33508 30200 33560 30252
rect 34520 30268 34572 30320
rect 35992 30268 36044 30320
rect 33692 30243 33744 30252
rect 33692 30209 33701 30243
rect 33701 30209 33735 30243
rect 33735 30209 33744 30243
rect 33968 30243 34020 30252
rect 33692 30200 33744 30209
rect 33968 30209 33977 30243
rect 33977 30209 34011 30243
rect 34011 30209 34020 30243
rect 33968 30200 34020 30209
rect 34612 30200 34664 30252
rect 27528 30132 27580 30184
rect 28448 30132 28500 30184
rect 32404 30175 32456 30184
rect 32404 30141 32413 30175
rect 32413 30141 32447 30175
rect 32447 30141 32456 30175
rect 32404 30132 32456 30141
rect 34152 30132 34204 30184
rect 46848 30132 46900 30184
rect 14924 29996 14976 30048
rect 19800 30039 19852 30048
rect 19800 30005 19809 30039
rect 19809 30005 19843 30039
rect 19843 30005 19852 30039
rect 19800 29996 19852 30005
rect 21272 30039 21324 30048
rect 21272 30005 21281 30039
rect 21281 30005 21315 30039
rect 21315 30005 21324 30039
rect 21272 29996 21324 30005
rect 24216 30039 24268 30048
rect 24216 30005 24225 30039
rect 24225 30005 24259 30039
rect 24259 30005 24268 30039
rect 24216 29996 24268 30005
rect 24492 29996 24544 30048
rect 26884 29996 26936 30048
rect 27528 29996 27580 30048
rect 28356 30039 28408 30048
rect 28356 30005 28365 30039
rect 28365 30005 28399 30039
rect 28399 30005 28408 30039
rect 28356 29996 28408 30005
rect 29184 29996 29236 30048
rect 29368 29996 29420 30048
rect 30104 29996 30156 30048
rect 30840 30039 30892 30048
rect 30840 30005 30849 30039
rect 30849 30005 30883 30039
rect 30883 30005 30892 30039
rect 30840 29996 30892 30005
rect 32036 29996 32088 30048
rect 33048 29996 33100 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 28080 29792 28132 29844
rect 28632 29835 28684 29844
rect 28632 29801 28641 29835
rect 28641 29801 28675 29835
rect 28675 29801 28684 29835
rect 28632 29792 28684 29801
rect 32496 29792 32548 29844
rect 33416 29792 33468 29844
rect 27528 29724 27580 29776
rect 14924 29699 14976 29708
rect 14924 29665 14933 29699
rect 14933 29665 14967 29699
rect 14967 29665 14976 29699
rect 14924 29656 14976 29665
rect 16488 29699 16540 29708
rect 16488 29665 16497 29699
rect 16497 29665 16531 29699
rect 16531 29665 16540 29699
rect 16488 29656 16540 29665
rect 21272 29656 21324 29708
rect 14096 29631 14148 29640
rect 14096 29597 14105 29631
rect 14105 29597 14139 29631
rect 14139 29597 14148 29631
rect 14096 29588 14148 29597
rect 14740 29631 14792 29640
rect 14740 29597 14749 29631
rect 14749 29597 14783 29631
rect 14783 29597 14792 29631
rect 14740 29588 14792 29597
rect 19156 29588 19208 29640
rect 23756 29656 23808 29708
rect 23204 29631 23256 29640
rect 23204 29597 23213 29631
rect 23213 29597 23247 29631
rect 23247 29597 23256 29631
rect 23204 29588 23256 29597
rect 19800 29520 19852 29572
rect 23388 29631 23440 29640
rect 23388 29597 23397 29631
rect 23397 29597 23431 29631
rect 23431 29597 23440 29631
rect 23388 29588 23440 29597
rect 23664 29588 23716 29640
rect 24768 29656 24820 29708
rect 24492 29631 24544 29640
rect 24492 29597 24501 29631
rect 24501 29597 24535 29631
rect 24535 29597 24544 29631
rect 24492 29588 24544 29597
rect 26056 29656 26108 29708
rect 25228 29588 25280 29640
rect 25596 29631 25648 29640
rect 25596 29597 25605 29631
rect 25605 29597 25639 29631
rect 25639 29597 25648 29631
rect 25596 29588 25648 29597
rect 30748 29724 30800 29776
rect 30932 29724 30984 29776
rect 27988 29656 28040 29708
rect 30472 29656 30524 29708
rect 30840 29656 30892 29708
rect 24768 29563 24820 29572
rect 24768 29529 24777 29563
rect 24777 29529 24811 29563
rect 24811 29529 24820 29563
rect 24768 29520 24820 29529
rect 28080 29588 28132 29640
rect 28172 29588 28224 29640
rect 30564 29631 30616 29640
rect 30564 29597 30573 29631
rect 30573 29597 30607 29631
rect 30607 29597 30616 29631
rect 30564 29588 30616 29597
rect 31484 29588 31536 29640
rect 32128 29588 32180 29640
rect 33876 29724 33928 29776
rect 32588 29699 32640 29708
rect 32588 29665 32597 29699
rect 32597 29665 32631 29699
rect 32631 29665 32640 29699
rect 32588 29656 32640 29665
rect 40224 29656 40276 29708
rect 47216 29656 47268 29708
rect 14464 29452 14516 29504
rect 21180 29452 21232 29504
rect 23572 29452 23624 29504
rect 23848 29452 23900 29504
rect 26700 29520 26752 29572
rect 27436 29520 27488 29572
rect 29276 29520 29328 29572
rect 32036 29520 32088 29572
rect 32956 29588 33008 29640
rect 33508 29631 33560 29640
rect 33508 29597 33517 29631
rect 33517 29597 33551 29631
rect 33551 29597 33560 29631
rect 33508 29588 33560 29597
rect 33600 29631 33652 29640
rect 33600 29597 33609 29631
rect 33609 29597 33643 29631
rect 33643 29597 33652 29631
rect 33876 29631 33928 29640
rect 33600 29588 33652 29597
rect 33876 29597 33885 29631
rect 33885 29597 33919 29631
rect 33919 29597 33928 29631
rect 33876 29588 33928 29597
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 24952 29452 25004 29504
rect 25688 29495 25740 29504
rect 25688 29461 25697 29495
rect 25697 29461 25731 29495
rect 25731 29461 25740 29495
rect 25688 29452 25740 29461
rect 26240 29452 26292 29504
rect 26976 29452 27028 29504
rect 27252 29452 27304 29504
rect 31484 29452 31536 29504
rect 32404 29452 32456 29504
rect 32496 29452 32548 29504
rect 34244 29452 34296 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 12440 29180 12492 29232
rect 14464 29223 14516 29232
rect 14464 29189 14473 29223
rect 14473 29189 14507 29223
rect 14507 29189 14516 29223
rect 14464 29180 14516 29189
rect 11060 29112 11112 29164
rect 18512 29112 18564 29164
rect 19340 29112 19392 29164
rect 20352 29248 20404 29300
rect 20996 29248 21048 29300
rect 24860 29248 24912 29300
rect 27712 29291 27764 29300
rect 27712 29257 27721 29291
rect 27721 29257 27755 29291
rect 27755 29257 27764 29291
rect 27712 29248 27764 29257
rect 28080 29248 28132 29300
rect 30748 29248 30800 29300
rect 31576 29291 31628 29300
rect 31576 29257 31585 29291
rect 31585 29257 31619 29291
rect 31619 29257 31628 29291
rect 31576 29248 31628 29257
rect 31760 29248 31812 29300
rect 32496 29248 32548 29300
rect 32956 29291 33008 29300
rect 32956 29257 32965 29291
rect 32965 29257 32999 29291
rect 32999 29257 33008 29291
rect 32956 29248 33008 29257
rect 33600 29248 33652 29300
rect 33784 29248 33836 29300
rect 23572 29223 23624 29232
rect 20904 29155 20956 29164
rect 10692 29087 10744 29096
rect 10692 29053 10701 29087
rect 10701 29053 10735 29087
rect 10735 29053 10744 29087
rect 10692 29044 10744 29053
rect 11520 29087 11572 29096
rect 11520 29053 11529 29087
rect 11529 29053 11563 29087
rect 11563 29053 11572 29087
rect 11520 29044 11572 29053
rect 8300 28976 8352 29028
rect 14464 29044 14516 29096
rect 14832 29044 14884 29096
rect 16856 29087 16908 29096
rect 16856 29053 16865 29087
rect 16865 29053 16899 29087
rect 16899 29053 16908 29087
rect 16856 29044 16908 29053
rect 11060 28908 11112 28960
rect 12164 28908 12216 28960
rect 16764 28976 16816 29028
rect 19984 29044 20036 29096
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 20904 29112 20956 29121
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 21732 29112 21784 29164
rect 23572 29189 23581 29223
rect 23581 29189 23615 29223
rect 23615 29189 23624 29223
rect 23572 29180 23624 29189
rect 25688 29180 25740 29232
rect 27436 29180 27488 29232
rect 20812 29044 20864 29096
rect 21180 29087 21232 29096
rect 21180 29053 21189 29087
rect 21189 29053 21223 29087
rect 21223 29053 21232 29087
rect 21180 29044 21232 29053
rect 25596 29112 25648 29164
rect 27804 29155 27856 29164
rect 19156 28976 19208 29028
rect 23664 29044 23716 29096
rect 27804 29121 27813 29155
rect 27813 29121 27847 29155
rect 27847 29121 27856 29155
rect 27804 29112 27856 29121
rect 34244 29223 34296 29232
rect 28356 29112 28408 29164
rect 30012 29112 30064 29164
rect 30748 29112 30800 29164
rect 31392 29155 31444 29164
rect 31392 29121 31401 29155
rect 31401 29121 31435 29155
rect 31435 29121 31444 29155
rect 31392 29112 31444 29121
rect 34244 29189 34253 29223
rect 34253 29189 34287 29223
rect 34287 29189 34296 29223
rect 34244 29180 34296 29189
rect 34796 29180 34848 29232
rect 32128 29112 32180 29164
rect 32404 29155 32456 29164
rect 32404 29121 32413 29155
rect 32413 29121 32447 29155
rect 32447 29121 32456 29155
rect 32404 29112 32456 29121
rect 33048 29112 33100 29164
rect 14832 28908 14884 28960
rect 20720 28951 20772 28960
rect 20720 28917 20729 28951
rect 20729 28917 20763 28951
rect 20763 28917 20772 28951
rect 20720 28908 20772 28917
rect 24216 28908 24268 28960
rect 24676 28908 24728 28960
rect 25964 28951 26016 28960
rect 25964 28917 25973 28951
rect 25973 28917 26007 28951
rect 26007 28917 26016 28951
rect 25964 28908 26016 28917
rect 27620 28976 27672 29028
rect 29736 29044 29788 29096
rect 29552 28951 29604 28960
rect 29552 28917 29561 28951
rect 29561 28917 29595 28951
rect 29595 28917 29604 28951
rect 29552 28908 29604 28917
rect 29644 28908 29696 28960
rect 33508 28908 33560 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 10692 28747 10744 28756
rect 10692 28713 10701 28747
rect 10701 28713 10735 28747
rect 10735 28713 10744 28747
rect 10692 28704 10744 28713
rect 12440 28747 12492 28756
rect 12440 28713 12449 28747
rect 12449 28713 12483 28747
rect 12483 28713 12492 28747
rect 12440 28704 12492 28713
rect 14464 28704 14516 28756
rect 16856 28704 16908 28756
rect 17592 28704 17644 28756
rect 20720 28704 20772 28756
rect 21732 28704 21784 28756
rect 23112 28704 23164 28756
rect 11520 28636 11572 28688
rect 20812 28636 20864 28688
rect 21272 28636 21324 28688
rect 26056 28704 26108 28756
rect 26976 28704 27028 28756
rect 27620 28704 27672 28756
rect 28908 28704 28960 28756
rect 31944 28704 31996 28756
rect 32404 28704 32456 28756
rect 34796 28747 34848 28756
rect 34796 28713 34805 28747
rect 34805 28713 34839 28747
rect 34839 28713 34848 28747
rect 34796 28704 34848 28713
rect 9956 28543 10008 28552
rect 9956 28509 9965 28543
rect 9965 28509 9999 28543
rect 9999 28509 10008 28543
rect 9956 28500 10008 28509
rect 11796 28568 11848 28620
rect 19156 28568 19208 28620
rect 21364 28568 21416 28620
rect 11244 28543 11296 28552
rect 11244 28509 11253 28543
rect 11253 28509 11287 28543
rect 11287 28509 11296 28543
rect 11244 28500 11296 28509
rect 11428 28543 11480 28552
rect 11428 28509 11437 28543
rect 11437 28509 11471 28543
rect 11471 28509 11480 28543
rect 11428 28500 11480 28509
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 14096 28543 14148 28552
rect 14096 28509 14105 28543
rect 14105 28509 14139 28543
rect 14139 28509 14148 28543
rect 14096 28500 14148 28509
rect 16580 28500 16632 28552
rect 17316 28543 17368 28552
rect 17316 28509 17325 28543
rect 17325 28509 17359 28543
rect 17359 28509 17368 28543
rect 17316 28500 17368 28509
rect 17868 28500 17920 28552
rect 18512 28543 18564 28552
rect 18512 28509 18521 28543
rect 18521 28509 18555 28543
rect 18555 28509 18564 28543
rect 18512 28500 18564 28509
rect 21732 28500 21784 28552
rect 24952 28611 25004 28620
rect 24952 28577 24961 28611
rect 24961 28577 24995 28611
rect 24995 28577 25004 28611
rect 24952 28568 25004 28577
rect 28632 28636 28684 28688
rect 29644 28636 29696 28688
rect 11980 28432 12032 28484
rect 13176 28432 13228 28484
rect 15384 28432 15436 28484
rect 19984 28432 20036 28484
rect 11336 28407 11388 28416
rect 11336 28373 11345 28407
rect 11345 28373 11379 28407
rect 11379 28373 11388 28407
rect 11336 28364 11388 28373
rect 11796 28364 11848 28416
rect 14740 28364 14792 28416
rect 19340 28364 19392 28416
rect 20352 28364 20404 28416
rect 22100 28432 22152 28484
rect 23020 28500 23072 28552
rect 24676 28543 24728 28552
rect 24676 28509 24685 28543
rect 24685 28509 24719 28543
rect 24719 28509 24728 28543
rect 24676 28500 24728 28509
rect 27068 28500 27120 28552
rect 27528 28500 27580 28552
rect 23940 28432 23992 28484
rect 25964 28432 26016 28484
rect 26976 28475 27028 28484
rect 26976 28441 26985 28475
rect 26985 28441 27019 28475
rect 27019 28441 27028 28475
rect 26976 28432 27028 28441
rect 30104 28500 30156 28552
rect 30380 28500 30432 28552
rect 31392 28568 31444 28620
rect 32128 28568 32180 28620
rect 32956 28611 33008 28620
rect 32956 28577 32965 28611
rect 32965 28577 32999 28611
rect 32999 28577 33008 28611
rect 32956 28568 33008 28577
rect 30932 28500 30984 28552
rect 30656 28432 30708 28484
rect 31668 28500 31720 28552
rect 31944 28543 31996 28552
rect 31944 28509 31953 28543
rect 31953 28509 31987 28543
rect 31987 28509 31996 28543
rect 31944 28500 31996 28509
rect 32680 28543 32732 28552
rect 32680 28509 32689 28543
rect 32689 28509 32723 28543
rect 32723 28509 32732 28543
rect 32680 28500 32732 28509
rect 34612 28500 34664 28552
rect 46940 28500 46992 28552
rect 31576 28432 31628 28484
rect 21824 28364 21876 28416
rect 23388 28364 23440 28416
rect 28632 28364 28684 28416
rect 29828 28364 29880 28416
rect 31024 28407 31076 28416
rect 31024 28373 31033 28407
rect 31033 28373 31067 28407
rect 31067 28373 31076 28407
rect 31024 28364 31076 28373
rect 32588 28364 32640 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3608 28160 3660 28212
rect 11796 28203 11848 28212
rect 3332 28024 3384 28076
rect 3608 28024 3660 28076
rect 9956 28024 10008 28076
rect 10508 27863 10560 27872
rect 10508 27829 10517 27863
rect 10517 27829 10551 27863
rect 10551 27829 10560 27863
rect 10508 27820 10560 27829
rect 11796 28169 11805 28203
rect 11805 28169 11839 28203
rect 11839 28169 11848 28203
rect 11796 28160 11848 28169
rect 13176 28203 13228 28212
rect 13176 28169 13185 28203
rect 13185 28169 13219 28203
rect 13219 28169 13228 28203
rect 13176 28160 13228 28169
rect 12164 28092 12216 28144
rect 11980 28024 12032 28076
rect 12348 28024 12400 28076
rect 13820 28092 13872 28144
rect 14464 28160 14516 28212
rect 15384 28160 15436 28212
rect 14004 28024 14056 28076
rect 11428 27956 11480 28008
rect 14832 28092 14884 28144
rect 14280 28067 14332 28076
rect 14280 28033 14289 28067
rect 14289 28033 14323 28067
rect 14323 28033 14332 28067
rect 14280 28024 14332 28033
rect 14740 28024 14792 28076
rect 15108 28067 15160 28076
rect 15108 28033 15117 28067
rect 15117 28033 15151 28067
rect 15151 28033 15160 28067
rect 15108 28024 15160 28033
rect 16580 28160 16632 28212
rect 17592 28160 17644 28212
rect 19156 28092 19208 28144
rect 27528 28203 27580 28212
rect 27528 28169 27537 28203
rect 27537 28169 27571 28203
rect 27571 28169 27580 28203
rect 27528 28160 27580 28169
rect 19340 28092 19392 28144
rect 21548 28092 21600 28144
rect 21824 28067 21876 28076
rect 21824 28033 21833 28067
rect 21833 28033 21867 28067
rect 21867 28033 21876 28067
rect 21824 28024 21876 28033
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 22836 28024 22888 28076
rect 23388 28024 23440 28076
rect 25504 28024 25556 28076
rect 26976 28067 27028 28076
rect 26976 28033 26985 28067
rect 26985 28033 27019 28067
rect 27019 28033 27028 28067
rect 26976 28024 27028 28033
rect 27068 28024 27120 28076
rect 28264 28024 28316 28076
rect 16580 27956 16632 28008
rect 11520 27931 11572 27940
rect 11520 27897 11529 27931
rect 11529 27897 11563 27931
rect 11563 27897 11572 27931
rect 11520 27888 11572 27897
rect 12624 27863 12676 27872
rect 12624 27829 12633 27863
rect 12633 27829 12667 27863
rect 12667 27829 12676 27863
rect 12624 27820 12676 27829
rect 20904 27956 20956 28008
rect 22192 27999 22244 28008
rect 22192 27965 22201 27999
rect 22201 27965 22235 27999
rect 22235 27965 22244 27999
rect 22192 27956 22244 27965
rect 28080 27956 28132 28008
rect 32036 28160 32088 28212
rect 32956 28160 33008 28212
rect 29552 28092 29604 28144
rect 30932 28092 30984 28144
rect 30840 28024 30892 28076
rect 31576 28067 31628 28076
rect 31576 28033 31585 28067
rect 31585 28033 31619 28067
rect 31619 28033 31628 28067
rect 32588 28135 32640 28144
rect 32588 28101 32597 28135
rect 32597 28101 32631 28135
rect 32631 28101 32640 28135
rect 32588 28092 32640 28101
rect 33600 28092 33652 28144
rect 32312 28067 32364 28076
rect 31576 28024 31628 28033
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 45836 28024 45888 28076
rect 29552 27956 29604 28008
rect 30380 27956 30432 28008
rect 14832 27820 14884 27872
rect 20720 27863 20772 27872
rect 20720 27829 20729 27863
rect 20729 27829 20763 27863
rect 20763 27829 20772 27863
rect 20720 27820 20772 27829
rect 27436 27820 27488 27872
rect 32128 27820 32180 27872
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 11336 27616 11388 27668
rect 11520 27616 11572 27668
rect 11888 27616 11940 27668
rect 14280 27616 14332 27668
rect 31944 27616 31996 27668
rect 42524 27616 42576 27668
rect 46204 27616 46256 27668
rect 7472 27548 7524 27600
rect 10508 27480 10560 27532
rect 14096 27548 14148 27600
rect 21364 27548 21416 27600
rect 23020 27548 23072 27600
rect 26516 27591 26568 27600
rect 26516 27557 26525 27591
rect 26525 27557 26559 27591
rect 26559 27557 26568 27591
rect 26516 27548 26568 27557
rect 29552 27591 29604 27600
rect 29552 27557 29561 27591
rect 29561 27557 29595 27591
rect 29595 27557 29604 27591
rect 29552 27548 29604 27557
rect 13912 27412 13964 27464
rect 14096 27412 14148 27464
rect 14832 27412 14884 27464
rect 20812 27455 20864 27464
rect 20812 27421 20821 27455
rect 20821 27421 20855 27455
rect 20855 27421 20864 27455
rect 20812 27412 20864 27421
rect 20996 27455 21048 27464
rect 20996 27421 21003 27455
rect 21003 27421 21048 27455
rect 20996 27412 21048 27421
rect 21916 27412 21968 27464
rect 22836 27455 22888 27464
rect 22836 27421 22845 27455
rect 22845 27421 22879 27455
rect 22879 27421 22888 27455
rect 22836 27412 22888 27421
rect 23388 27455 23440 27464
rect 12624 27344 12676 27396
rect 14004 27344 14056 27396
rect 21088 27387 21140 27396
rect 21088 27353 21097 27387
rect 21097 27353 21131 27387
rect 21131 27353 21140 27387
rect 21088 27344 21140 27353
rect 22008 27344 22060 27396
rect 23388 27421 23397 27455
rect 23397 27421 23431 27455
rect 23431 27421 23440 27455
rect 23388 27412 23440 27421
rect 23664 27344 23716 27396
rect 21272 27276 21324 27328
rect 23572 27319 23624 27328
rect 23572 27285 23581 27319
rect 23581 27285 23615 27319
rect 23615 27285 23624 27319
rect 23572 27276 23624 27285
rect 27252 27412 27304 27464
rect 31024 27548 31076 27600
rect 33600 27591 33652 27600
rect 33600 27557 33609 27591
rect 33609 27557 33643 27591
rect 33643 27557 33652 27591
rect 33600 27548 33652 27557
rect 29828 27455 29880 27464
rect 29828 27421 29837 27455
rect 29837 27421 29871 27455
rect 29871 27421 29880 27455
rect 29828 27412 29880 27421
rect 29368 27344 29420 27396
rect 45652 27480 45704 27532
rect 46940 27548 46992 27600
rect 47676 27480 47728 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 31944 27412 31996 27464
rect 31208 27344 31260 27396
rect 31668 27344 31720 27396
rect 32128 27455 32180 27464
rect 32128 27421 32137 27455
rect 32137 27421 32171 27455
rect 32171 27421 32180 27455
rect 32128 27412 32180 27421
rect 34612 27412 34664 27464
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 11244 27072 11296 27124
rect 26884 27072 26936 27124
rect 27528 27072 27580 27124
rect 11704 27004 11756 27056
rect 11520 26979 11572 26988
rect 11520 26945 11529 26979
rect 11529 26945 11563 26979
rect 11563 26945 11572 26979
rect 11520 26936 11572 26945
rect 11888 26979 11940 26988
rect 11888 26945 11897 26979
rect 11897 26945 11931 26979
rect 11931 26945 11940 26979
rect 11888 26936 11940 26945
rect 13820 26936 13872 26988
rect 15108 26936 15160 26988
rect 15292 26936 15344 26988
rect 21272 27004 21324 27056
rect 21916 27004 21968 27056
rect 23388 27004 23440 27056
rect 30656 27004 30708 27056
rect 20720 26979 20772 26988
rect 20720 26945 20729 26979
rect 20729 26945 20763 26979
rect 20763 26945 20772 26979
rect 20720 26936 20772 26945
rect 22468 26936 22520 26988
rect 24124 26979 24176 26988
rect 12164 26868 12216 26920
rect 22100 26911 22152 26920
rect 22100 26877 22109 26911
rect 22109 26877 22143 26911
rect 22143 26877 22152 26911
rect 22100 26868 22152 26877
rect 23664 26868 23716 26920
rect 14188 26775 14240 26784
rect 14188 26741 14197 26775
rect 14197 26741 14231 26775
rect 14231 26741 14240 26775
rect 14188 26732 14240 26741
rect 21180 26800 21232 26852
rect 21364 26800 21416 26852
rect 24124 26945 24133 26979
rect 24133 26945 24167 26979
rect 24167 26945 24176 26979
rect 24124 26936 24176 26945
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 28172 26979 28224 26988
rect 28172 26945 28181 26979
rect 28181 26945 28215 26979
rect 28215 26945 28224 26979
rect 28172 26936 28224 26945
rect 28908 26936 28960 26988
rect 31116 26979 31168 26988
rect 31116 26945 31125 26979
rect 31125 26945 31159 26979
rect 31159 26945 31168 26979
rect 31116 26936 31168 26945
rect 32220 26936 32272 26988
rect 25780 26911 25832 26920
rect 25780 26877 25789 26911
rect 25789 26877 25823 26911
rect 25823 26877 25832 26911
rect 25780 26868 25832 26877
rect 24400 26800 24452 26852
rect 25596 26800 25648 26852
rect 21548 26732 21600 26784
rect 23848 26732 23900 26784
rect 26240 26732 26292 26784
rect 27068 26732 27120 26784
rect 31208 26732 31260 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2044 26528 2096 26580
rect 11520 26460 11572 26512
rect 12256 26503 12308 26512
rect 12256 26469 12265 26503
rect 12265 26469 12299 26503
rect 12299 26469 12308 26503
rect 12256 26460 12308 26469
rect 14096 26460 14148 26512
rect 14004 26392 14056 26444
rect 20352 26460 20404 26512
rect 21180 26460 21232 26512
rect 21548 26503 21600 26512
rect 21548 26469 21557 26503
rect 21557 26469 21591 26503
rect 21591 26469 21600 26503
rect 21548 26460 21600 26469
rect 21732 26460 21784 26512
rect 24124 26460 24176 26512
rect 9956 26324 10008 26376
rect 11980 26324 12032 26376
rect 14096 26324 14148 26376
rect 14280 26367 14332 26376
rect 14280 26333 14289 26367
rect 14289 26333 14323 26367
rect 14323 26333 14332 26367
rect 14280 26324 14332 26333
rect 15016 26324 15068 26376
rect 16580 26367 16632 26376
rect 14740 26256 14792 26308
rect 16580 26333 16589 26367
rect 16589 26333 16623 26367
rect 16623 26333 16632 26367
rect 16580 26324 16632 26333
rect 16856 26367 16908 26376
rect 16856 26333 16865 26367
rect 16865 26333 16899 26367
rect 16899 26333 16908 26367
rect 16856 26324 16908 26333
rect 16948 26324 17000 26376
rect 20904 26392 20956 26444
rect 21364 26392 21416 26444
rect 22560 26392 22612 26444
rect 23388 26435 23440 26444
rect 23388 26401 23397 26435
rect 23397 26401 23431 26435
rect 23431 26401 23440 26435
rect 23388 26392 23440 26401
rect 19984 26324 20036 26376
rect 21548 26324 21600 26376
rect 24400 26367 24452 26376
rect 18880 26256 18932 26308
rect 20352 26256 20404 26308
rect 20996 26256 21048 26308
rect 21272 26299 21324 26308
rect 10232 26231 10284 26240
rect 10232 26197 10241 26231
rect 10241 26197 10275 26231
rect 10275 26197 10284 26231
rect 10232 26188 10284 26197
rect 13820 26188 13872 26240
rect 16672 26188 16724 26240
rect 17132 26188 17184 26240
rect 18144 26231 18196 26240
rect 18144 26197 18153 26231
rect 18153 26197 18187 26231
rect 18187 26197 18196 26231
rect 18144 26188 18196 26197
rect 21272 26265 21281 26299
rect 21281 26265 21315 26299
rect 21315 26265 21324 26299
rect 21272 26256 21324 26265
rect 21732 26256 21784 26308
rect 21824 26256 21876 26308
rect 24400 26333 24409 26367
rect 24409 26333 24443 26367
rect 24443 26333 24452 26367
rect 24400 26324 24452 26333
rect 25688 26392 25740 26444
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 26516 26460 26568 26512
rect 27528 26392 27580 26444
rect 26516 26367 26568 26376
rect 26516 26333 26525 26367
rect 26525 26333 26559 26367
rect 26559 26333 26568 26367
rect 27068 26367 27120 26376
rect 26516 26324 26568 26333
rect 27068 26333 27077 26367
rect 27077 26333 27111 26367
rect 27111 26333 27120 26367
rect 27068 26324 27120 26333
rect 27252 26324 27304 26376
rect 28908 26528 28960 26580
rect 32680 26571 32732 26580
rect 23664 26256 23716 26308
rect 26976 26256 27028 26308
rect 28264 26256 28316 26308
rect 30380 26392 30432 26444
rect 29184 26324 29236 26376
rect 29552 26256 29604 26308
rect 30840 26299 30892 26308
rect 30840 26265 30849 26299
rect 30849 26265 30883 26299
rect 30883 26265 30892 26299
rect 30840 26256 30892 26265
rect 32680 26537 32689 26571
rect 32689 26537 32723 26571
rect 32723 26537 32732 26571
rect 32680 26528 32732 26537
rect 32772 26528 32824 26580
rect 33508 26528 33560 26580
rect 33968 26460 34020 26512
rect 32588 26392 32640 26444
rect 33692 26392 33744 26444
rect 31760 26324 31812 26376
rect 32036 26367 32088 26376
rect 32036 26333 32045 26367
rect 32045 26333 32079 26367
rect 32079 26333 32088 26367
rect 32036 26324 32088 26333
rect 33784 26367 33836 26376
rect 33784 26333 33793 26367
rect 33793 26333 33827 26367
rect 33827 26333 33836 26367
rect 33784 26324 33836 26333
rect 31944 26299 31996 26308
rect 31944 26265 31953 26299
rect 31953 26265 31987 26299
rect 31987 26265 31996 26299
rect 31944 26256 31996 26265
rect 32128 26256 32180 26308
rect 33048 26256 33100 26308
rect 46388 26324 46440 26376
rect 23020 26188 23072 26240
rect 26240 26188 26292 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 12256 25984 12308 26036
rect 18880 26027 18932 26036
rect 11796 25848 11848 25900
rect 10968 25780 11020 25832
rect 13820 25916 13872 25968
rect 14188 25916 14240 25968
rect 18880 25993 18889 26027
rect 18889 25993 18923 26027
rect 18923 25993 18932 26027
rect 18880 25984 18932 25993
rect 20812 25984 20864 26036
rect 16580 25916 16632 25968
rect 19984 25916 20036 25968
rect 20628 25916 20680 25968
rect 16856 25848 16908 25900
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 19340 25848 19392 25900
rect 20352 25848 20404 25900
rect 20720 25891 20772 25900
rect 20720 25857 20729 25891
rect 20729 25857 20763 25891
rect 20763 25857 20772 25891
rect 20720 25848 20772 25857
rect 20904 25891 20956 25900
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 21180 25891 21232 25900
rect 21180 25857 21189 25891
rect 21189 25857 21223 25891
rect 21223 25857 21232 25891
rect 21180 25848 21232 25857
rect 13912 25780 13964 25832
rect 14924 25780 14976 25832
rect 15660 25823 15712 25832
rect 15660 25789 15669 25823
rect 15669 25789 15703 25823
rect 15703 25789 15712 25823
rect 15660 25780 15712 25789
rect 18144 25780 18196 25832
rect 19524 25823 19576 25832
rect 19524 25789 19533 25823
rect 19533 25789 19567 25823
rect 19567 25789 19576 25823
rect 19524 25780 19576 25789
rect 21548 25780 21600 25832
rect 21272 25712 21324 25764
rect 24492 25916 24544 25968
rect 30840 25984 30892 26036
rect 31116 25984 31168 26036
rect 32220 26027 32272 26036
rect 25780 25891 25832 25900
rect 25780 25857 25789 25891
rect 25789 25857 25823 25891
rect 25823 25857 25832 25891
rect 25780 25848 25832 25857
rect 26516 25848 26568 25900
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 29552 25916 29604 25968
rect 32220 25993 32229 26027
rect 32229 25993 32263 26027
rect 32263 25993 32272 26027
rect 32220 25984 32272 25993
rect 27712 25848 27764 25900
rect 28632 25891 28684 25900
rect 28632 25857 28641 25891
rect 28641 25857 28675 25891
rect 28675 25857 28684 25891
rect 28632 25848 28684 25857
rect 10508 25644 10560 25696
rect 14096 25644 14148 25696
rect 14280 25644 14332 25696
rect 15108 25644 15160 25696
rect 16948 25644 17000 25696
rect 23572 25780 23624 25832
rect 23664 25780 23716 25832
rect 24032 25712 24084 25764
rect 26240 25823 26292 25832
rect 26240 25789 26274 25823
rect 26274 25789 26292 25823
rect 26240 25780 26292 25789
rect 27436 25780 27488 25832
rect 29920 25848 29972 25900
rect 33048 25916 33100 25968
rect 30472 25848 30524 25900
rect 31392 25891 31444 25900
rect 31392 25857 31401 25891
rect 31401 25857 31435 25891
rect 31435 25857 31444 25891
rect 31392 25848 31444 25857
rect 32128 25891 32180 25900
rect 32128 25857 32137 25891
rect 32137 25857 32171 25891
rect 32171 25857 32180 25891
rect 32128 25848 32180 25857
rect 32588 25848 32640 25900
rect 32680 25848 32732 25900
rect 33692 25848 33744 25900
rect 33968 25891 34020 25900
rect 33968 25857 33977 25891
rect 33977 25857 34011 25891
rect 34011 25857 34020 25891
rect 33968 25848 34020 25857
rect 33048 25823 33100 25832
rect 33048 25789 33057 25823
rect 33057 25789 33091 25823
rect 33091 25789 33100 25823
rect 33048 25780 33100 25789
rect 23480 25644 23532 25696
rect 24860 25644 24912 25696
rect 28172 25712 28224 25764
rect 31668 25712 31720 25764
rect 32220 25712 32272 25764
rect 32496 25712 32548 25764
rect 26884 25644 26936 25696
rect 29552 25644 29604 25696
rect 33324 25644 33376 25696
rect 46296 25644 46348 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 15568 25440 15620 25492
rect 17408 25440 17460 25492
rect 19340 25483 19392 25492
rect 19340 25449 19349 25483
rect 19349 25449 19383 25483
rect 19383 25449 19392 25483
rect 19340 25440 19392 25449
rect 23020 25483 23072 25492
rect 23020 25449 23029 25483
rect 23029 25449 23063 25483
rect 23063 25449 23072 25483
rect 23020 25440 23072 25449
rect 24492 25483 24544 25492
rect 24492 25449 24501 25483
rect 24501 25449 24535 25483
rect 24535 25449 24544 25483
rect 24492 25440 24544 25449
rect 21548 25372 21600 25424
rect 21916 25372 21968 25424
rect 22836 25372 22888 25424
rect 10232 25347 10284 25356
rect 10232 25313 10241 25347
rect 10241 25313 10275 25347
rect 10275 25313 10284 25347
rect 10232 25304 10284 25313
rect 10508 25347 10560 25356
rect 10508 25313 10517 25347
rect 10517 25313 10551 25347
rect 10551 25313 10560 25347
rect 10508 25304 10560 25313
rect 11796 25304 11848 25356
rect 15476 25304 15528 25356
rect 16948 25347 17000 25356
rect 11612 25236 11664 25288
rect 14740 25279 14792 25288
rect 14740 25245 14749 25279
rect 14749 25245 14783 25279
rect 14783 25245 14792 25279
rect 14740 25236 14792 25245
rect 14832 25236 14884 25288
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 14096 25168 14148 25220
rect 15016 25168 15068 25220
rect 15108 25168 15160 25220
rect 2044 25100 2096 25152
rect 14832 25100 14884 25152
rect 15200 25100 15252 25152
rect 16948 25313 16957 25347
rect 16957 25313 16991 25347
rect 16991 25313 17000 25347
rect 16948 25304 17000 25313
rect 19524 25304 19576 25356
rect 24860 25304 24912 25356
rect 16672 25279 16724 25288
rect 16672 25245 16681 25279
rect 16681 25245 16715 25279
rect 16715 25245 16724 25279
rect 16672 25236 16724 25245
rect 18236 25236 18288 25288
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 15844 25100 15896 25152
rect 16580 25100 16632 25152
rect 17040 25100 17092 25152
rect 18328 25168 18380 25220
rect 21272 25279 21324 25288
rect 21272 25245 21282 25279
rect 21282 25245 21316 25279
rect 21316 25245 21324 25279
rect 21548 25279 21600 25288
rect 21272 25236 21324 25245
rect 21548 25245 21557 25279
rect 21557 25245 21591 25279
rect 21591 25245 21600 25279
rect 21548 25236 21600 25245
rect 22008 25236 22060 25288
rect 23112 25236 23164 25288
rect 23848 25236 23900 25288
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 21088 25168 21140 25220
rect 26240 25372 26292 25424
rect 29276 25372 29328 25424
rect 33692 25440 33744 25492
rect 32220 25372 32272 25424
rect 25872 25304 25924 25356
rect 28632 25304 28684 25356
rect 25596 25279 25648 25288
rect 25596 25245 25605 25279
rect 25605 25245 25639 25279
rect 25639 25245 25648 25279
rect 25596 25236 25648 25245
rect 25780 25279 25832 25288
rect 25780 25245 25789 25279
rect 25789 25245 25823 25279
rect 25823 25245 25832 25279
rect 25780 25236 25832 25245
rect 26608 25279 26660 25288
rect 26608 25245 26617 25279
rect 26617 25245 26651 25279
rect 26651 25245 26660 25279
rect 26608 25236 26660 25245
rect 26884 25279 26936 25288
rect 26884 25245 26893 25279
rect 26893 25245 26927 25279
rect 26927 25245 26936 25279
rect 26884 25236 26936 25245
rect 26976 25279 27028 25288
rect 26976 25245 26985 25279
rect 26985 25245 27019 25279
rect 27019 25245 27028 25279
rect 29552 25279 29604 25288
rect 26976 25236 27028 25245
rect 29552 25245 29561 25279
rect 29561 25245 29595 25279
rect 29595 25245 29604 25279
rect 29552 25236 29604 25245
rect 31392 25304 31444 25356
rect 31116 25279 31168 25288
rect 31116 25245 31125 25279
rect 31125 25245 31159 25279
rect 31159 25245 31168 25279
rect 31116 25236 31168 25245
rect 27528 25168 27580 25220
rect 32312 25304 32364 25356
rect 33324 25304 33376 25356
rect 46296 25347 46348 25356
rect 46296 25313 46305 25347
rect 46305 25313 46339 25347
rect 46339 25313 46348 25347
rect 46296 25304 46348 25313
rect 22100 25100 22152 25152
rect 25412 25100 25464 25152
rect 26240 25100 26292 25152
rect 30840 25100 30892 25152
rect 32588 25168 32640 25220
rect 33140 25168 33192 25220
rect 35164 25211 35216 25220
rect 35164 25177 35173 25211
rect 35173 25177 35207 25211
rect 35207 25177 35216 25211
rect 35164 25168 35216 25177
rect 47676 25168 47728 25220
rect 48136 25211 48188 25220
rect 48136 25177 48145 25211
rect 48145 25177 48179 25211
rect 48179 25177 48188 25211
rect 48136 25168 48188 25177
rect 31300 25143 31352 25152
rect 31300 25109 31309 25143
rect 31309 25109 31343 25143
rect 31343 25109 31352 25143
rect 31300 25100 31352 25109
rect 34796 25100 34848 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 14740 24896 14792 24948
rect 15660 24896 15712 24948
rect 17040 24939 17092 24948
rect 17040 24905 17049 24939
rect 17049 24905 17083 24939
rect 17083 24905 17092 24939
rect 17040 24896 17092 24905
rect 21272 24939 21324 24948
rect 21272 24905 21281 24939
rect 21281 24905 21315 24939
rect 21315 24905 21324 24939
rect 21272 24896 21324 24905
rect 10968 24803 11020 24812
rect 10968 24769 10977 24803
rect 10977 24769 11011 24803
rect 11011 24769 11020 24803
rect 10968 24760 11020 24769
rect 11336 24692 11388 24744
rect 11612 24803 11664 24812
rect 11612 24769 11621 24803
rect 11621 24769 11655 24803
rect 11655 24769 11664 24803
rect 11612 24760 11664 24769
rect 16948 24871 17000 24880
rect 16948 24837 16957 24871
rect 16957 24837 16991 24871
rect 16991 24837 17000 24871
rect 23480 24896 23532 24948
rect 24676 24896 24728 24948
rect 25044 24896 25096 24948
rect 25780 24896 25832 24948
rect 26516 24896 26568 24948
rect 16948 24828 17000 24837
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 15568 24760 15620 24812
rect 15844 24803 15896 24812
rect 15844 24769 15853 24803
rect 15853 24769 15887 24803
rect 15887 24769 15896 24803
rect 15844 24760 15896 24769
rect 12348 24692 12400 24744
rect 14556 24735 14608 24744
rect 14556 24701 14565 24735
rect 14565 24701 14599 24735
rect 14599 24701 14608 24735
rect 14556 24692 14608 24701
rect 15200 24692 15252 24744
rect 16764 24760 16816 24812
rect 18236 24803 18288 24812
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 18328 24803 18380 24812
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 21548 24760 21600 24812
rect 31300 24828 31352 24880
rect 34796 24828 34848 24880
rect 23204 24760 23256 24812
rect 26976 24803 27028 24812
rect 20720 24692 20772 24744
rect 20996 24735 21048 24744
rect 20996 24701 21005 24735
rect 21005 24701 21039 24735
rect 21039 24701 21048 24735
rect 20996 24692 21048 24701
rect 22100 24735 22152 24744
rect 22100 24701 22109 24735
rect 22109 24701 22143 24735
rect 22143 24701 22152 24735
rect 24676 24735 24728 24744
rect 22100 24692 22152 24701
rect 24676 24701 24685 24735
rect 24685 24701 24719 24735
rect 24719 24701 24728 24735
rect 24676 24692 24728 24701
rect 26976 24769 26985 24803
rect 26985 24769 27019 24803
rect 27019 24769 27028 24803
rect 26976 24760 27028 24769
rect 28080 24803 28132 24812
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 28080 24760 28132 24769
rect 29644 24760 29696 24812
rect 31208 24803 31260 24812
rect 28356 24735 28408 24744
rect 28356 24701 28365 24735
rect 28365 24701 28399 24735
rect 28399 24701 28408 24735
rect 28356 24692 28408 24701
rect 30380 24692 30432 24744
rect 31208 24769 31217 24803
rect 31217 24769 31251 24803
rect 31251 24769 31260 24803
rect 31208 24760 31260 24769
rect 32220 24803 32272 24812
rect 32220 24769 32229 24803
rect 32229 24769 32263 24803
rect 32263 24769 32272 24803
rect 32220 24760 32272 24769
rect 32404 24803 32456 24812
rect 32404 24769 32413 24803
rect 32413 24769 32447 24803
rect 32447 24769 32456 24803
rect 32404 24760 32456 24769
rect 32496 24760 32548 24812
rect 33140 24760 33192 24812
rect 35164 24803 35216 24812
rect 35164 24769 35173 24803
rect 35173 24769 35207 24803
rect 35207 24769 35216 24803
rect 35164 24760 35216 24769
rect 45008 24760 45060 24812
rect 47584 24803 47636 24812
rect 47584 24769 47593 24803
rect 47593 24769 47627 24803
rect 47627 24769 47636 24803
rect 47584 24760 47636 24769
rect 47676 24803 47728 24812
rect 47676 24769 47685 24803
rect 47685 24769 47719 24803
rect 47719 24769 47728 24803
rect 47676 24760 47728 24769
rect 32128 24692 32180 24744
rect 44364 24692 44416 24744
rect 45100 24692 45152 24744
rect 45376 24735 45428 24744
rect 45376 24701 45385 24735
rect 45385 24701 45419 24735
rect 45419 24701 45428 24735
rect 45376 24692 45428 24701
rect 46756 24735 46808 24744
rect 46756 24701 46765 24735
rect 46765 24701 46799 24735
rect 46799 24701 46808 24735
rect 46756 24692 46808 24701
rect 26240 24624 26292 24676
rect 10600 24556 10652 24608
rect 21916 24556 21968 24608
rect 27344 24556 27396 24608
rect 46848 24624 46900 24676
rect 30380 24599 30432 24608
rect 30380 24565 30389 24599
rect 30389 24565 30423 24599
rect 30423 24565 30432 24599
rect 30380 24556 30432 24565
rect 30656 24556 30708 24608
rect 32128 24556 32180 24608
rect 32220 24556 32272 24608
rect 34796 24556 34848 24608
rect 40040 24599 40092 24608
rect 40040 24565 40049 24599
rect 40049 24565 40083 24599
rect 40083 24565 40092 24599
rect 40040 24556 40092 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 16672 24352 16724 24404
rect 19340 24352 19392 24404
rect 23112 24352 23164 24404
rect 23204 24352 23256 24404
rect 26056 24352 26108 24404
rect 10600 24259 10652 24268
rect 10600 24225 10609 24259
rect 10609 24225 10643 24259
rect 10643 24225 10652 24259
rect 10600 24216 10652 24225
rect 10324 24191 10376 24200
rect 10324 24157 10333 24191
rect 10333 24157 10367 24191
rect 10367 24157 10376 24191
rect 10324 24148 10376 24157
rect 12348 24148 12400 24200
rect 14924 24148 14976 24200
rect 16856 24148 16908 24200
rect 20536 24284 20588 24336
rect 27160 24352 27212 24404
rect 29644 24395 29696 24404
rect 29644 24361 29653 24395
rect 29653 24361 29687 24395
rect 29687 24361 29696 24395
rect 29644 24352 29696 24361
rect 30380 24352 30432 24404
rect 32588 24352 32640 24404
rect 45376 24352 45428 24404
rect 30656 24284 30708 24336
rect 17776 24216 17828 24268
rect 19064 24148 19116 24200
rect 24676 24216 24728 24268
rect 25412 24259 25464 24268
rect 25412 24225 25421 24259
rect 25421 24225 25455 24259
rect 25455 24225 25464 24259
rect 25412 24216 25464 24225
rect 32312 24216 32364 24268
rect 35348 24216 35400 24268
rect 45652 24284 45704 24336
rect 40040 24259 40092 24268
rect 40040 24225 40049 24259
rect 40049 24225 40083 24259
rect 40083 24225 40092 24259
rect 40040 24216 40092 24225
rect 40316 24259 40368 24268
rect 40316 24225 40325 24259
rect 40325 24225 40359 24259
rect 40359 24225 40368 24259
rect 40316 24216 40368 24225
rect 44364 24216 44416 24268
rect 22836 24148 22888 24200
rect 24400 24148 24452 24200
rect 28632 24148 28684 24200
rect 32128 24148 32180 24200
rect 34612 24148 34664 24200
rect 45008 24191 45060 24200
rect 11888 24012 11940 24064
rect 14372 24012 14424 24064
rect 17684 24012 17736 24064
rect 17868 24055 17920 24064
rect 17868 24021 17877 24055
rect 17877 24021 17911 24055
rect 17911 24021 17920 24055
rect 17868 24012 17920 24021
rect 20076 24055 20128 24064
rect 20076 24021 20085 24055
rect 20085 24021 20119 24055
rect 20119 24021 20128 24055
rect 20076 24012 20128 24021
rect 25964 24080 26016 24132
rect 34520 24080 34572 24132
rect 45008 24157 45017 24191
rect 45017 24157 45051 24191
rect 45051 24157 45060 24191
rect 45008 24148 45060 24157
rect 46480 24216 46532 24268
rect 45836 24148 45888 24200
rect 46296 24191 46348 24200
rect 46296 24157 46305 24191
rect 46305 24157 46339 24191
rect 46339 24157 46348 24191
rect 46296 24148 46348 24157
rect 40040 24080 40092 24132
rect 41052 24080 41104 24132
rect 47768 24012 47820 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3516 23808 3568 23860
rect 17592 23851 17644 23860
rect 3884 23740 3936 23792
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 9956 23672 10008 23724
rect 10324 23740 10376 23792
rect 11796 23647 11848 23656
rect 11796 23613 11805 23647
rect 11805 23613 11839 23647
rect 11839 23613 11848 23647
rect 11796 23604 11848 23613
rect 11980 23647 12032 23656
rect 11980 23613 11989 23647
rect 11989 23613 12023 23647
rect 12023 23613 12032 23647
rect 11980 23604 12032 23613
rect 14372 23740 14424 23792
rect 17592 23817 17601 23851
rect 17601 23817 17635 23851
rect 17635 23817 17644 23851
rect 17592 23808 17644 23817
rect 17684 23808 17736 23860
rect 19340 23808 19392 23860
rect 23480 23808 23532 23860
rect 24400 23808 24452 23860
rect 25964 23851 26016 23860
rect 25964 23817 25973 23851
rect 25973 23817 26007 23851
rect 26007 23817 26016 23851
rect 25964 23808 26016 23817
rect 32128 23808 32180 23860
rect 34520 23851 34572 23860
rect 34520 23817 34529 23851
rect 34529 23817 34563 23851
rect 34563 23817 34572 23851
rect 34520 23808 34572 23817
rect 41052 23851 41104 23860
rect 41052 23817 41061 23851
rect 41061 23817 41095 23851
rect 41095 23817 41104 23851
rect 41052 23808 41104 23817
rect 20076 23740 20128 23792
rect 26792 23740 26844 23792
rect 40316 23740 40368 23792
rect 14924 23715 14976 23724
rect 14924 23681 14933 23715
rect 14933 23681 14967 23715
rect 14967 23681 14976 23715
rect 14924 23672 14976 23681
rect 15292 23672 15344 23724
rect 17960 23672 18012 23724
rect 19340 23672 19392 23724
rect 23112 23672 23164 23724
rect 24400 23672 24452 23724
rect 26976 23672 27028 23724
rect 28632 23672 28684 23724
rect 32496 23672 32548 23724
rect 35348 23672 35400 23724
rect 39672 23715 39724 23724
rect 39672 23681 39681 23715
rect 39681 23681 39715 23715
rect 39715 23681 39724 23715
rect 39672 23672 39724 23681
rect 47492 23740 47544 23792
rect 13912 23604 13964 23656
rect 16396 23604 16448 23656
rect 19064 23604 19116 23656
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 13820 23468 13872 23520
rect 14924 23468 14976 23520
rect 17132 23468 17184 23520
rect 19340 23468 19392 23520
rect 27160 23536 27212 23588
rect 35992 23536 36044 23588
rect 39396 23604 39448 23656
rect 42616 23672 42668 23724
rect 43260 23715 43312 23724
rect 43260 23681 43269 23715
rect 43269 23681 43303 23715
rect 43303 23681 43312 23715
rect 43260 23672 43312 23681
rect 43904 23672 43956 23724
rect 44088 23715 44140 23724
rect 44088 23681 44097 23715
rect 44097 23681 44131 23715
rect 44131 23681 44140 23715
rect 44088 23672 44140 23681
rect 45744 23715 45796 23724
rect 45744 23681 45753 23715
rect 45753 23681 45787 23715
rect 45787 23681 45796 23715
rect 45744 23672 45796 23681
rect 47032 23672 47084 23724
rect 46204 23647 46256 23656
rect 46204 23613 46213 23647
rect 46213 23613 46247 23647
rect 46247 23613 46256 23647
rect 46204 23604 46256 23613
rect 45652 23536 45704 23588
rect 24584 23468 24636 23520
rect 43812 23468 43864 23520
rect 46940 23468 46992 23520
rect 47676 23511 47728 23520
rect 47676 23477 47685 23511
rect 47685 23477 47719 23511
rect 47719 23477 47728 23511
rect 47676 23468 47728 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 11336 23307 11388 23316
rect 11336 23273 11345 23307
rect 11345 23273 11379 23307
rect 11379 23273 11388 23307
rect 11336 23264 11388 23273
rect 11980 23264 12032 23316
rect 12256 23264 12308 23316
rect 14556 23264 14608 23316
rect 14740 23264 14792 23316
rect 16856 23264 16908 23316
rect 19248 23264 19300 23316
rect 21824 23264 21876 23316
rect 22008 23264 22060 23316
rect 22560 23264 22612 23316
rect 22652 23264 22704 23316
rect 25872 23264 25924 23316
rect 35716 23264 35768 23316
rect 42340 23264 42392 23316
rect 3608 23128 3660 23180
rect 14096 23171 14148 23180
rect 14096 23137 14105 23171
rect 14105 23137 14139 23171
rect 14139 23137 14148 23171
rect 14096 23128 14148 23137
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 16396 23171 16448 23180
rect 16396 23137 16405 23171
rect 16405 23137 16439 23171
rect 16439 23137 16448 23171
rect 16396 23128 16448 23137
rect 19340 23196 19392 23248
rect 20536 23196 20588 23248
rect 35716 23171 35768 23180
rect 35716 23137 35725 23171
rect 35725 23137 35759 23171
rect 35759 23137 35768 23171
rect 35716 23128 35768 23137
rect 40500 23171 40552 23180
rect 40500 23137 40509 23171
rect 40509 23137 40543 23171
rect 40543 23137 40552 23171
rect 40500 23128 40552 23137
rect 9956 23060 10008 23112
rect 11060 23060 11112 23112
rect 11612 23103 11664 23112
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 11796 22992 11848 23044
rect 9864 22967 9916 22976
rect 9864 22933 9873 22967
rect 9873 22933 9907 22967
rect 9907 22933 9916 22967
rect 9864 22924 9916 22933
rect 10784 22967 10836 22976
rect 10784 22933 10793 22967
rect 10793 22933 10827 22967
rect 10827 22933 10836 22967
rect 10784 22924 10836 22933
rect 12256 22924 12308 22976
rect 13084 22967 13136 22976
rect 13084 22933 13109 22967
rect 13109 22933 13136 22967
rect 19340 23103 19392 23112
rect 19340 23069 19349 23103
rect 19349 23069 19383 23103
rect 19383 23069 19392 23103
rect 19340 23060 19392 23069
rect 20076 23060 20128 23112
rect 21364 23060 21416 23112
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 23480 23103 23532 23112
rect 23480 23069 23489 23103
rect 23489 23069 23523 23103
rect 23523 23069 23532 23103
rect 23480 23060 23532 23069
rect 25504 23103 25556 23112
rect 25504 23069 25513 23103
rect 25513 23069 25547 23103
rect 25547 23069 25556 23103
rect 25504 23060 25556 23069
rect 28264 23103 28316 23112
rect 28264 23069 28273 23103
rect 28273 23069 28307 23103
rect 28307 23069 28316 23103
rect 28264 23060 28316 23069
rect 30196 23103 30248 23112
rect 30196 23069 30205 23103
rect 30205 23069 30239 23103
rect 30239 23069 30248 23103
rect 30196 23060 30248 23069
rect 33140 23060 33192 23112
rect 14280 23035 14332 23044
rect 14280 23001 14289 23035
rect 14289 23001 14323 23035
rect 14323 23001 14332 23035
rect 14280 22992 14332 23001
rect 14464 22992 14516 23044
rect 15292 22992 15344 23044
rect 15476 22992 15528 23044
rect 17132 22992 17184 23044
rect 18420 22992 18472 23044
rect 20720 22992 20772 23044
rect 22560 22992 22612 23044
rect 32220 22992 32272 23044
rect 13084 22924 13136 22933
rect 16580 22924 16632 22976
rect 16856 22924 16908 22976
rect 22928 22967 22980 22976
rect 22928 22933 22937 22967
rect 22937 22933 22971 22967
rect 22971 22933 22980 22967
rect 22928 22924 22980 22933
rect 23388 22924 23440 22976
rect 28724 22924 28776 22976
rect 33784 22967 33836 22976
rect 33784 22933 33793 22967
rect 33793 22933 33827 22967
rect 33827 22933 33836 22967
rect 33784 22924 33836 22933
rect 35348 23060 35400 23112
rect 39856 23103 39908 23112
rect 39856 23069 39865 23103
rect 39865 23069 39899 23103
rect 39899 23069 39908 23103
rect 39856 23060 39908 23069
rect 42432 23060 42484 23112
rect 39488 22992 39540 23044
rect 39580 22924 39632 22976
rect 45928 23196 45980 23248
rect 46388 23196 46440 23248
rect 43628 23171 43680 23180
rect 43628 23137 43637 23171
rect 43637 23137 43671 23171
rect 43671 23137 43680 23171
rect 43628 23128 43680 23137
rect 47676 23128 47728 23180
rect 48228 23128 48280 23180
rect 43812 23103 43864 23112
rect 43812 23069 43821 23103
rect 43821 23069 43855 23103
rect 43855 23069 43864 23103
rect 43812 23060 43864 23069
rect 45560 22992 45612 23044
rect 45376 22924 45428 22976
rect 47768 22992 47820 23044
rect 46296 22924 46348 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9956 22720 10008 22772
rect 11888 22763 11940 22772
rect 11888 22729 11897 22763
rect 11897 22729 11931 22763
rect 11931 22729 11940 22763
rect 11888 22720 11940 22729
rect 12256 22720 12308 22772
rect 11244 22652 11296 22704
rect 12164 22652 12216 22704
rect 14740 22720 14792 22772
rect 11336 22584 11388 22636
rect 13820 22584 13872 22636
rect 14464 22652 14516 22704
rect 22008 22720 22060 22772
rect 32220 22763 32272 22772
rect 22928 22652 22980 22704
rect 15844 22584 15896 22636
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 21824 22627 21876 22636
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 28264 22652 28316 22704
rect 29644 22652 29696 22704
rect 32220 22729 32229 22763
rect 32229 22729 32263 22763
rect 32263 22729 32272 22763
rect 32220 22720 32272 22729
rect 37280 22720 37332 22772
rect 39488 22763 39540 22772
rect 39488 22729 39497 22763
rect 39497 22729 39531 22763
rect 39531 22729 39540 22763
rect 39488 22720 39540 22729
rect 33784 22695 33836 22704
rect 33784 22661 33793 22695
rect 33793 22661 33827 22695
rect 33827 22661 33836 22695
rect 33784 22652 33836 22661
rect 43996 22652 44048 22704
rect 45376 22695 45428 22704
rect 45376 22661 45385 22695
rect 45385 22661 45419 22695
rect 45419 22661 45428 22695
rect 45376 22652 45428 22661
rect 8392 22559 8444 22568
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 15200 22559 15252 22568
rect 3700 22448 3752 22500
rect 15200 22525 15209 22559
rect 15209 22525 15243 22559
rect 15243 22525 15252 22559
rect 15200 22516 15252 22525
rect 15476 22559 15528 22568
rect 15476 22525 15485 22559
rect 15485 22525 15519 22559
rect 15519 22525 15528 22559
rect 15476 22516 15528 22525
rect 17040 22559 17092 22568
rect 17040 22525 17049 22559
rect 17049 22525 17083 22559
rect 17083 22525 17092 22559
rect 17040 22516 17092 22525
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 11060 22448 11112 22500
rect 13084 22448 13136 22500
rect 11704 22423 11756 22432
rect 11704 22389 11713 22423
rect 11713 22389 11747 22423
rect 11747 22389 11756 22423
rect 11704 22380 11756 22389
rect 11980 22380 12032 22432
rect 12348 22380 12400 22432
rect 15660 22448 15712 22500
rect 19984 22516 20036 22568
rect 21272 22559 21324 22568
rect 21272 22525 21281 22559
rect 21281 22525 21315 22559
rect 21315 22525 21324 22559
rect 21272 22516 21324 22525
rect 23296 22559 23348 22568
rect 23296 22525 23305 22559
rect 23305 22525 23339 22559
rect 23339 22525 23348 22559
rect 23296 22516 23348 22525
rect 23112 22448 23164 22500
rect 27344 22584 27396 22636
rect 28724 22627 28776 22636
rect 27988 22559 28040 22568
rect 27988 22525 27997 22559
rect 27997 22525 28031 22559
rect 28031 22525 28040 22559
rect 27988 22516 28040 22525
rect 14464 22423 14516 22432
rect 14464 22389 14473 22423
rect 14473 22389 14507 22423
rect 14507 22389 14516 22423
rect 14464 22380 14516 22389
rect 19340 22380 19392 22432
rect 25964 22423 26016 22432
rect 25964 22389 25973 22423
rect 25973 22389 26007 22423
rect 26007 22389 26016 22423
rect 25964 22380 26016 22389
rect 27068 22380 27120 22432
rect 28724 22593 28733 22627
rect 28733 22593 28767 22627
rect 28767 22593 28776 22627
rect 28724 22584 28776 22593
rect 33140 22584 33192 22636
rect 39580 22584 39632 22636
rect 40040 22627 40092 22636
rect 40040 22593 40049 22627
rect 40049 22593 40083 22627
rect 40083 22593 40092 22627
rect 40040 22584 40092 22593
rect 42432 22627 42484 22636
rect 42432 22593 42441 22627
rect 42441 22593 42475 22627
rect 42475 22593 42484 22627
rect 42432 22584 42484 22593
rect 43536 22627 43588 22636
rect 43536 22593 43545 22627
rect 43545 22593 43579 22627
rect 43579 22593 43588 22627
rect 43536 22584 43588 22593
rect 43628 22627 43680 22636
rect 43628 22593 43637 22627
rect 43637 22593 43671 22627
rect 43671 22593 43680 22627
rect 43628 22584 43680 22593
rect 43904 22584 43956 22636
rect 44272 22627 44324 22636
rect 44272 22593 44281 22627
rect 44281 22593 44315 22627
rect 44315 22593 44324 22627
rect 44272 22584 44324 22593
rect 29092 22516 29144 22568
rect 40224 22559 40276 22568
rect 40224 22525 40233 22559
rect 40233 22525 40267 22559
rect 40267 22525 40276 22559
rect 40224 22516 40276 22525
rect 42524 22448 42576 22500
rect 42616 22448 42668 22500
rect 44088 22491 44140 22500
rect 44088 22457 44097 22491
rect 44097 22457 44131 22491
rect 44131 22457 44140 22491
rect 44088 22448 44140 22457
rect 45560 22516 45612 22568
rect 47676 22720 47728 22772
rect 46940 22652 46992 22704
rect 47124 22584 47176 22636
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 47860 22627 47912 22636
rect 47860 22593 47869 22627
rect 47869 22593 47903 22627
rect 47903 22593 47912 22627
rect 47860 22584 47912 22593
rect 47216 22516 47268 22568
rect 47492 22448 47544 22500
rect 30196 22380 30248 22432
rect 43260 22380 43312 22432
rect 44272 22380 44324 22432
rect 48136 22423 48188 22432
rect 48136 22389 48145 22423
rect 48145 22389 48179 22423
rect 48179 22389 48188 22423
rect 48136 22380 48188 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 8392 22176 8444 22228
rect 14280 22176 14332 22228
rect 16580 22176 16632 22228
rect 18236 22176 18288 22228
rect 20628 22176 20680 22228
rect 21272 22176 21324 22228
rect 39856 22176 39908 22228
rect 40132 22219 40184 22228
rect 40132 22185 40141 22219
rect 40141 22185 40175 22219
rect 40175 22185 40184 22219
rect 40132 22176 40184 22185
rect 40224 22176 40276 22228
rect 43536 22176 43588 22228
rect 44456 22176 44508 22228
rect 48044 22176 48096 22228
rect 11244 22151 11296 22160
rect 11244 22117 11253 22151
rect 11253 22117 11287 22151
rect 11287 22117 11296 22151
rect 11244 22108 11296 22117
rect 14924 22108 14976 22160
rect 20076 22108 20128 22160
rect 9864 22040 9916 22092
rect 11336 22040 11388 22092
rect 8944 21972 8996 22024
rect 11888 22015 11940 22024
rect 11888 21981 11894 22015
rect 11894 21981 11928 22015
rect 11928 21981 11940 22015
rect 11888 21972 11940 21981
rect 12808 21972 12860 22024
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 17592 22040 17644 22092
rect 19892 22083 19944 22092
rect 19892 22049 19901 22083
rect 19901 22049 19935 22083
rect 19935 22049 19944 22083
rect 19892 22040 19944 22049
rect 17960 21972 18012 22024
rect 19432 21972 19484 22024
rect 10784 21904 10836 21956
rect 12900 21947 12952 21956
rect 12900 21913 12909 21947
rect 12909 21913 12943 21947
rect 12943 21913 12952 21947
rect 12900 21904 12952 21913
rect 14464 21904 14516 21956
rect 19064 21904 19116 21956
rect 20076 21972 20128 22024
rect 21364 22108 21416 22160
rect 20628 21972 20680 22024
rect 21088 22040 21140 22092
rect 27988 22108 28040 22160
rect 43168 22108 43220 22160
rect 43904 22108 43956 22160
rect 20996 21972 21048 22024
rect 22100 21972 22152 22024
rect 25964 22040 26016 22092
rect 26700 22040 26752 22092
rect 27344 22040 27396 22092
rect 29644 22083 29696 22092
rect 29644 22049 29653 22083
rect 29653 22049 29687 22083
rect 29687 22049 29696 22083
rect 29644 22040 29696 22049
rect 30012 22040 30064 22092
rect 31576 22040 31628 22092
rect 20904 21904 20956 21956
rect 21180 21947 21232 21956
rect 21180 21913 21189 21947
rect 21189 21913 21223 21947
rect 21223 21913 21232 21947
rect 21180 21904 21232 21913
rect 23296 21904 23348 21956
rect 11612 21836 11664 21888
rect 11888 21879 11940 21888
rect 11888 21845 11897 21879
rect 11897 21845 11931 21879
rect 11931 21845 11940 21879
rect 11888 21836 11940 21845
rect 13912 21836 13964 21888
rect 16212 21879 16264 21888
rect 16212 21845 16221 21879
rect 16221 21845 16255 21879
rect 16255 21845 16264 21879
rect 16212 21836 16264 21845
rect 20536 21836 20588 21888
rect 20812 21836 20864 21888
rect 22560 21836 22612 21888
rect 23664 21879 23716 21888
rect 23664 21845 23673 21879
rect 23673 21845 23707 21879
rect 23707 21845 23716 21879
rect 23664 21836 23716 21845
rect 25504 21879 25556 21888
rect 25504 21845 25513 21879
rect 25513 21845 25547 21879
rect 25547 21845 25556 21879
rect 25504 21836 25556 21845
rect 28172 21972 28224 22024
rect 29184 21972 29236 22024
rect 29460 21972 29512 22024
rect 26332 21947 26384 21956
rect 26332 21913 26341 21947
rect 26341 21913 26375 21947
rect 26375 21913 26384 21947
rect 26332 21904 26384 21913
rect 27068 21904 27120 21956
rect 26700 21836 26752 21888
rect 27160 21836 27212 21888
rect 29000 21904 29052 21956
rect 28724 21836 28776 21888
rect 29092 21836 29144 21888
rect 32404 21947 32456 21956
rect 32404 21913 32413 21947
rect 32413 21913 32447 21947
rect 32447 21913 32456 21947
rect 32404 21904 32456 21913
rect 33968 21972 34020 22024
rect 40040 22015 40092 22024
rect 40040 21981 40049 22015
rect 40049 21981 40083 22015
rect 40083 21981 40092 22015
rect 40040 21972 40092 21981
rect 43168 22015 43220 22024
rect 34060 21904 34112 21956
rect 35808 21947 35860 21956
rect 35808 21913 35817 21947
rect 35817 21913 35851 21947
rect 35851 21913 35860 21947
rect 35808 21904 35860 21913
rect 43168 21981 43177 22015
rect 43177 21981 43211 22015
rect 43211 21981 43220 22015
rect 43168 21972 43220 21981
rect 43260 21972 43312 22024
rect 43904 21947 43956 21956
rect 43904 21913 43913 21947
rect 43913 21913 43947 21947
rect 43947 21913 43956 21947
rect 43904 21904 43956 21913
rect 43996 21904 44048 21956
rect 47400 22040 47452 22092
rect 47676 22040 47728 22092
rect 45192 22015 45244 22024
rect 45192 21981 45201 22015
rect 45201 21981 45235 22015
rect 45235 21981 45244 22015
rect 45192 21972 45244 21981
rect 45284 21972 45336 22024
rect 48044 21972 48096 22024
rect 45560 21904 45612 21956
rect 44272 21879 44324 21888
rect 44272 21845 44281 21879
rect 44281 21845 44315 21879
rect 44315 21845 44324 21879
rect 44272 21836 44324 21845
rect 45468 21836 45520 21888
rect 47124 21904 47176 21956
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 12164 21632 12216 21684
rect 12900 21632 12952 21684
rect 17040 21632 17092 21684
rect 19340 21632 19392 21684
rect 19984 21632 20036 21684
rect 21272 21632 21324 21684
rect 21732 21632 21784 21684
rect 11428 21564 11480 21616
rect 12440 21607 12492 21616
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 12440 21573 12449 21607
rect 12449 21573 12483 21607
rect 12483 21573 12492 21607
rect 12440 21564 12492 21573
rect 21180 21564 21232 21616
rect 22560 21607 22612 21616
rect 22560 21573 22569 21607
rect 22569 21573 22603 21607
rect 22603 21573 22612 21607
rect 22560 21564 22612 21573
rect 25504 21564 25556 21616
rect 11704 21496 11756 21505
rect 11888 21496 11940 21548
rect 12348 21496 12400 21548
rect 14924 21539 14976 21548
rect 9036 21428 9088 21480
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 16212 21496 16264 21548
rect 17316 21539 17368 21548
rect 17316 21505 17325 21539
rect 17325 21505 17359 21539
rect 17359 21505 17368 21539
rect 17316 21496 17368 21505
rect 17960 21496 18012 21548
rect 19432 21539 19484 21548
rect 19432 21505 19441 21539
rect 19441 21505 19475 21539
rect 19475 21505 19484 21539
rect 19432 21496 19484 21505
rect 20076 21539 20128 21548
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 7932 21360 7984 21412
rect 8944 21292 8996 21344
rect 18236 21428 18288 21480
rect 18604 21428 18656 21480
rect 20812 21496 20864 21548
rect 20536 21428 20588 21480
rect 20996 21428 21048 21480
rect 12808 21403 12860 21412
rect 12808 21369 12817 21403
rect 12817 21369 12851 21403
rect 12851 21369 12860 21403
rect 12808 21360 12860 21369
rect 14096 21360 14148 21412
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 12164 21292 12216 21344
rect 14280 21292 14332 21344
rect 14372 21292 14424 21344
rect 18236 21292 18288 21344
rect 20628 21360 20680 21412
rect 23664 21496 23716 21548
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 28172 21607 28224 21616
rect 28172 21573 28197 21607
rect 28197 21573 28224 21607
rect 28172 21564 28224 21573
rect 28724 21564 28776 21616
rect 28908 21496 28960 21548
rect 29184 21564 29236 21616
rect 30288 21564 30340 21616
rect 31576 21607 31628 21616
rect 29736 21539 29788 21548
rect 22284 21471 22336 21480
rect 22284 21437 22293 21471
rect 22293 21437 22327 21471
rect 22327 21437 22336 21471
rect 22284 21428 22336 21437
rect 23296 21428 23348 21480
rect 24124 21428 24176 21480
rect 25320 21428 25372 21480
rect 21456 21292 21508 21344
rect 26332 21360 26384 21412
rect 28356 21403 28408 21412
rect 28356 21369 28365 21403
rect 28365 21369 28399 21403
rect 28399 21369 28408 21403
rect 28356 21360 28408 21369
rect 29736 21505 29745 21539
rect 29745 21505 29779 21539
rect 29779 21505 29788 21539
rect 29736 21496 29788 21505
rect 31576 21573 31585 21607
rect 31585 21573 31619 21607
rect 31619 21573 31628 21607
rect 31576 21564 31628 21573
rect 32404 21632 32456 21684
rect 33968 21675 34020 21684
rect 33968 21641 33977 21675
rect 33977 21641 34011 21675
rect 34011 21641 34020 21675
rect 33968 21632 34020 21641
rect 42708 21632 42760 21684
rect 35072 21607 35124 21616
rect 35072 21573 35081 21607
rect 35081 21573 35115 21607
rect 35115 21573 35124 21607
rect 35072 21564 35124 21573
rect 36360 21564 36412 21616
rect 38384 21564 38436 21616
rect 46112 21632 46164 21684
rect 47768 21632 47820 21684
rect 45100 21564 45152 21616
rect 45192 21564 45244 21616
rect 47676 21564 47728 21616
rect 34796 21496 34848 21548
rect 39948 21539 40000 21548
rect 39948 21505 39957 21539
rect 39957 21505 39991 21539
rect 39991 21505 40000 21539
rect 39948 21496 40000 21505
rect 40132 21539 40184 21548
rect 40132 21505 40141 21539
rect 40141 21505 40175 21539
rect 40175 21505 40184 21539
rect 40132 21496 40184 21505
rect 42892 21496 42944 21548
rect 43260 21496 43312 21548
rect 43536 21496 43588 21548
rect 44180 21496 44232 21548
rect 44548 21496 44600 21548
rect 46204 21539 46256 21548
rect 46204 21505 46213 21539
rect 46213 21505 46247 21539
rect 46247 21505 46256 21539
rect 46204 21496 46256 21505
rect 22008 21292 22060 21344
rect 26240 21335 26292 21344
rect 26240 21301 26249 21335
rect 26249 21301 26283 21335
rect 26283 21301 26292 21335
rect 26240 21292 26292 21301
rect 28724 21292 28776 21344
rect 29000 21292 29052 21344
rect 32404 21335 32456 21344
rect 32404 21301 32413 21335
rect 32413 21301 32447 21335
rect 32447 21301 32456 21335
rect 32404 21292 32456 21301
rect 35808 21471 35860 21480
rect 33600 21335 33652 21344
rect 33600 21301 33609 21335
rect 33609 21301 33643 21335
rect 33643 21301 33652 21335
rect 33600 21292 33652 21301
rect 35808 21437 35817 21471
rect 35817 21437 35851 21471
rect 35851 21437 35860 21471
rect 35808 21428 35860 21437
rect 43904 21428 43956 21480
rect 44456 21428 44508 21480
rect 47032 21496 47084 21548
rect 47584 21539 47636 21548
rect 47584 21505 47593 21539
rect 47593 21505 47627 21539
rect 47627 21505 47636 21539
rect 47584 21496 47636 21505
rect 46480 21471 46532 21480
rect 46480 21437 46489 21471
rect 46489 21437 46523 21471
rect 46523 21437 46532 21471
rect 46480 21428 46532 21437
rect 47860 21471 47912 21480
rect 47860 21437 47869 21471
rect 47869 21437 47903 21471
rect 47903 21437 47912 21471
rect 47860 21428 47912 21437
rect 37004 21360 37056 21412
rect 46020 21360 46072 21412
rect 38384 21292 38436 21344
rect 40132 21292 40184 21344
rect 43628 21292 43680 21344
rect 45468 21292 45520 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 9036 21131 9088 21140
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 2872 21020 2924 21072
rect 11520 21063 11572 21072
rect 11520 21029 11529 21063
rect 11529 21029 11563 21063
rect 11563 21029 11572 21063
rect 11520 21020 11572 21029
rect 19340 21088 19392 21140
rect 20628 21088 20680 21140
rect 20996 21131 21048 21140
rect 20996 21097 21005 21131
rect 21005 21097 21039 21131
rect 21039 21097 21048 21131
rect 20996 21088 21048 21097
rect 22284 21088 22336 21140
rect 25320 21131 25372 21140
rect 25320 21097 25329 21131
rect 25329 21097 25363 21131
rect 25363 21097 25372 21131
rect 25320 21088 25372 21097
rect 31116 21088 31168 21140
rect 46480 21088 46532 21140
rect 47216 21088 47268 21140
rect 47860 21088 47912 21140
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 14280 20995 14332 21004
rect 14280 20961 14289 20995
rect 14289 20961 14323 20995
rect 14323 20961 14332 20995
rect 14280 20952 14332 20961
rect 33600 21020 33652 21072
rect 43720 21020 43772 21072
rect 17316 20952 17368 21004
rect 17960 20995 18012 21004
rect 14096 20927 14148 20936
rect 20 20816 72 20868
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 21456 20995 21508 21004
rect 21456 20961 21465 20995
rect 21465 20961 21499 20995
rect 21499 20961 21508 20995
rect 21456 20952 21508 20961
rect 22100 20952 22152 21004
rect 28172 20952 28224 21004
rect 28540 20952 28592 21004
rect 19340 20884 19392 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 21364 20884 21416 20936
rect 12808 20816 12860 20868
rect 16580 20859 16632 20868
rect 16580 20825 16589 20859
rect 16589 20825 16623 20859
rect 16623 20825 16632 20859
rect 16580 20816 16632 20825
rect 19248 20816 19300 20868
rect 11796 20748 11848 20800
rect 19432 20748 19484 20800
rect 20720 20816 20772 20868
rect 20996 20816 21048 20868
rect 23204 20884 23256 20936
rect 26240 20884 26292 20936
rect 28264 20927 28316 20936
rect 28264 20893 28273 20927
rect 28273 20893 28307 20927
rect 28307 20893 28316 20927
rect 28264 20884 28316 20893
rect 29460 20884 29512 20936
rect 30380 20884 30432 20936
rect 34060 20952 34112 21004
rect 33140 20927 33192 20936
rect 33140 20893 33149 20927
rect 33149 20893 33183 20927
rect 33183 20893 33192 20927
rect 33140 20884 33192 20893
rect 43260 20952 43312 21004
rect 43352 20995 43404 21004
rect 43352 20961 43361 20995
rect 43361 20961 43395 20995
rect 43395 20961 43404 20995
rect 43628 20995 43680 21004
rect 43352 20952 43404 20961
rect 43628 20961 43637 20995
rect 43637 20961 43671 20995
rect 43671 20961 43680 20995
rect 43628 20952 43680 20961
rect 43444 20927 43496 20936
rect 28448 20859 28500 20868
rect 28448 20825 28457 20859
rect 28457 20825 28491 20859
rect 28491 20825 28500 20859
rect 28448 20816 28500 20825
rect 31024 20859 31076 20868
rect 31024 20825 31033 20859
rect 31033 20825 31067 20859
rect 31067 20825 31076 20859
rect 31024 20816 31076 20825
rect 37004 20816 37056 20868
rect 43444 20893 43453 20927
rect 43453 20893 43487 20927
rect 43487 20893 43496 20927
rect 43444 20884 43496 20893
rect 42984 20816 43036 20868
rect 43904 20884 43956 20936
rect 45468 20927 45520 20936
rect 43996 20816 44048 20868
rect 45468 20893 45477 20927
rect 45477 20893 45511 20927
rect 45511 20893 45520 20927
rect 45468 20884 45520 20893
rect 46940 21020 46992 21072
rect 47584 21020 47636 21072
rect 47860 20952 47912 21004
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 46480 20859 46532 20868
rect 46480 20825 46489 20859
rect 46489 20825 46523 20859
rect 46523 20825 46532 20859
rect 46480 20816 46532 20825
rect 23296 20791 23348 20800
rect 23296 20757 23305 20791
rect 23305 20757 23339 20791
rect 23339 20757 23348 20791
rect 23296 20748 23348 20757
rect 29736 20748 29788 20800
rect 33232 20791 33284 20800
rect 33232 20757 33241 20791
rect 33241 20757 33275 20791
rect 33275 20757 33284 20791
rect 33232 20748 33284 20757
rect 43076 20748 43128 20800
rect 43444 20748 43496 20800
rect 44088 20748 44140 20800
rect 45836 20791 45888 20800
rect 45836 20757 45845 20791
rect 45845 20757 45879 20791
rect 45879 20757 45888 20791
rect 45836 20748 45888 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2964 20544 3016 20596
rect 11796 20519 11848 20528
rect 11796 20485 11805 20519
rect 11805 20485 11839 20519
rect 11839 20485 11848 20519
rect 11796 20476 11848 20485
rect 12072 20476 12124 20528
rect 16580 20544 16632 20596
rect 19156 20544 19208 20596
rect 21824 20544 21876 20596
rect 23112 20544 23164 20596
rect 17960 20476 18012 20528
rect 18236 20519 18288 20528
rect 18236 20485 18245 20519
rect 18245 20485 18279 20519
rect 18279 20485 18288 20519
rect 18236 20476 18288 20485
rect 18972 20476 19024 20528
rect 16212 20408 16264 20460
rect 16764 20408 16816 20460
rect 17868 20408 17920 20460
rect 20812 20408 20864 20460
rect 22008 20476 22060 20528
rect 24124 20519 24176 20528
rect 24124 20485 24133 20519
rect 24133 20485 24167 20519
rect 24167 20485 24176 20519
rect 24124 20476 24176 20485
rect 23204 20408 23256 20460
rect 23296 20408 23348 20460
rect 10692 20340 10744 20392
rect 12440 20340 12492 20392
rect 15476 20340 15528 20392
rect 16120 20383 16172 20392
rect 16120 20349 16129 20383
rect 16129 20349 16163 20383
rect 16163 20349 16172 20383
rect 16120 20340 16172 20349
rect 17960 20383 18012 20392
rect 17960 20349 17969 20383
rect 17969 20349 18003 20383
rect 18003 20349 18012 20383
rect 17960 20340 18012 20349
rect 18604 20340 18656 20392
rect 20536 20383 20588 20392
rect 19340 20272 19392 20324
rect 20536 20349 20545 20383
rect 20545 20349 20579 20383
rect 20579 20349 20588 20383
rect 20536 20340 20588 20349
rect 29000 20476 29052 20528
rect 29736 20476 29788 20528
rect 33232 20476 33284 20528
rect 43260 20476 43312 20528
rect 28448 20451 28500 20460
rect 28448 20417 28457 20451
rect 28457 20417 28491 20451
rect 28491 20417 28500 20451
rect 28448 20408 28500 20417
rect 32128 20451 32180 20460
rect 32128 20417 32137 20451
rect 32137 20417 32171 20451
rect 32171 20417 32180 20451
rect 32128 20408 32180 20417
rect 43076 20451 43128 20460
rect 43076 20417 43085 20451
rect 43085 20417 43119 20451
rect 43119 20417 43128 20451
rect 43076 20408 43128 20417
rect 43444 20451 43496 20460
rect 43444 20417 43453 20451
rect 43453 20417 43487 20451
rect 43487 20417 43496 20451
rect 43444 20408 43496 20417
rect 44364 20408 44416 20460
rect 44732 20451 44784 20460
rect 44732 20417 44741 20451
rect 44741 20417 44775 20451
rect 44775 20417 44784 20451
rect 44732 20408 44784 20417
rect 46480 20544 46532 20596
rect 48044 20587 48096 20596
rect 48044 20553 48053 20587
rect 48053 20553 48087 20587
rect 48087 20553 48096 20587
rect 48044 20544 48096 20553
rect 45836 20408 45888 20460
rect 47400 20408 47452 20460
rect 29092 20340 29144 20392
rect 34428 20383 34480 20392
rect 34428 20349 34437 20383
rect 34437 20349 34471 20383
rect 34471 20349 34480 20383
rect 34428 20340 34480 20349
rect 43904 20340 43956 20392
rect 45744 20340 45796 20392
rect 17040 20204 17092 20256
rect 19892 20204 19944 20256
rect 21916 20247 21968 20256
rect 21916 20213 21925 20247
rect 21925 20213 21959 20247
rect 21959 20213 21968 20247
rect 21916 20204 21968 20213
rect 32220 20247 32272 20256
rect 32220 20213 32229 20247
rect 32229 20213 32263 20247
rect 32263 20213 32272 20247
rect 32220 20204 32272 20213
rect 47676 20247 47728 20256
rect 47676 20213 47685 20247
rect 47685 20213 47719 20247
rect 47719 20213 47728 20247
rect 47676 20204 47728 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3424 20000 3476 20052
rect 27252 20000 27304 20052
rect 28632 20000 28684 20052
rect 31024 20000 31076 20052
rect 42984 20043 43036 20052
rect 42984 20009 42993 20043
rect 42993 20009 43027 20043
rect 43027 20009 43036 20043
rect 42984 20000 43036 20009
rect 43352 20000 43404 20052
rect 47860 20000 47912 20052
rect 10692 19975 10744 19984
rect 10692 19941 10701 19975
rect 10701 19941 10735 19975
rect 10735 19941 10744 19975
rect 10692 19932 10744 19941
rect 12072 19975 12124 19984
rect 12072 19941 12081 19975
rect 12081 19941 12115 19975
rect 12115 19941 12124 19975
rect 12072 19932 12124 19941
rect 15476 19975 15528 19984
rect 15476 19941 15485 19975
rect 15485 19941 15519 19975
rect 15519 19941 15528 19975
rect 15476 19932 15528 19941
rect 23296 19932 23348 19984
rect 27344 19932 27396 19984
rect 16856 19907 16908 19916
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 17040 19907 17092 19916
rect 17040 19873 17049 19907
rect 17049 19873 17083 19907
rect 17083 19873 17092 19907
rect 17040 19864 17092 19873
rect 19432 19864 19484 19916
rect 19892 19907 19944 19916
rect 19892 19873 19901 19907
rect 19901 19873 19935 19907
rect 19935 19873 19944 19907
rect 19892 19864 19944 19873
rect 19984 19864 20036 19916
rect 1768 19796 1820 19848
rect 11336 19796 11388 19848
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 14372 19839 14424 19848
rect 10876 19728 10928 19780
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 15108 19796 15160 19848
rect 16764 19796 16816 19848
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 23388 19796 23440 19848
rect 26332 19796 26384 19848
rect 27252 19864 27304 19916
rect 27344 19796 27396 19848
rect 13268 19728 13320 19780
rect 19984 19728 20036 19780
rect 21916 19728 21968 19780
rect 22284 19771 22336 19780
rect 22284 19737 22293 19771
rect 22293 19737 22327 19771
rect 22327 19737 22336 19771
rect 22284 19728 22336 19737
rect 24584 19728 24636 19780
rect 30472 19796 30524 19848
rect 31300 19839 31352 19848
rect 31300 19805 31309 19839
rect 31309 19805 31343 19839
rect 31343 19805 31352 19839
rect 31300 19796 31352 19805
rect 44180 19932 44232 19984
rect 43904 19864 43956 19916
rect 45744 19907 45796 19916
rect 45744 19873 45753 19907
rect 45753 19873 45787 19907
rect 45787 19873 45796 19907
rect 45744 19864 45796 19873
rect 46940 19907 46992 19916
rect 46940 19873 46949 19907
rect 46949 19873 46983 19907
rect 46983 19873 46992 19907
rect 46940 19864 46992 19873
rect 47124 19864 47176 19916
rect 42892 19839 42944 19848
rect 42892 19805 42901 19839
rect 42901 19805 42935 19839
rect 42935 19805 42944 19839
rect 42892 19796 42944 19805
rect 43076 19839 43128 19848
rect 43076 19805 43085 19839
rect 43085 19805 43119 19839
rect 43119 19805 43128 19839
rect 43076 19796 43128 19805
rect 43536 19796 43588 19848
rect 43812 19839 43864 19848
rect 43812 19805 43821 19839
rect 43821 19805 43855 19839
rect 43855 19805 43864 19839
rect 43812 19796 43864 19805
rect 43996 19839 44048 19848
rect 43996 19805 44005 19839
rect 44005 19805 44039 19839
rect 44039 19805 44048 19839
rect 43996 19796 44048 19805
rect 12900 19660 12952 19712
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 20628 19660 20680 19712
rect 27068 19660 27120 19712
rect 46572 19728 46624 19780
rect 32220 19660 32272 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 14096 19456 14148 19508
rect 14464 19388 14516 19440
rect 17960 19456 18012 19508
rect 18972 19456 19024 19508
rect 22284 19456 22336 19508
rect 26332 19499 26384 19508
rect 26332 19465 26341 19499
rect 26341 19465 26375 19499
rect 26375 19465 26384 19499
rect 26332 19456 26384 19465
rect 31300 19456 31352 19508
rect 31944 19456 31996 19508
rect 43444 19499 43496 19508
rect 43444 19465 43453 19499
rect 43453 19465 43487 19499
rect 43487 19465 43496 19499
rect 43444 19456 43496 19465
rect 44548 19456 44600 19508
rect 46020 19456 46072 19508
rect 47308 19456 47360 19508
rect 16856 19388 16908 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 11980 19320 12032 19372
rect 12900 19363 12952 19372
rect 12900 19329 12909 19363
rect 12909 19329 12943 19363
rect 12943 19329 12952 19363
rect 12900 19320 12952 19329
rect 14740 19320 14792 19372
rect 19340 19388 19392 19440
rect 22008 19388 22060 19440
rect 34060 19388 34112 19440
rect 46388 19388 46440 19440
rect 47400 19388 47452 19440
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 13176 19295 13228 19304
rect 13176 19261 13185 19295
rect 13185 19261 13219 19295
rect 13219 19261 13228 19295
rect 13176 19252 13228 19261
rect 14372 19252 14424 19304
rect 19156 19320 19208 19372
rect 23296 19320 23348 19372
rect 26148 19363 26200 19372
rect 26148 19329 26157 19363
rect 26157 19329 26191 19363
rect 26191 19329 26200 19363
rect 26148 19320 26200 19329
rect 26516 19320 26568 19372
rect 15660 19295 15712 19304
rect 15660 19261 15669 19295
rect 15669 19261 15703 19295
rect 15703 19261 15712 19295
rect 15660 19252 15712 19261
rect 19064 19252 19116 19304
rect 19524 19252 19576 19304
rect 25596 19252 25648 19304
rect 28264 19363 28316 19372
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 28632 19320 28684 19372
rect 31208 19320 31260 19372
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 43352 19363 43404 19372
rect 43352 19329 43361 19363
rect 43361 19329 43395 19363
rect 43395 19329 43404 19363
rect 43352 19320 43404 19329
rect 44088 19363 44140 19372
rect 44088 19329 44097 19363
rect 44097 19329 44131 19363
rect 44131 19329 44140 19363
rect 44088 19320 44140 19329
rect 44272 19363 44324 19372
rect 44272 19329 44281 19363
rect 44281 19329 44315 19363
rect 44315 19329 44324 19363
rect 44272 19320 44324 19329
rect 46756 19320 46808 19372
rect 35348 19184 35400 19236
rect 47032 19184 47084 19236
rect 10416 19116 10468 19168
rect 11704 19116 11756 19168
rect 26792 19116 26844 19168
rect 28908 19159 28960 19168
rect 28908 19125 28917 19159
rect 28917 19125 28951 19159
rect 28951 19125 28960 19159
rect 28908 19116 28960 19125
rect 32220 19159 32272 19168
rect 32220 19125 32229 19159
rect 32229 19125 32263 19159
rect 32263 19125 32272 19159
rect 32220 19116 32272 19125
rect 47768 19159 47820 19168
rect 47768 19125 47777 19159
rect 47777 19125 47811 19159
rect 47811 19125 47820 19159
rect 47768 19116 47820 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 4988 18912 5040 18964
rect 29000 18912 29052 18964
rect 13176 18844 13228 18896
rect 13820 18844 13872 18896
rect 22376 18844 22428 18896
rect 10416 18819 10468 18828
rect 10416 18785 10425 18819
rect 10425 18785 10459 18819
rect 10459 18785 10468 18819
rect 10416 18776 10468 18785
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 12348 18708 12400 18760
rect 14096 18708 14148 18760
rect 14740 18708 14792 18760
rect 19524 18708 19576 18760
rect 20812 18708 20864 18760
rect 10968 18640 11020 18692
rect 11704 18640 11756 18692
rect 14464 18683 14516 18692
rect 12164 18615 12216 18624
rect 12164 18581 12173 18615
rect 12173 18581 12207 18615
rect 12207 18581 12216 18615
rect 12164 18572 12216 18581
rect 14464 18649 14473 18683
rect 14473 18649 14507 18683
rect 14507 18649 14516 18683
rect 14464 18640 14516 18649
rect 19340 18640 19392 18692
rect 23112 18776 23164 18828
rect 21824 18708 21876 18760
rect 23664 18776 23716 18828
rect 24492 18776 24544 18828
rect 13360 18572 13412 18624
rect 14372 18572 14424 18624
rect 14924 18572 14976 18624
rect 15016 18572 15068 18624
rect 16764 18572 16816 18624
rect 19432 18572 19484 18624
rect 24584 18708 24636 18760
rect 25596 18776 25648 18828
rect 26792 18819 26844 18828
rect 26792 18785 26801 18819
rect 26801 18785 26835 18819
rect 26835 18785 26844 18819
rect 26792 18776 26844 18785
rect 27068 18819 27120 18828
rect 27068 18785 27077 18819
rect 27077 18785 27111 18819
rect 27111 18785 27120 18819
rect 27068 18776 27120 18785
rect 35348 18912 35400 18964
rect 32220 18776 32272 18828
rect 32312 18819 32364 18828
rect 32312 18785 32321 18819
rect 32321 18785 32355 18819
rect 32355 18785 32364 18819
rect 32312 18776 32364 18785
rect 47768 18776 47820 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 25964 18751 26016 18760
rect 25964 18717 25973 18751
rect 25973 18717 26007 18751
rect 26007 18717 26016 18751
rect 25964 18708 26016 18717
rect 30012 18708 30064 18760
rect 30104 18751 30156 18760
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 31116 18708 31168 18760
rect 33508 18751 33560 18760
rect 33508 18717 33517 18751
rect 33517 18717 33551 18751
rect 33551 18717 33560 18751
rect 33508 18708 33560 18717
rect 35532 18708 35584 18760
rect 45836 18751 45888 18760
rect 45836 18717 45845 18751
rect 45845 18717 45879 18751
rect 45879 18717 45888 18751
rect 45836 18708 45888 18717
rect 19984 18572 20036 18624
rect 23296 18572 23348 18624
rect 24768 18572 24820 18624
rect 27252 18572 27304 18624
rect 28908 18640 28960 18692
rect 34612 18640 34664 18692
rect 47676 18640 47728 18692
rect 30196 18572 30248 18624
rect 34796 18572 34848 18624
rect 45652 18615 45704 18624
rect 45652 18581 45661 18615
rect 45661 18581 45695 18615
rect 45695 18581 45704 18615
rect 45652 18572 45704 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3424 18368 3476 18420
rect 47676 18411 47728 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 12348 18300 12400 18352
rect 14464 18300 14516 18352
rect 11520 18232 11572 18284
rect 12164 18232 12216 18284
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 16856 18300 16908 18352
rect 19432 18300 19484 18352
rect 23940 18300 23992 18352
rect 25504 18300 25556 18352
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 13820 18164 13872 18216
rect 15108 18232 15160 18284
rect 15660 18232 15712 18284
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 17040 18232 17092 18284
rect 19340 18232 19392 18284
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 23848 18232 23900 18284
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24768 18275 24820 18284
rect 24216 18232 24268 18241
rect 24768 18241 24777 18275
rect 24777 18241 24811 18275
rect 24811 18241 24820 18275
rect 24768 18232 24820 18241
rect 25688 18232 25740 18284
rect 26148 18300 26200 18352
rect 27252 18343 27304 18352
rect 27252 18309 27261 18343
rect 27261 18309 27295 18343
rect 27295 18309 27304 18343
rect 27252 18300 27304 18309
rect 28264 18300 28316 18352
rect 30012 18343 30064 18352
rect 30012 18309 30021 18343
rect 30021 18309 30055 18343
rect 30055 18309 30064 18343
rect 30012 18300 30064 18309
rect 30104 18300 30156 18352
rect 31208 18343 31260 18352
rect 31208 18309 31217 18343
rect 31217 18309 31251 18343
rect 31251 18309 31260 18343
rect 31208 18300 31260 18309
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 32312 18300 32364 18352
rect 33508 18300 33560 18352
rect 26424 18232 26476 18284
rect 34796 18275 34848 18284
rect 34796 18241 34805 18275
rect 34805 18241 34839 18275
rect 34839 18241 34848 18275
rect 34796 18232 34848 18241
rect 43904 18300 43956 18352
rect 46020 18275 46072 18284
rect 46020 18241 46029 18275
rect 46029 18241 46063 18275
rect 46063 18241 46072 18275
rect 46020 18232 46072 18241
rect 46388 18275 46440 18284
rect 46388 18241 46397 18275
rect 46397 18241 46431 18275
rect 46431 18241 46440 18275
rect 46388 18232 46440 18241
rect 46756 18275 46808 18284
rect 46756 18241 46765 18275
rect 46765 18241 46799 18275
rect 46799 18241 46808 18275
rect 46756 18232 46808 18241
rect 47032 18275 47084 18284
rect 47032 18241 47041 18275
rect 47041 18241 47075 18275
rect 47075 18241 47084 18275
rect 47032 18232 47084 18241
rect 47584 18275 47636 18284
rect 47584 18241 47593 18275
rect 47593 18241 47627 18275
rect 47627 18241 47636 18275
rect 47584 18232 47636 18241
rect 14556 18164 14608 18216
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 14924 18164 14976 18216
rect 15016 18096 15068 18148
rect 13820 18028 13872 18080
rect 15476 18028 15528 18080
rect 16580 18028 16632 18080
rect 19248 18028 19300 18080
rect 20628 18164 20680 18216
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 22100 18164 22152 18173
rect 23388 18164 23440 18216
rect 23940 18207 23992 18216
rect 23940 18173 23949 18207
rect 23949 18173 23983 18207
rect 23983 18173 23992 18207
rect 23940 18164 23992 18173
rect 24492 18164 24544 18216
rect 26976 18207 27028 18216
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 30288 18164 30340 18216
rect 31944 18164 31996 18216
rect 34060 18207 34112 18216
rect 34060 18173 34069 18207
rect 34069 18173 34103 18207
rect 34103 18173 34112 18207
rect 34060 18164 34112 18173
rect 43536 18207 43588 18216
rect 43536 18173 43545 18207
rect 43545 18173 43579 18207
rect 43579 18173 43588 18207
rect 43536 18164 43588 18173
rect 45192 18207 45244 18216
rect 45192 18173 45201 18207
rect 45201 18173 45235 18207
rect 45235 18173 45244 18207
rect 45192 18164 45244 18173
rect 47860 18164 47912 18216
rect 25688 18096 25740 18148
rect 22652 18028 22704 18080
rect 23480 18028 23532 18080
rect 24676 18028 24728 18080
rect 24860 18071 24912 18080
rect 24860 18037 24869 18071
rect 24869 18037 24903 18071
rect 24903 18037 24912 18071
rect 24860 18028 24912 18037
rect 25964 18028 26016 18080
rect 30380 18096 30432 18148
rect 35532 18096 35584 18148
rect 46756 18096 46808 18148
rect 33140 18028 33192 18080
rect 46296 18071 46348 18080
rect 46296 18037 46305 18071
rect 46305 18037 46339 18071
rect 46339 18037 46348 18071
rect 46296 18028 46348 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 14372 17824 14424 17876
rect 14648 17824 14700 17876
rect 16856 17824 16908 17876
rect 17040 17824 17092 17876
rect 23296 17824 23348 17876
rect 25596 17867 25648 17876
rect 14648 17688 14700 17740
rect 15016 17688 15068 17740
rect 15476 17731 15528 17740
rect 15476 17697 15485 17731
rect 15485 17697 15519 17731
rect 15519 17697 15528 17731
rect 15476 17688 15528 17697
rect 18420 17731 18472 17740
rect 18420 17697 18429 17731
rect 18429 17697 18463 17731
rect 18463 17697 18472 17731
rect 18420 17688 18472 17697
rect 13268 17620 13320 17672
rect 16580 17620 16632 17672
rect 19248 17663 19300 17672
rect 14740 17552 14792 17604
rect 15016 17552 15068 17604
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 21824 17620 21876 17672
rect 23204 17620 23256 17672
rect 24032 17756 24084 17808
rect 23848 17688 23900 17740
rect 25596 17833 25605 17867
rect 25605 17833 25639 17867
rect 25639 17833 25648 17867
rect 25596 17824 25648 17833
rect 26976 17824 27028 17876
rect 43536 17824 43588 17876
rect 44180 17824 44232 17876
rect 24676 17799 24728 17808
rect 24676 17765 24685 17799
rect 24685 17765 24719 17799
rect 24719 17765 24728 17799
rect 24676 17756 24728 17765
rect 30288 17731 30340 17740
rect 23664 17620 23716 17672
rect 30288 17697 30297 17731
rect 30297 17697 30331 17731
rect 30331 17697 30340 17731
rect 30288 17688 30340 17697
rect 31116 17688 31168 17740
rect 33140 17688 33192 17740
rect 25504 17663 25556 17672
rect 20536 17552 20588 17604
rect 21548 17595 21600 17604
rect 21548 17561 21557 17595
rect 21557 17561 21591 17595
rect 21591 17561 21600 17595
rect 21548 17552 21600 17561
rect 21916 17595 21968 17604
rect 21916 17561 21925 17595
rect 21925 17561 21959 17595
rect 21959 17561 21968 17595
rect 21916 17552 21968 17561
rect 13452 17484 13504 17536
rect 14924 17484 14976 17536
rect 19064 17484 19116 17536
rect 21824 17527 21876 17536
rect 21824 17493 21833 17527
rect 21833 17493 21867 17527
rect 21867 17493 21876 17527
rect 21824 17484 21876 17493
rect 23204 17484 23256 17536
rect 23388 17484 23440 17536
rect 23756 17552 23808 17604
rect 23940 17484 23992 17536
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 25688 17663 25740 17672
rect 25688 17629 25697 17663
rect 25697 17629 25731 17663
rect 25731 17629 25740 17663
rect 25688 17620 25740 17629
rect 26516 17663 26568 17672
rect 26516 17629 26525 17663
rect 26525 17629 26559 17663
rect 26559 17629 26568 17663
rect 26516 17620 26568 17629
rect 30196 17663 30248 17672
rect 30196 17629 30205 17663
rect 30205 17629 30239 17663
rect 30239 17629 30248 17663
rect 30196 17620 30248 17629
rect 35532 17688 35584 17740
rect 35348 17663 35400 17672
rect 35348 17629 35357 17663
rect 35357 17629 35391 17663
rect 35391 17629 35400 17663
rect 35348 17620 35400 17629
rect 46388 17756 46440 17808
rect 34060 17595 34112 17604
rect 34060 17561 34069 17595
rect 34069 17561 34103 17595
rect 34103 17561 34112 17595
rect 34060 17552 34112 17561
rect 35072 17552 35124 17604
rect 26884 17484 26936 17536
rect 42800 17620 42852 17672
rect 43536 17620 43588 17672
rect 45744 17688 45796 17740
rect 46848 17688 46900 17740
rect 44916 17620 44968 17672
rect 46940 17552 46992 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 44364 17527 44416 17536
rect 44364 17493 44373 17527
rect 44373 17493 44407 17527
rect 44407 17493 44416 17527
rect 44364 17484 44416 17493
rect 45008 17527 45060 17536
rect 45008 17493 45017 17527
rect 45017 17493 45051 17527
rect 45051 17493 45060 17527
rect 45008 17484 45060 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1584 17280 1636 17332
rect 26884 17280 26936 17332
rect 30288 17280 30340 17332
rect 34060 17280 34112 17332
rect 13820 17212 13872 17264
rect 20536 17212 20588 17264
rect 21824 17212 21876 17264
rect 23480 17255 23532 17264
rect 23480 17221 23489 17255
rect 23489 17221 23523 17255
rect 23523 17221 23532 17255
rect 23480 17212 23532 17221
rect 24860 17212 24912 17264
rect 3424 17144 3476 17196
rect 7932 17144 7984 17196
rect 13452 17187 13504 17196
rect 11060 17076 11112 17128
rect 13452 17153 13461 17187
rect 13461 17153 13495 17187
rect 13495 17153 13504 17187
rect 13452 17144 13504 17153
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 20628 17144 20680 17196
rect 15016 17076 15068 17128
rect 16948 17119 17000 17128
rect 16948 17085 16957 17119
rect 16957 17085 16991 17119
rect 16991 17085 17000 17119
rect 16948 17076 17000 17085
rect 19156 17076 19208 17128
rect 16672 17008 16724 17060
rect 22652 17144 22704 17196
rect 23204 17187 23256 17196
rect 23204 17153 23213 17187
rect 23213 17153 23247 17187
rect 23247 17153 23256 17187
rect 23204 17144 23256 17153
rect 27988 17144 28040 17196
rect 28264 17187 28316 17196
rect 28264 17153 28273 17187
rect 28273 17153 28307 17187
rect 28307 17153 28316 17187
rect 28264 17144 28316 17153
rect 28540 17144 28592 17196
rect 35072 17255 35124 17264
rect 35072 17221 35081 17255
rect 35081 17221 35115 17255
rect 35115 17221 35124 17255
rect 35072 17212 35124 17221
rect 24032 17076 24084 17128
rect 1400 16940 1452 16992
rect 11888 16940 11940 16992
rect 14372 16940 14424 16992
rect 21548 16940 21600 16992
rect 22100 17008 22152 17060
rect 27712 17008 27764 17060
rect 29000 17119 29052 17128
rect 29000 17085 29009 17119
rect 29009 17085 29043 17119
rect 29043 17085 29052 17119
rect 29000 17076 29052 17085
rect 29460 17076 29512 17128
rect 44916 17280 44968 17332
rect 45008 17280 45060 17332
rect 44456 17255 44508 17264
rect 44456 17221 44465 17255
rect 44465 17221 44499 17255
rect 44499 17221 44508 17255
rect 44456 17212 44508 17221
rect 43720 17187 43772 17196
rect 43720 17153 43729 17187
rect 43729 17153 43763 17187
rect 43763 17153 43772 17187
rect 43720 17144 43772 17153
rect 44364 17144 44416 17196
rect 46296 17212 46348 17264
rect 30012 17008 30064 17060
rect 30656 17008 30708 17060
rect 41420 17076 41472 17128
rect 42800 17008 42852 17060
rect 45652 17076 45704 17128
rect 46664 17144 46716 17196
rect 47032 17076 47084 17128
rect 22008 16940 22060 16992
rect 28080 16983 28132 16992
rect 28080 16949 28089 16983
rect 28089 16949 28123 16983
rect 28123 16949 28132 16983
rect 28080 16940 28132 16949
rect 29184 16983 29236 16992
rect 29184 16949 29193 16983
rect 29193 16949 29227 16983
rect 29227 16949 29236 16983
rect 29184 16940 29236 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 14372 16736 14424 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 16948 16736 17000 16788
rect 22284 16736 22336 16788
rect 11888 16643 11940 16652
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 11060 16585 11112 16594
rect 11060 16551 11069 16585
rect 11069 16551 11103 16585
rect 11103 16551 11112 16585
rect 11060 16542 11112 16551
rect 15016 16600 15068 16652
rect 17224 16668 17276 16720
rect 18604 16668 18656 16720
rect 21824 16668 21876 16720
rect 28540 16736 28592 16788
rect 45744 16779 45796 16788
rect 45744 16745 45753 16779
rect 45753 16745 45787 16779
rect 45787 16745 45796 16779
rect 45744 16736 45796 16745
rect 14924 16532 14976 16584
rect 18420 16600 18472 16652
rect 2136 16464 2188 16516
rect 3516 16464 3568 16516
rect 22100 16600 22152 16652
rect 23296 16600 23348 16652
rect 22008 16532 22060 16584
rect 27160 16575 27212 16584
rect 27160 16541 27169 16575
rect 27169 16541 27203 16575
rect 27203 16541 27212 16575
rect 27160 16532 27212 16541
rect 27252 16532 27304 16584
rect 27712 16532 27764 16584
rect 28080 16600 28132 16652
rect 30656 16643 30708 16652
rect 30656 16609 30665 16643
rect 30665 16609 30699 16643
rect 30699 16609 30708 16643
rect 30656 16600 30708 16609
rect 45652 16668 45704 16720
rect 43720 16600 43772 16652
rect 29828 16575 29880 16584
rect 22376 16464 22428 16516
rect 23664 16464 23716 16516
rect 28632 16507 28684 16516
rect 28632 16473 28641 16507
rect 28641 16473 28675 16507
rect 28675 16473 28684 16507
rect 28632 16464 28684 16473
rect 29828 16541 29837 16575
rect 29837 16541 29871 16575
rect 29871 16541 29880 16575
rect 29828 16532 29880 16541
rect 35992 16532 36044 16584
rect 36544 16532 36596 16584
rect 47492 16600 47544 16652
rect 11704 16396 11756 16448
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 21548 16396 21600 16448
rect 23848 16396 23900 16448
rect 27804 16396 27856 16448
rect 28724 16439 28776 16448
rect 28724 16405 28733 16439
rect 28733 16405 28767 16439
rect 28767 16405 28776 16439
rect 28724 16396 28776 16405
rect 28908 16396 28960 16448
rect 47676 16464 47728 16516
rect 48136 16507 48188 16516
rect 48136 16473 48145 16507
rect 48145 16473 48179 16507
rect 48179 16473 48188 16507
rect 48136 16464 48188 16473
rect 46572 16396 46624 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 1952 16056 2004 16108
rect 11704 16167 11756 16176
rect 11704 16133 11713 16167
rect 11713 16133 11747 16167
rect 11747 16133 11756 16167
rect 11704 16124 11756 16133
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 11520 16056 11572 16065
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 15660 15988 15712 16040
rect 18604 16124 18656 16176
rect 19248 16124 19300 16176
rect 18420 16056 18472 16108
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 21916 16192 21968 16244
rect 22376 16192 22428 16244
rect 20720 16124 20772 16176
rect 22468 16124 22520 16176
rect 19064 16056 19116 16065
rect 20628 16056 20680 16108
rect 22008 16056 22060 16108
rect 27988 16192 28040 16244
rect 28264 16192 28316 16244
rect 29828 16192 29880 16244
rect 36544 16192 36596 16244
rect 46940 16235 46992 16244
rect 24768 16124 24820 16176
rect 28908 16124 28960 16176
rect 46940 16201 46949 16235
rect 46949 16201 46983 16235
rect 46983 16201 46992 16235
rect 46940 16192 46992 16201
rect 47676 16235 47728 16244
rect 47676 16201 47685 16235
rect 47685 16201 47719 16235
rect 47719 16201 47728 16235
rect 47676 16192 47728 16201
rect 23848 16099 23900 16108
rect 19984 15988 20036 16040
rect 23848 16065 23857 16099
rect 23857 16065 23891 16099
rect 23891 16065 23900 16099
rect 23848 16056 23900 16065
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27252 16056 27304 16108
rect 27804 16056 27856 16108
rect 28632 16056 28684 16108
rect 29184 16056 29236 16108
rect 44456 16099 44508 16108
rect 23756 15988 23808 16040
rect 19156 15920 19208 15972
rect 14556 15852 14608 15904
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 17592 15852 17644 15904
rect 19340 15852 19392 15904
rect 19432 15852 19484 15904
rect 20628 15895 20680 15904
rect 20628 15861 20637 15895
rect 20637 15861 20671 15895
rect 20671 15861 20680 15895
rect 20628 15852 20680 15861
rect 22100 15963 22152 15972
rect 22100 15929 22109 15963
rect 22109 15929 22143 15963
rect 22143 15929 22152 15963
rect 22100 15920 22152 15929
rect 24584 15988 24636 16040
rect 28724 15988 28776 16040
rect 29460 15988 29512 16040
rect 44456 16065 44465 16099
rect 44465 16065 44499 16099
rect 44499 16065 44508 16099
rect 44456 16056 44508 16065
rect 47124 16056 47176 16108
rect 47400 16056 47452 16108
rect 45560 15988 45612 16040
rect 46112 16031 46164 16040
rect 46112 15997 46121 16031
rect 46121 15997 46155 16031
rect 46155 15997 46164 16031
rect 46112 15988 46164 15997
rect 47124 15920 47176 15972
rect 25504 15852 25556 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 5448 15512 5500 15564
rect 24584 15648 24636 15700
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 25504 15648 25556 15700
rect 45560 15648 45612 15700
rect 47492 15648 47544 15700
rect 18604 15623 18656 15632
rect 18604 15589 18613 15623
rect 18613 15589 18647 15623
rect 18647 15589 18656 15623
rect 18604 15580 18656 15589
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 16856 15555 16908 15564
rect 16856 15521 16865 15555
rect 16865 15521 16899 15555
rect 16899 15521 16908 15555
rect 16856 15512 16908 15521
rect 19340 15555 19392 15564
rect 19340 15521 19349 15555
rect 19349 15521 19383 15555
rect 19383 15521 19392 15555
rect 19340 15512 19392 15521
rect 21548 15555 21600 15564
rect 21548 15521 21557 15555
rect 21557 15521 21591 15555
rect 21591 15521 21600 15555
rect 21548 15512 21600 15521
rect 1768 15444 1820 15496
rect 19984 15444 20036 15496
rect 24676 15487 24728 15496
rect 24676 15453 24685 15487
rect 24685 15453 24719 15487
rect 24719 15453 24728 15487
rect 24676 15444 24728 15453
rect 43536 15487 43588 15496
rect 43536 15453 43545 15487
rect 43545 15453 43579 15487
rect 43579 15453 43588 15487
rect 43536 15444 43588 15453
rect 14832 15419 14884 15428
rect 14832 15385 14841 15419
rect 14841 15385 14875 15419
rect 14875 15385 14884 15419
rect 14832 15376 14884 15385
rect 15568 15376 15620 15428
rect 17132 15419 17184 15428
rect 17132 15385 17141 15419
rect 17141 15385 17175 15419
rect 17175 15385 17184 15419
rect 17132 15376 17184 15385
rect 17592 15376 17644 15428
rect 19340 15376 19392 15428
rect 22284 15376 22336 15428
rect 16304 15351 16356 15360
rect 16304 15317 16313 15351
rect 16313 15317 16347 15351
rect 16347 15317 16356 15351
rect 16304 15308 16356 15317
rect 19432 15308 19484 15360
rect 22468 15308 22520 15360
rect 43812 15308 43864 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 15568 15147 15620 15156
rect 15568 15113 15577 15147
rect 15577 15113 15611 15147
rect 15611 15113 15620 15147
rect 15568 15104 15620 15113
rect 17132 15104 17184 15156
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 14740 15036 14792 15088
rect 16304 15036 16356 15088
rect 15660 14968 15712 15020
rect 22284 15104 22336 15156
rect 18420 15079 18472 15088
rect 18420 15045 18429 15079
rect 18429 15045 18463 15079
rect 18463 15045 18472 15079
rect 18420 15036 18472 15045
rect 18880 15036 18932 15088
rect 19432 15036 19484 15088
rect 43812 15079 43864 15088
rect 43812 15045 43821 15079
rect 43821 15045 43855 15079
rect 43855 15045 43864 15079
rect 43812 15036 43864 15045
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 14832 14900 14884 14952
rect 14924 14832 14976 14884
rect 18512 14968 18564 15020
rect 20628 14968 20680 15020
rect 22008 14968 22060 15020
rect 24676 14968 24728 15020
rect 42800 14968 42852 15020
rect 46848 14968 46900 15020
rect 18604 14900 18656 14952
rect 45284 14943 45336 14952
rect 45284 14909 45293 14943
rect 45293 14909 45327 14943
rect 45327 14909 45336 14943
rect 45284 14900 45336 14909
rect 18420 14832 18472 14884
rect 19064 14764 19116 14816
rect 19340 14764 19392 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 2688 14356 2740 14408
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 17684 14356 17736 14408
rect 19984 14492 20036 14544
rect 19248 14467 19300 14476
rect 19248 14433 19257 14467
rect 19257 14433 19291 14467
rect 19291 14433 19300 14467
rect 19248 14424 19300 14433
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 22468 14424 22520 14476
rect 23388 14467 23440 14476
rect 23388 14433 23397 14467
rect 23397 14433 23431 14467
rect 23431 14433 23440 14467
rect 23388 14424 23440 14433
rect 17592 14288 17644 14340
rect 16856 14220 16908 14272
rect 47124 14356 47176 14408
rect 22100 14288 22152 14340
rect 21640 14220 21692 14272
rect 47308 14263 47360 14272
rect 47308 14229 47317 14263
rect 47317 14229 47351 14263
rect 47351 14229 47360 14263
rect 47308 14220 47360 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 17592 14016 17644 14068
rect 20628 14016 20680 14068
rect 22100 14059 22152 14068
rect 22100 14025 22109 14059
rect 22109 14025 22143 14059
rect 22143 14025 22152 14059
rect 22100 14016 22152 14025
rect 16856 13991 16908 14000
rect 16856 13957 16865 13991
rect 16865 13957 16899 13991
rect 16899 13957 16908 13991
rect 16856 13948 16908 13957
rect 16304 13880 16356 13932
rect 19064 13880 19116 13932
rect 21640 13880 21692 13932
rect 30472 13880 30524 13932
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 19616 13855 19668 13864
rect 19616 13821 19625 13855
rect 19625 13821 19659 13855
rect 19659 13821 19668 13855
rect 19616 13812 19668 13821
rect 21364 13812 21416 13864
rect 3424 13744 3476 13796
rect 15752 13744 15804 13796
rect 16304 13744 16356 13796
rect 18420 13744 18472 13796
rect 47768 13719 47820 13728
rect 47768 13685 47777 13719
rect 47777 13685 47811 13719
rect 47811 13685 47820 13719
rect 47768 13676 47820 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 14832 13472 14884 13524
rect 19616 13472 19668 13524
rect 47768 13336 47820 13388
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 17684 13268 17736 13320
rect 47308 13200 47360 13252
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 17224 13132 17276 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 22376 12860 22428 12912
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 3608 12656 3660 12708
rect 32036 12588 32088 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 22008 12384 22060 12436
rect 17224 12180 17276 12232
rect 45928 12180 45980 12232
rect 46480 12044 46532 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 46480 11203 46532 11212
rect 46480 11169 46489 11203
rect 46489 11169 46523 11203
rect 46523 11169 46532 11203
rect 46480 11160 46532 11169
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 2964 10956 3016 11008
rect 12440 10956 12492 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 47400 10616 47452 10668
rect 46296 10412 46348 10464
rect 47676 10455 47728 10464
rect 47676 10421 47685 10455
rect 47685 10421 47719 10455
rect 47719 10421 47728 10455
rect 47676 10412 47728 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 47676 10072 47728 10124
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 47952 9392 48004 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47768 8891 47820 8900
rect 47768 8857 47777 8891
rect 47777 8857 47811 8891
rect 47811 8857 47820 8891
rect 47768 8848 47820 8857
rect 29920 8780 29972 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 46848 8440 46900 8492
rect 18512 8236 18564 8288
rect 46848 8236 46900 8288
rect 47124 8236 47176 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3516 8032 3568 8084
rect 20720 8032 20772 8084
rect 19340 7896 19392 7948
rect 20168 7896 20220 7948
rect 45652 7896 45704 7948
rect 20168 7760 20220 7812
rect 20444 7760 20496 7812
rect 46204 7760 46256 7812
rect 46572 7803 46624 7812
rect 46572 7769 46581 7803
rect 46581 7769 46615 7803
rect 46615 7769 46624 7803
rect 47124 7939 47176 7948
rect 47124 7905 47133 7939
rect 47133 7905 47167 7939
rect 47167 7905 47176 7939
rect 47124 7896 47176 7905
rect 46572 7760 46624 7769
rect 47584 7760 47636 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 47584 7531 47636 7540
rect 47584 7497 47593 7531
rect 47593 7497 47627 7531
rect 47627 7497 47636 7531
rect 47584 7488 47636 7497
rect 46204 7352 46256 7404
rect 2044 7216 2096 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3332 6808 3384 6860
rect 23388 6808 23440 6860
rect 39396 6808 39448 6860
rect 47308 6851 47360 6860
rect 47308 6817 47317 6851
rect 47317 6817 47351 6851
rect 47351 6817 47360 6851
rect 47308 6808 47360 6817
rect 47216 6740 47268 6792
rect 6644 6604 6696 6656
rect 37740 6715 37792 6724
rect 37740 6681 37749 6715
rect 37749 6681 37783 6715
rect 37783 6681 37792 6715
rect 37740 6672 37792 6681
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 37740 6400 37792 6452
rect 43996 6400 44048 6452
rect 38476 6375 38528 6384
rect 38476 6341 38485 6375
rect 38485 6341 38519 6375
rect 38519 6341 38528 6375
rect 38476 6332 38528 6341
rect 39396 6375 39448 6384
rect 39396 6341 39405 6375
rect 39405 6341 39439 6375
rect 39439 6341 39448 6375
rect 39396 6332 39448 6341
rect 37740 6307 37792 6316
rect 37740 6273 37749 6307
rect 37749 6273 37783 6307
rect 37783 6273 37792 6307
rect 37740 6264 37792 6273
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 38384 6239 38436 6248
rect 38384 6205 38393 6239
rect 38393 6205 38427 6239
rect 38427 6205 38436 6239
rect 38384 6196 38436 6205
rect 39212 6196 39264 6248
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 37740 5355 37792 5364
rect 37740 5321 37749 5355
rect 37749 5321 37783 5355
rect 37783 5321 37792 5355
rect 37740 5312 37792 5321
rect 38476 5176 38528 5228
rect 39672 5219 39724 5228
rect 39672 5185 39681 5219
rect 39681 5185 39715 5219
rect 39715 5185 39724 5219
rect 39672 5176 39724 5185
rect 47952 5176 48004 5228
rect 26608 5040 26660 5092
rect 37372 5015 37424 5024
rect 37372 4981 37381 5015
rect 37381 4981 37415 5015
rect 37415 4981 37424 5015
rect 37372 4972 37424 4981
rect 39120 4972 39172 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 20076 4700 20128 4752
rect 26240 4700 26292 4752
rect 46296 4700 46348 4752
rect 3976 4632 4028 4684
rect 43260 4675 43312 4684
rect 43260 4641 43269 4675
rect 43269 4641 43303 4675
rect 43303 4641 43312 4675
rect 43260 4632 43312 4641
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 39120 4607 39172 4616
rect 39120 4573 39129 4607
rect 39129 4573 39163 4607
rect 39163 4573 39172 4607
rect 39120 4564 39172 4573
rect 40132 4564 40184 4616
rect 40868 4607 40920 4616
rect 40868 4573 40877 4607
rect 40877 4573 40911 4607
rect 40911 4573 40920 4607
rect 40868 4564 40920 4573
rect 47492 4632 47544 4684
rect 46848 4564 46900 4616
rect 15660 4496 15712 4548
rect 15844 4428 15896 4480
rect 16672 4428 16724 4480
rect 23388 4428 23440 4480
rect 24860 4428 24912 4480
rect 26240 4539 26292 4548
rect 26240 4505 26249 4539
rect 26249 4505 26283 4539
rect 26283 4505 26292 4539
rect 26240 4496 26292 4505
rect 26976 4496 27028 4548
rect 27712 4496 27764 4548
rect 39948 4496 40000 4548
rect 44088 4496 44140 4548
rect 38384 4428 38436 4480
rect 38660 4428 38712 4480
rect 40224 4471 40276 4480
rect 40224 4437 40233 4471
rect 40233 4437 40267 4471
rect 40267 4437 40276 4471
rect 40224 4428 40276 4437
rect 41052 4428 41104 4480
rect 46480 4428 46532 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 14464 4224 14516 4276
rect 20904 4224 20956 4276
rect 39488 4224 39540 4276
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 8116 4020 8168 4072
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 13360 4088 13412 4140
rect 13820 4088 13872 4140
rect 8208 4020 8260 4029
rect 15752 4020 15804 4072
rect 17500 4088 17552 4140
rect 18236 4088 18288 4140
rect 19432 4088 19484 4140
rect 20444 4131 20496 4140
rect 20444 4097 20453 4131
rect 20453 4097 20487 4131
rect 20487 4097 20496 4131
rect 20444 4088 20496 4097
rect 20812 4088 20864 4140
rect 21180 4088 21232 4140
rect 17224 4020 17276 4072
rect 17316 4020 17368 4072
rect 20168 4020 20220 4072
rect 20628 4020 20680 4072
rect 22284 4088 22336 4140
rect 28724 4088 28776 4140
rect 38660 4088 38712 4140
rect 40224 4156 40276 4208
rect 42892 4199 42944 4208
rect 42892 4165 42901 4199
rect 42901 4165 42935 4199
rect 42935 4165 42944 4199
rect 42892 4156 42944 4165
rect 43260 4156 43312 4208
rect 46388 4156 46440 4208
rect 46664 4156 46716 4208
rect 32220 4020 32272 4072
rect 44456 4131 44508 4140
rect 44456 4097 44465 4131
rect 44465 4097 44499 4131
rect 44499 4097 44508 4131
rect 44456 4088 44508 4097
rect 39580 4020 39632 4072
rect 41420 4063 41472 4072
rect 41420 4029 41429 4063
rect 41429 4029 41463 4063
rect 41463 4029 41472 4063
rect 41420 4020 41472 4029
rect 41512 4020 41564 4072
rect 45652 4020 45704 4072
rect 1584 3884 1636 3936
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 3792 3884 3844 3936
rect 21732 3952 21784 4004
rect 21916 3952 21968 4004
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 13728 3884 13780 3936
rect 15108 3884 15160 3936
rect 15936 3927 15988 3936
rect 15936 3893 15945 3927
rect 15945 3893 15979 3927
rect 15979 3893 15988 3927
rect 15936 3884 15988 3893
rect 17960 3884 18012 3936
rect 19248 3884 19300 3936
rect 20076 3884 20128 3936
rect 20720 3884 20772 3936
rect 22100 3927 22152 3936
rect 22100 3893 22109 3927
rect 22109 3893 22143 3927
rect 22143 3893 22152 3927
rect 22100 3884 22152 3893
rect 22192 3884 22244 3936
rect 39488 3952 39540 4004
rect 29460 3884 29512 3936
rect 36544 3884 36596 3936
rect 39580 3884 39632 3936
rect 44088 3884 44140 3936
rect 46296 3884 46348 3936
rect 47860 3927 47912 3936
rect 47860 3893 47869 3927
rect 47869 3893 47903 3927
rect 47903 3893 47912 3927
rect 47860 3884 47912 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8116 3723 8168 3732
rect 8116 3689 8125 3723
rect 8125 3689 8159 3723
rect 8159 3689 8168 3723
rect 8116 3680 8168 3689
rect 17500 3723 17552 3732
rect 1768 3544 1820 3596
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 6552 3476 6604 3528
rect 10416 3612 10468 3664
rect 12992 3612 13044 3664
rect 10692 3587 10744 3596
rect 1308 3408 1360 3460
rect 7288 3408 7340 3460
rect 9128 3476 9180 3528
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 15108 3587 15160 3596
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 13176 3408 13228 3460
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 2780 3340 2832 3349
rect 6736 3340 6788 3392
rect 9312 3340 9364 3392
rect 10416 3340 10468 3392
rect 13544 3476 13596 3528
rect 14004 3408 14056 3460
rect 15108 3553 15117 3587
rect 15117 3553 15151 3587
rect 15151 3553 15160 3587
rect 15108 3544 15160 3553
rect 15936 3544 15988 3596
rect 17500 3689 17509 3723
rect 17509 3689 17543 3723
rect 17543 3689 17552 3723
rect 17500 3680 17552 3689
rect 18328 3680 18380 3732
rect 19340 3680 19392 3732
rect 21732 3723 21784 3732
rect 16304 3612 16356 3664
rect 21180 3612 21232 3664
rect 19984 3544 20036 3596
rect 21732 3689 21741 3723
rect 21741 3689 21775 3723
rect 21775 3689 21784 3723
rect 21732 3680 21784 3689
rect 24860 3680 24912 3732
rect 39672 3680 39724 3732
rect 40132 3723 40184 3732
rect 40132 3689 40141 3723
rect 40141 3689 40175 3723
rect 40175 3689 40184 3723
rect 40132 3680 40184 3689
rect 40868 3680 40920 3732
rect 21364 3612 21416 3664
rect 30932 3612 30984 3664
rect 32956 3612 33008 3664
rect 36544 3612 36596 3664
rect 47860 3612 47912 3664
rect 16764 3476 16816 3528
rect 17960 3476 18012 3528
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 19340 3476 19392 3528
rect 20168 3476 20220 3528
rect 22192 3476 22244 3528
rect 16948 3408 17000 3460
rect 13360 3340 13412 3392
rect 13636 3340 13688 3392
rect 22284 3408 22336 3460
rect 23664 3544 23716 3596
rect 27712 3544 27764 3596
rect 32772 3544 32824 3596
rect 36452 3544 36504 3596
rect 41052 3587 41104 3596
rect 41052 3553 41061 3587
rect 41061 3553 41095 3587
rect 41095 3553 41104 3587
rect 41052 3544 41104 3553
rect 41420 3587 41472 3596
rect 41420 3553 41429 3587
rect 41429 3553 41463 3587
rect 41463 3553 41472 3587
rect 41420 3544 41472 3553
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 23388 3476 23440 3528
rect 39120 3519 39172 3528
rect 24584 3408 24636 3460
rect 26240 3451 26292 3460
rect 26240 3417 26249 3451
rect 26249 3417 26283 3451
rect 26283 3417 26292 3451
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 39948 3476 40000 3528
rect 40592 3476 40644 3528
rect 40868 3519 40920 3528
rect 40868 3485 40877 3519
rect 40877 3485 40911 3519
rect 40911 3485 40920 3519
rect 40868 3476 40920 3485
rect 26240 3408 26292 3417
rect 35716 3408 35768 3460
rect 45192 3519 45244 3528
rect 42800 3408 42852 3460
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 47400 3408 47452 3460
rect 48964 3408 49016 3460
rect 17592 3340 17644 3392
rect 18788 3340 18840 3392
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 20260 3340 20312 3392
rect 24768 3340 24820 3392
rect 33140 3383 33192 3392
rect 33140 3349 33149 3383
rect 33149 3349 33183 3383
rect 33183 3349 33192 3383
rect 33140 3340 33192 3349
rect 34428 3340 34480 3392
rect 42432 3340 42484 3392
rect 42984 3340 43036 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3884 3136 3936 3188
rect 16764 3179 16816 3188
rect 2780 3068 2832 3120
rect 6736 3111 6788 3120
rect 6736 3077 6745 3111
rect 6745 3077 6779 3111
rect 6779 3077 6788 3111
rect 6736 3068 6788 3077
rect 7288 3068 7340 3120
rect 9312 3111 9364 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 664 2932 716 2984
rect 6460 2932 6512 2984
rect 7748 2864 7800 2916
rect 9312 3077 9321 3111
rect 9321 3077 9355 3111
rect 9355 3077 9364 3111
rect 9312 3068 9364 3077
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 9036 2932 9088 2984
rect 12348 2932 12400 2984
rect 13452 3068 13504 3120
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 13452 2932 13504 2984
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 14188 2975 14240 2984
rect 13728 2932 13780 2941
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 15660 3068 15712 3120
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 18236 3179 18288 3188
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 17592 3068 17644 3120
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 19340 3136 19392 3188
rect 19432 3136 19484 3188
rect 20168 3179 20220 3188
rect 20168 3145 20177 3179
rect 20177 3145 20211 3179
rect 20211 3145 20220 3179
rect 20168 3136 20220 3145
rect 20812 3179 20864 3188
rect 20812 3145 20821 3179
rect 20821 3145 20855 3179
rect 20855 3145 20864 3179
rect 20812 3136 20864 3145
rect 20904 3136 20956 3188
rect 32772 3136 32824 3188
rect 33140 3111 33192 3120
rect 33140 3077 33149 3111
rect 33149 3077 33183 3111
rect 33183 3077 33192 3111
rect 33140 3068 33192 3077
rect 39120 3136 39172 3188
rect 40868 3136 40920 3188
rect 45100 3136 45152 3188
rect 47676 3136 47728 3188
rect 42984 3111 43036 3120
rect 42984 3077 42993 3111
rect 42993 3077 43027 3111
rect 43027 3077 43036 3111
rect 42984 3068 43036 3077
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 19984 3000 20036 3052
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20720 3043 20772 3052
rect 20076 3000 20128 3009
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 21916 3043 21968 3052
rect 21916 3009 21925 3043
rect 21925 3009 21959 3043
rect 21959 3009 21968 3043
rect 21916 3000 21968 3009
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 27068 3000 27120 3052
rect 29368 3000 29420 3052
rect 32956 3043 33008 3052
rect 32956 3009 32965 3043
rect 32965 3009 32999 3043
rect 32999 3009 33008 3043
rect 32956 3000 33008 3009
rect 39120 3000 39172 3052
rect 39948 3000 40000 3052
rect 18328 2932 18380 2984
rect 19340 2932 19392 2984
rect 21272 2932 21324 2984
rect 22100 2975 22152 2984
rect 22100 2941 22109 2975
rect 22109 2941 22143 2975
rect 22143 2941 22152 2975
rect 22100 2932 22152 2941
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 24768 2975 24820 2984
rect 24768 2941 24777 2975
rect 24777 2941 24811 2975
rect 24811 2941 24820 2975
rect 24768 2932 24820 2941
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 26424 2932 26476 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 39212 2975 39264 2984
rect 39212 2941 39221 2975
rect 39221 2941 39255 2975
rect 39255 2941 39264 2975
rect 39212 2932 39264 2941
rect 41512 3000 41564 3052
rect 42800 3043 42852 3052
rect 42800 3009 42809 3043
rect 42809 3009 42843 3043
rect 42843 3009 42852 3043
rect 42800 3000 42852 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 48320 3000 48372 3052
rect 40592 2975 40644 2984
rect 40592 2941 40601 2975
rect 40601 2941 40635 2975
rect 40635 2941 40644 2975
rect 40592 2932 40644 2941
rect 41696 2932 41748 2984
rect 43168 2932 43220 2984
rect 47676 2932 47728 2984
rect 7104 2796 7156 2848
rect 8208 2796 8260 2848
rect 41420 2864 41472 2916
rect 12992 2796 13044 2848
rect 14096 2796 14148 2848
rect 15752 2796 15804 2848
rect 20904 2796 20956 2848
rect 33140 2796 33192 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2872 2592 2924 2644
rect 4620 2592 4672 2644
rect 7196 2592 7248 2644
rect 10508 2592 10560 2644
rect 13820 2592 13872 2644
rect 14004 2592 14056 2644
rect 20444 2592 20496 2644
rect 20536 2592 20588 2644
rect 22192 2592 22244 2644
rect 23664 2592 23716 2644
rect 25044 2592 25096 2644
rect 26240 2635 26292 2644
rect 26240 2601 26249 2635
rect 26249 2601 26283 2635
rect 26283 2601 26292 2635
rect 26240 2592 26292 2601
rect 28816 2592 28868 2644
rect 33140 2592 33192 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 39120 2635 39172 2644
rect 39120 2601 39129 2635
rect 39129 2601 39163 2635
rect 39163 2601 39172 2635
rect 39120 2592 39172 2601
rect 41696 2635 41748 2644
rect 41696 2601 41705 2635
rect 41705 2601 41739 2635
rect 41739 2601 41748 2635
rect 41696 2592 41748 2601
rect 42524 2635 42576 2644
rect 42524 2601 42533 2635
rect 42533 2601 42567 2635
rect 42567 2601 42576 2635
rect 42524 2592 42576 2601
rect 44456 2592 44508 2644
rect 37372 2524 37424 2576
rect 43076 2524 43128 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 27252 2499 27304 2508
rect 5172 2388 5224 2440
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 16120 2388 16172 2440
rect 20260 2388 20312 2440
rect 23204 2388 23256 2440
rect 26424 2431 26476 2440
rect 26424 2397 26433 2431
rect 26433 2397 26467 2431
rect 26467 2397 26476 2431
rect 26424 2388 26476 2397
rect 26516 2388 26568 2440
rect 27252 2465 27261 2499
rect 27261 2465 27295 2499
rect 27295 2465 27304 2499
rect 27252 2456 27304 2465
rect 34244 2456 34296 2508
rect 27896 2388 27948 2440
rect 28356 2388 28408 2440
rect 29644 2388 29696 2440
rect 35440 2388 35492 2440
rect 2596 2252 2648 2304
rect 8392 2320 8444 2372
rect 15476 2320 15528 2372
rect 20628 2320 20680 2372
rect 21916 2320 21968 2372
rect 24492 2320 24544 2372
rect 32404 2320 32456 2372
rect 39948 2388 40000 2440
rect 41236 2388 41288 2440
rect 42892 2456 42944 2508
rect 46756 2456 46808 2508
rect 43812 2388 43864 2440
rect 36084 2320 36136 2372
rect 38016 2320 38068 2372
rect 39396 2320 39448 2372
rect 40592 2320 40644 2372
rect 47032 2388 47084 2440
rect 48044 2388 48096 2440
rect 12348 2252 12400 2304
rect 25228 2252 25280 2304
rect 29736 2295 29788 2304
rect 29736 2261 29745 2295
rect 29745 2261 29779 2295
rect 29779 2261 29788 2295
rect 29736 2252 29788 2261
rect 38476 2252 38528 2304
rect 46756 2320 46808 2372
rect 41788 2252 41840 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 29736 1980 29788 2032
rect 42524 1980 42576 2032
rect 32864 1912 32916 1964
rect 41788 1912 41840 1964
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 32 20874 60 49200
rect 1858 47696 1914 47705
rect 1858 47631 1914 47640
rect 1872 46646 1900 47631
rect 1964 47054 1992 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2608 46918 2636 49200
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3514 47016 3570 47025
rect 3514 46951 3570 46960
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 2872 46912 2924 46918
rect 2872 46854 2924 46860
rect 1860 46640 1912 46646
rect 1860 46582 1912 46588
rect 2044 46436 2096 46442
rect 2044 46378 2096 46384
rect 1400 46368 1452 46374
rect 1400 46310 1452 46316
rect 1412 46034 1440 46310
rect 1400 46028 1452 46034
rect 1400 45970 1452 45976
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1492 43240 1544 43246
rect 1492 43182 1544 43188
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1398 33416 1454 33425
rect 1398 33351 1454 33360
rect 1412 32978 1440 33351
rect 1400 32972 1452 32978
rect 1400 32914 1452 32920
rect 1504 26234 1532 43182
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1584 41540 1636 41546
rect 1858 41511 1914 41520
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35465 1624 35634
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1964 34066 1992 40326
rect 1952 34060 2004 34066
rect 1952 34002 2004 34008
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1596 32745 1624 33458
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1676 32360 1728 32366
rect 1676 32302 1728 32308
rect 1688 32026 1716 32302
rect 1676 32020 1728 32026
rect 1676 31962 1728 31968
rect 2056 26586 2084 46378
rect 2778 46336 2834 46345
rect 2778 46271 2834 46280
rect 2792 46034 2820 46271
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2228 45892 2280 45898
rect 2228 45834 2280 45840
rect 2240 45626 2268 45834
rect 2228 45620 2280 45626
rect 2228 45562 2280 45568
rect 2320 45484 2372 45490
rect 2320 45426 2372 45432
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2136 36168 2188 36174
rect 2136 36110 2188 36116
rect 2044 26580 2096 26586
rect 2044 26522 2096 26528
rect 1504 26206 1624 26234
rect 20 20868 72 20874
rect 20 20810 72 20816
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1596 17338 1624 26206
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1964 6914 1992 16050
rect 2056 7274 2084 25094
rect 2148 18766 2176 36110
rect 2228 35488 2280 35494
rect 2228 35430 2280 35436
rect 2240 33522 2268 35430
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 2228 32360 2280 32366
rect 2228 32302 2280 32308
rect 2240 32026 2268 32302
rect 2228 32020 2280 32026
rect 2228 31962 2280 31968
rect 2332 31822 2360 45426
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2780 33312 2832 33318
rect 2780 33254 2832 33260
rect 2792 33114 2820 33254
rect 2780 33108 2832 33114
rect 2780 33050 2832 33056
rect 2688 32904 2740 32910
rect 2688 32846 2740 32852
rect 2700 31890 2728 32846
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2792 32065 2820 32302
rect 2778 32056 2834 32065
rect 2778 31991 2834 32000
rect 2688 31884 2740 31890
rect 2688 31826 2740 31832
rect 2320 31816 2372 31822
rect 2320 31758 2372 31764
rect 2884 21078 2912 46854
rect 3422 44976 3478 44985
rect 3422 44911 3478 44920
rect 3330 31376 3386 31385
rect 3330 31311 3386 31320
rect 3344 28082 3372 31311
rect 3332 28076 3384 28082
rect 3332 28018 3384 28024
rect 2872 21072 2924 21078
rect 2872 21014 2924 21020
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2976 19825 3004 20538
rect 3436 20058 3464 44911
rect 3528 23866 3556 46951
rect 3896 46646 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 47054 4752 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7328 49314
rect 7074 49200 7186 49286
rect 5828 47054 5856 49200
rect 7300 47054 7328 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 4712 47048 4764 47054
rect 4712 46990 4764 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7288 47048 7340 47054
rect 7288 46990 7340 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 4988 46980 5040 46986
rect 4988 46922 5040 46928
rect 6644 46980 6696 46986
rect 6644 46922 6696 46928
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3988 46170 4016 46446
rect 3976 46164 4028 46170
rect 3976 46106 4028 46112
rect 3698 43616 3754 43625
rect 3698 43551 3754 43560
rect 3606 28656 3662 28665
rect 3606 28591 3662 28600
rect 3620 28218 3648 28591
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3620 23186 3648 28018
rect 3608 23180 3660 23186
rect 3608 23122 3660 23128
rect 3712 22506 3740 43551
rect 3882 39536 3938 39545
rect 3882 39471 3938 39480
rect 3792 33448 3844 33454
rect 3792 33390 3844 33396
rect 3804 33114 3832 33390
rect 3792 33108 3844 33114
rect 3792 33050 3844 33056
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3700 22500 3752 22506
rect 3700 22442 3752 22448
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 2962 19816 3018 19825
rect 2962 19751 3018 19760
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 3422 18456 3478 18465
rect 3422 18391 3424 18400
rect 3476 18391 3478 18400
rect 3424 18362 3476 18368
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3436 17105 3464 17138
rect 3422 17096 3478 17105
rect 3422 17031 3478 17040
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1964 6886 2084 6914
rect 2056 4146 2084 6886
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3402
rect 1596 2514 1624 3878
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3058 1808 3538
rect 2700 3534 2728 14350
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 13705 3464 13738
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3528 11642 3556 16458
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3436 11614 3556 11642
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10305 3004 10950
rect 2962 10296 3018 10305
rect 2962 10231 3018 10240
rect 3330 6896 3386 6905
rect 3330 6831 3332 6840
rect 3384 6831 3386 6840
rect 3332 6802 3384 6808
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2792 3126 2820 3334
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2884 2650 2912 3878
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2884 785 2912 2450
rect 3436 1465 3464 11614
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3528 7585 3556 8026
rect 3514 7576 3570 7585
rect 3514 7511 3570 7520
rect 3620 6914 3648 12650
rect 3528 6886 3648 6914
rect 3528 3505 3556 6886
rect 3804 3942 3832 31758
rect 3896 23798 3924 39471
rect 3884 23792 3936 23798
rect 3884 23734 3936 23740
rect 4080 6914 4108 46922
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4632 31890 4660 33390
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4620 30388 4672 30394
rect 4620 30330 4672 30336
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3988 6886 4108 6914
rect 3988 4690 4016 6886
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3514 3496 3570 3505
rect 3514 3431 3570 3440
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 3896 800 3924 3130
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 2650 4660 30330
rect 5000 18970 5028 46922
rect 5172 46504 5224 46510
rect 5172 46446 5224 46452
rect 5184 46170 5212 46446
rect 5172 46164 5224 46170
rect 5172 46106 5224 46112
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 5460 15570 5488 31826
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 6656 6662 6684 46922
rect 7472 46912 7524 46918
rect 7472 46854 7524 46860
rect 7484 27606 7512 46854
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 8312 29034 8340 45526
rect 9508 36378 9536 46922
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 46034 10456 46310
rect 10980 46034 11008 49200
rect 11624 47054 11652 49200
rect 12268 47054 12296 49200
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 12256 47048 12308 47054
rect 12256 46990 12308 46996
rect 12624 47048 12676 47054
rect 12624 46990 12676 46996
rect 11796 46980 11848 46986
rect 11796 46922 11848 46928
rect 10416 46028 10468 46034
rect 10416 45970 10468 45976
rect 10968 46028 11020 46034
rect 10968 45970 11020 45976
rect 10600 45892 10652 45898
rect 10600 45834 10652 45840
rect 10612 45626 10640 45834
rect 10600 45620 10652 45626
rect 10600 45562 10652 45568
rect 11808 36854 11836 46922
rect 12636 38418 12664 46990
rect 12912 46918 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 14200 47954 14228 49200
rect 14200 47926 14320 47954
rect 13740 47110 13860 47138
rect 13832 47054 13860 47110
rect 13820 47048 13872 47054
rect 13820 46990 13872 46996
rect 12900 46912 12952 46918
rect 12900 46854 12952 46860
rect 14292 46510 14320 47926
rect 15488 47138 15516 49200
rect 15488 47110 16160 47138
rect 15568 46980 15620 46986
rect 15568 46922 15620 46928
rect 14648 46912 14700 46918
rect 14648 46854 14700 46860
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 14200 46170 14228 46446
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 14108 41138 14136 45902
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 12624 38412 12676 38418
rect 12624 38354 12676 38360
rect 14660 37262 14688 46854
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 11796 36848 11848 36854
rect 11796 36790 11848 36796
rect 9496 36372 9548 36378
rect 9496 36314 9548 36320
rect 14200 35894 14228 37198
rect 14200 35866 14412 35894
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14108 29646 14136 30194
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 12440 29232 12492 29238
rect 12440 29174 12492 29180
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 10704 28762 10732 29038
rect 11072 28966 11100 29106
rect 11520 29096 11572 29102
rect 11520 29038 11572 29044
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 10692 28756 10744 28762
rect 10692 28698 10744 28704
rect 11532 28694 11560 29038
rect 12164 28960 12216 28966
rect 12164 28902 12216 28908
rect 11520 28688 11572 28694
rect 11520 28630 11572 28636
rect 11796 28620 11848 28626
rect 11796 28562 11848 28568
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 11244 28552 11296 28558
rect 11244 28494 11296 28500
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 9968 28082 9996 28494
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 9968 26382 9996 28018
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 10520 27538 10548 27814
rect 10508 27532 10560 27538
rect 10508 27474 10560 27480
rect 11256 27130 11284 28494
rect 11336 28416 11388 28422
rect 11336 28358 11388 28364
rect 11348 27674 11376 28358
rect 11440 28014 11468 28494
rect 11808 28422 11836 28562
rect 11980 28484 12032 28490
rect 11980 28426 12032 28432
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11808 28218 11836 28358
rect 11796 28212 11848 28218
rect 11716 28172 11796 28200
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 11520 27940 11572 27946
rect 11520 27882 11572 27888
rect 11532 27674 11560 27882
rect 11336 27668 11388 27674
rect 11336 27610 11388 27616
rect 11520 27668 11572 27674
rect 11520 27610 11572 27616
rect 11532 27282 11560 27610
rect 11440 27254 11560 27282
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9968 23730 9996 26318
rect 10232 26240 10284 26246
rect 10232 26182 10284 26188
rect 10244 25362 10272 26182
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10520 25362 10548 25638
rect 10232 25356 10284 25362
rect 10232 25298 10284 25304
rect 10508 25356 10560 25362
rect 10508 25298 10560 25304
rect 10980 24818 11008 25774
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 10600 24608 10652 24614
rect 10600 24550 10652 24556
rect 10612 24274 10640 24550
rect 10600 24268 10652 24274
rect 10600 24210 10652 24216
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10336 23798 10364 24142
rect 10324 23792 10376 23798
rect 10324 23734 10376 23740
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 9968 23118 9996 23666
rect 11348 23322 11376 24686
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8404 22234 8432 22510
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 9876 22098 9904 22918
rect 9968 22778 9996 23054
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 7932 21412 7984 21418
rect 7932 21354 7984 21360
rect 7944 17202 7972 21354
rect 8956 21350 8984 21966
rect 10796 21962 10824 22918
rect 11072 22506 11100 23054
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 11256 22166 11284 22646
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11348 22098 11376 22578
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 10784 21956 10836 21962
rect 10784 21898 10836 21904
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8956 20942 8984 21286
rect 9048 21146 9076 21422
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10704 19990 10732 20334
rect 10692 19984 10744 19990
rect 10692 19926 10744 19932
rect 11348 19854 11376 22034
rect 11440 21622 11468 27254
rect 11716 27062 11744 28172
rect 11796 28154 11848 28160
rect 11992 28082 12020 28426
rect 12176 28150 12204 28902
rect 12452 28762 12480 29174
rect 12440 28756 12492 28762
rect 12440 28698 12492 28704
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 12164 28144 12216 28150
rect 12164 28086 12216 28092
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 11888 27668 11940 27674
rect 11888 27610 11940 27616
rect 11704 27056 11756 27062
rect 11704 26998 11756 27004
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11532 26518 11560 26930
rect 11520 26512 11572 26518
rect 11520 26454 11572 26460
rect 11716 26234 11744 26998
rect 11900 26994 11928 27610
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11992 26382 12020 28018
rect 12176 26926 12204 28086
rect 12360 28082 12388 28494
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 13188 28218 13216 28426
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12624 27872 12676 27878
rect 12624 27814 12676 27820
rect 12636 27402 12664 27814
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 13832 26994 13860 28086
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13912 27464 13964 27470
rect 13912 27406 13964 27412
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 12164 26920 12216 26926
rect 12164 26862 12216 26868
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 11716 26206 11836 26234
rect 11808 25906 11836 26206
rect 12268 26042 12296 26454
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 13832 25974 13860 26182
rect 13820 25968 13872 25974
rect 13820 25910 13872 25916
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11808 25362 11836 25842
rect 13924 25838 13952 27406
rect 14016 27402 14044 28018
rect 14108 27606 14136 28494
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14292 27674 14320 28018
rect 14280 27668 14332 27674
rect 14280 27610 14332 27616
rect 14096 27600 14148 27606
rect 14096 27542 14148 27548
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 14016 26450 14044 27338
rect 14108 26518 14136 27406
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14096 26512 14148 26518
rect 14096 26454 14148 26460
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 14108 26382 14136 26454
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14200 25974 14228 26726
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 14292 25702 14320 26318
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11624 24818 11652 25230
rect 14108 25226 14136 25638
rect 14096 25220 14148 25226
rect 14096 25162 14148 25168
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12360 24206 12388 24686
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11900 23746 11928 24006
rect 11808 23718 11928 23746
rect 11808 23662 11836 23718
rect 11796 23656 11848 23662
rect 11796 23598 11848 23604
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11624 21894 11652 23054
rect 11808 23050 11836 23598
rect 11992 23322 12020 23598
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 12268 22982 12296 23258
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 12268 22778 12296 22918
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11428 21616 11480 21622
rect 11428 21558 11480 21564
rect 11716 21554 11744 22374
rect 11900 22030 11928 22714
rect 12164 22704 12216 22710
rect 12164 22646 12216 22652
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11900 21554 11928 21830
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 21078 11560 21286
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11808 20534 11836 20742
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11992 19854 12020 22374
rect 12176 21690 12204 22646
rect 12360 22438 12388 24142
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13096 22506 13124 22918
rect 13832 22642 13860 23462
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13084 22500 13136 22506
rect 13084 22442 13136 22448
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12176 21350 12204 21626
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 12084 19990 12112 20470
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10888 19378 10916 19722
rect 11992 19378 12020 19790
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 10428 18834 10456 19110
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 11716 18698 11744 19110
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 10980 18222 11008 18634
rect 12176 18630 12204 21286
rect 12360 18766 12388 21490
rect 12452 20398 12480 21558
rect 12820 21418 12848 21966
rect 12900 21956 12952 21962
rect 12900 21898 12952 21904
rect 12912 21690 12940 21898
rect 13924 21894 13952 23598
rect 14108 23186 14136 25162
rect 14384 24070 14412 35866
rect 15580 31754 15608 46922
rect 16132 45554 16160 47110
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49314 21354 50000
rect 21242 49286 21680 49314
rect 21242 49200 21354 49286
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 17420 45554 17448 49200
rect 18708 46918 18736 49200
rect 19996 46918 20024 49200
rect 20076 46980 20128 46986
rect 20076 46922 20128 46928
rect 18696 46912 18748 46918
rect 18696 46854 18748 46860
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19616 46504 19668 46510
rect 19616 46446 19668 46452
rect 19628 46170 19656 46446
rect 19616 46164 19668 46170
rect 19616 46106 19668 46112
rect 18420 45960 18472 45966
rect 18420 45902 18472 45908
rect 18604 45960 18656 45966
rect 18604 45902 18656 45908
rect 16132 45526 16528 45554
rect 15488 31726 15608 31754
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 14936 29714 14964 29990
rect 14924 29708 14976 29714
rect 14924 29650 14976 29656
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14476 29238 14504 29446
rect 14464 29232 14516 29238
rect 14464 29174 14516 29180
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 14476 28762 14504 29038
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14476 28218 14504 28698
rect 14752 28422 14780 29582
rect 14832 29096 14884 29102
rect 14832 29038 14884 29044
rect 14844 28966 14872 29038
rect 14832 28960 14884 28966
rect 14832 28902 14884 28908
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 14752 28082 14780 28358
rect 14844 28150 14872 28902
rect 15384 28484 15436 28490
rect 15384 28426 15436 28432
rect 15396 28218 15424 28426
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 14832 28144 14884 28150
rect 14832 28086 14884 28092
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 15108 28076 15160 28082
rect 15108 28018 15160 28024
rect 14832 27872 14884 27878
rect 14832 27814 14884 27820
rect 14844 27470 14872 27814
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14740 26308 14792 26314
rect 14740 26250 14792 26256
rect 14752 25294 14780 26250
rect 14844 25294 14872 27406
rect 15120 26994 15148 28018
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 14740 25288 14792 25294
rect 14740 25230 14792 25236
rect 14832 25288 14884 25294
rect 14832 25230 14884 25236
rect 14752 24954 14780 25230
rect 14844 25158 14872 25230
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23798 14412 24006
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14568 23322 14596 24686
rect 14752 23322 14780 24754
rect 14936 24206 14964 25774
rect 15028 25226 15056 26318
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 15120 25226 15148 25638
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14936 23730 14964 24142
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14096 23180 14148 23186
rect 14096 23122 14148 23128
rect 14280 23044 14332 23050
rect 14280 22986 14332 22992
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14292 22234 14320 22986
rect 14476 22710 14504 22986
rect 14752 22778 14780 23258
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 12900 21684 12952 21690
rect 12900 21626 12952 21632
rect 14108 21418 14136 21966
rect 14476 21962 14504 22374
rect 14936 22166 14964 23462
rect 14924 22160 14976 22166
rect 14924 22102 14976 22108
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14936 21554 14964 22102
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 12820 20874 12848 21354
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14292 21010 14320 21286
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 19378 12940 19654
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13188 18902 13216 19246
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 18290 12204 18566
rect 12360 18358 12388 18702
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 13280 18290 13308 19722
rect 14108 19514 14136 20878
rect 14384 19854 14412 21286
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16600 11100 17070
rect 11060 16594 11112 16600
rect 11060 16536 11112 16542
rect 11532 16114 11560 18226
rect 13280 17678 13308 18226
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16658 11928 16934
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16182 11744 16390
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12452 11014 12480 15982
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 13372 4146 13400 18566
rect 13832 18222 13860 18838
rect 14108 18766 14136 19450
rect 14476 19446 14504 19654
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14384 18630 14412 19246
rect 14752 18766 14780 19314
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17202 13492 17478
rect 13832 17270 13860 18022
rect 14384 17882 14412 18566
rect 14476 18358 14504 18634
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16794 14412 16934
rect 14568 16794 14596 18158
rect 14660 17882 14688 18158
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14660 16402 14688 17682
rect 14752 17610 14780 18702
rect 15028 18630 15056 25162
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24750 15240 25094
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15212 22574 15240 24686
rect 15304 23730 15332 26930
rect 15488 25362 15516 31726
rect 16500 29714 16528 45526
rect 16776 45526 17448 45554
rect 16488 29708 16540 29714
rect 16488 29650 16540 29656
rect 16776 29034 16804 45526
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 18156 32434 18184 32846
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 18144 31816 18196 31822
rect 18144 31758 18196 31764
rect 18156 31346 18184 31758
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 16764 29028 16816 29034
rect 16764 28970 16816 28976
rect 16868 28762 16896 29038
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 17328 28558 17356 30194
rect 17408 30184 17460 30190
rect 17408 30126 17460 30132
rect 17592 30184 17644 30190
rect 17592 30126 17644 30132
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 16592 28218 16620 28494
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16580 28008 16632 28014
rect 16580 27950 16632 27956
rect 16592 26382 16620 27950
rect 16580 26376 16632 26382
rect 16856 26376 16908 26382
rect 16632 26336 16804 26364
rect 16580 26318 16632 26324
rect 16672 26240 16724 26246
rect 16592 26188 16672 26194
rect 16592 26182 16724 26188
rect 16592 26166 16712 26182
rect 16592 25974 16620 26166
rect 16580 25968 16632 25974
rect 16580 25910 16632 25916
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 15580 24818 15608 25434
rect 15672 24954 15700 25774
rect 16592 25158 16620 25910
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15856 24818 15884 25094
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15304 23050 15332 23666
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 15476 23044 15528 23050
rect 15476 22986 15528 22992
rect 15488 22574 15516 22986
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15660 22500 15712 22506
rect 15660 22442 15712 22448
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15488 19990 15516 20334
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14936 18222 14964 18566
rect 15120 18290 15148 19790
rect 15672 19310 15700 22442
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 14936 17542 14964 18158
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 15028 17746 15056 18090
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 17746 15516 18022
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14936 16590 14964 17478
rect 15028 17134 15056 17546
rect 15672 17202 15700 18226
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 15028 16658 15056 17070
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14740 16448 14792 16454
rect 14660 16396 14740 16402
rect 14660 16390 14792 16396
rect 14660 16374 14780 16390
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 15570 14596 15846
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14752 15094 14780 16374
rect 14832 15428 14884 15434
rect 14832 15370 14884 15376
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14844 14958 14872 15370
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14936 14890 14964 16526
rect 15672 16046 15700 17138
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 15162 15608 15370
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15672 15026 15700 15982
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 15764 13802 15792 23122
rect 15856 22642 15884 24754
rect 16684 24410 16712 25230
rect 16776 24818 16804 26336
rect 16856 26318 16908 26324
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16868 25906 16896 26318
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16960 25786 16988 26318
rect 17132 26240 17184 26246
rect 17132 26182 17184 26188
rect 17144 25906 17172 26182
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 16868 25758 16988 25786
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 16868 24206 16896 25758
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 16960 25362 16988 25638
rect 17420 25498 17448 30126
rect 17604 28762 17632 30126
rect 17592 28756 17644 28762
rect 17592 28698 17644 28704
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 17592 28212 17644 28218
rect 17592 28154 17644 28160
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 16948 25356 17000 25362
rect 16948 25298 17000 25304
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24954 17080 25094
rect 17040 24948 17092 24954
rect 17040 24890 17092 24896
rect 16948 24880 17000 24886
rect 16948 24822 17000 24828
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16408 23186 16436 23598
rect 16856 23316 16908 23322
rect 16960 23304 16988 24822
rect 17604 24290 17632 28154
rect 17604 24274 17816 24290
rect 17604 24268 17828 24274
rect 17604 24262 17776 24268
rect 17604 23866 17632 24262
rect 17776 24210 17828 24216
rect 17880 24070 17908 28494
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18156 25838 18184 26182
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18248 24818 18276 25230
rect 18328 25220 18380 25226
rect 18328 25162 18380 25168
rect 18340 24818 18368 25162
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17696 23866 17724 24006
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 16908 23276 16988 23304
rect 16856 23258 16908 23264
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16960 22930 16988 23276
rect 17144 23050 17172 23462
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 16592 22234 16620 22918
rect 16868 22642 16896 22918
rect 16960 22902 17172 22930
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 17040 22568 17092 22574
rect 17040 22510 17092 22516
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16592 22094 16620 22170
rect 16592 22066 16712 22094
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 21554 16252 21830
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16224 20466 16252 21490
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16592 20602 16620 20810
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14476 4282 14504 4558
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 3058 6592 3470
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3126 6776 3334
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5184 800 5212 2382
rect 6472 800 6500 2926
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 800 7144 2790
rect 7208 2650 7236 4014
rect 8128 3738 8156 4014
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7300 3126 7328 3402
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7760 800 7788 2858
rect 8220 2854 8248 4014
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 3058 9168 3470
rect 10428 3398 10456 3606
rect 10704 3602 10732 3878
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 9324 3126 9352 3334
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9048 800 9076 2926
rect 10520 2650 10548 3470
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10980 800 11008 3538
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 2310 12388 2926
rect 13004 2854 13032 3606
rect 13544 3528 13596 3534
rect 13176 3460 13228 3466
rect 13280 3454 13492 3482
rect 13544 3470 13596 3476
rect 13280 3448 13308 3454
rect 13228 3420 13308 3448
rect 13176 3402 13228 3408
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13372 2446 13400 3334
rect 13464 3126 13492 3454
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13556 3058 13584 3470
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13452 2984 13504 2990
rect 13648 2938 13676 3334
rect 13740 2990 13768 3878
rect 13504 2932 13676 2938
rect 13452 2926 13676 2932
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13464 2910 13676 2926
rect 13832 2650 13860 4082
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 14016 2650 14044 3402
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14108 2446 14136 2790
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 14200 800 14228 2926
rect 14844 800 14872 13466
rect 16132 12434 16160 20334
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17678 16620 18022
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16684 17066 16712 22066
rect 17052 21690 17080 22510
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16776 19854 16804 20402
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 19922 17080 20198
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16868 19446 16896 19858
rect 16856 19440 16908 19446
rect 16856 19382 16908 19388
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18290 16804 18566
rect 16868 18358 16896 19382
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16868 17882 16896 18294
rect 17040 18284 17092 18290
rect 17144 18272 17172 22902
rect 17604 22098 17632 23802
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17328 21010 17356 21490
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17880 20466 17908 24006
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17972 22030 18000 23666
rect 18432 23050 18460 45902
rect 18616 45554 18644 45902
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 18524 45526 18644 45554
rect 18524 45490 18552 45526
rect 18512 45484 18564 45490
rect 18512 45426 18564 45432
rect 18524 38282 18552 45426
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 19444 38350 19472 38898
rect 19432 38344 19484 38350
rect 19432 38286 19484 38292
rect 18512 38276 18564 38282
rect 18512 38218 18564 38224
rect 18524 31822 18552 38218
rect 19444 38010 19472 38286
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19432 38004 19484 38010
rect 19432 37946 19484 37952
rect 19444 37874 19472 37946
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 19432 37868 19484 37874
rect 19432 37810 19484 37816
rect 19616 37868 19668 37874
rect 19616 37810 19668 37816
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 18616 34542 18644 35566
rect 18604 34536 18656 34542
rect 18604 34478 18656 34484
rect 18616 32910 18644 34478
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18524 31414 18552 31622
rect 18512 31408 18564 31414
rect 18512 31350 18564 31356
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18524 28558 18552 29106
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18880 26308 18932 26314
rect 18880 26250 18932 26256
rect 18892 26042 18920 26250
rect 18880 26036 18932 26042
rect 18880 25978 18932 25984
rect 19076 24206 19104 37810
rect 19432 37732 19484 37738
rect 19432 37674 19484 37680
rect 19156 36236 19208 36242
rect 19156 36178 19208 36184
rect 19168 35630 19196 36178
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 19352 30258 19380 36110
rect 19444 36106 19472 37674
rect 19628 37466 19656 37810
rect 19616 37460 19668 37466
rect 19616 37402 19668 37408
rect 19984 37460 20036 37466
rect 19984 37402 20036 37408
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36174 20024 37402
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19432 36100 19484 36106
rect 19432 36042 19484 36048
rect 19444 32774 19472 36042
rect 19984 36032 20036 36038
rect 19984 35974 20036 35980
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19996 35766 20024 35974
rect 19984 35760 20036 35766
rect 19984 35702 20036 35708
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19616 34672 19668 34678
rect 19616 34614 19668 34620
rect 19628 34202 19656 34614
rect 19616 34196 19668 34202
rect 19616 34138 19668 34144
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 19996 32842 20024 33254
rect 19984 32836 20036 32842
rect 19984 32778 20036 32784
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19984 32564 20036 32570
rect 19984 32506 20036 32512
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19444 32026 19472 32438
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19996 31822 20024 32506
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 19168 29034 19196 29582
rect 19352 29170 19380 30194
rect 19800 30048 19852 30054
rect 19800 29990 19852 29996
rect 19812 29578 19840 29990
rect 19800 29572 19852 29578
rect 19800 29514 19852 29520
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19984 29096 20036 29102
rect 19984 29038 20036 29044
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19168 28626 19196 28970
rect 19156 28620 19208 28626
rect 19156 28562 19208 28568
rect 19168 28150 19196 28562
rect 19996 28490 20024 29038
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19352 28150 19380 28358
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19156 28144 19208 28150
rect 19156 28086 19208 28092
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19996 25974 20024 26318
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19352 25498 19380 25842
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19340 25492 19392 25498
rect 19340 25434 19392 25440
rect 19536 25362 19564 25774
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19076 23662 19104 24142
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 19260 23322 19288 25230
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19352 23866 19380 24346
rect 20088 24177 20116 46922
rect 20640 46510 20668 49200
rect 20720 47048 20772 47054
rect 20720 46990 20772 46996
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20732 46102 20760 46990
rect 20720 46096 20772 46102
rect 20720 46038 20772 46044
rect 21652 45966 21680 49286
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49314 27150 50000
rect 26712 49286 27150 49314
rect 22284 47184 22336 47190
rect 22284 47126 22336 47132
rect 21824 46912 21876 46918
rect 21824 46854 21876 46860
rect 21640 45960 21692 45966
rect 21640 45902 21692 45908
rect 20168 39568 20220 39574
rect 20168 39510 20220 39516
rect 20180 39030 20208 39510
rect 21836 39030 21864 46854
rect 20168 39024 20220 39030
rect 20168 38966 20220 38972
rect 20444 39024 20496 39030
rect 20444 38966 20496 38972
rect 21824 39024 21876 39030
rect 21824 38966 21876 38972
rect 20168 38480 20220 38486
rect 20168 38422 20220 38428
rect 20180 38282 20208 38422
rect 20168 38276 20220 38282
rect 20168 38218 20220 38224
rect 20074 24168 20130 24177
rect 20074 24103 20130 24112
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 20088 23798 20116 24006
rect 20076 23792 20128 23798
rect 19522 23760 19578 23769
rect 19340 23724 19392 23730
rect 19392 23704 19522 23712
rect 20076 23734 20128 23740
rect 19392 23695 19578 23704
rect 19392 23684 19564 23695
rect 19340 23666 19392 23672
rect 19338 23624 19394 23633
rect 19338 23559 19394 23568
rect 19352 23526 19380 23559
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19352 23118 19380 23190
rect 19340 23112 19392 23118
rect 20076 23112 20128 23118
rect 19392 23072 19472 23100
rect 19340 23054 19392 23060
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17972 21554 18000 21966
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 18248 21486 18276 22170
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17972 20534 18000 20946
rect 18248 20534 18276 21286
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 18616 20398 18644 21422
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 17972 19514 18000 20334
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17092 18244 17172 18272
rect 17040 18226 17092 18232
rect 17052 17882 17080 18226
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16672 17060 16724 17066
rect 16672 17002 16724 17008
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16316 15094 16344 15302
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16316 13938 16344 15030
rect 16684 14414 16712 17002
rect 16960 16794 16988 17070
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15570 16896 15846
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17144 15162 17172 15370
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16868 14006 16896 14214
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16316 13326 16344 13738
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 17236 13190 17264 16662
rect 18432 16658 18460 17682
rect 18616 16726 18644 20334
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18432 16114 18460 16594
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15434 17632 15846
rect 18616 15638 18644 16118
rect 18604 15632 18656 15638
rect 18604 15574 18656 15580
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 18420 15088 18472 15094
rect 18616 15042 18644 15574
rect 18420 15030 18472 15036
rect 18432 14890 18460 15030
rect 18524 15026 18644 15042
rect 18512 15020 18644 15026
rect 18564 15014 18644 15020
rect 18512 14962 18564 14968
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17604 14074 17632 14282
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17696 13326 17724 14350
rect 18432 13802 18460 14826
rect 18616 14618 18644 14894
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 16132 12406 16344 12434
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15120 3602 15148 3878
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15672 3126 15700 4490
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15764 2854 15792 4014
rect 15856 3058 15884 4422
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 3602 15976 3878
rect 16316 3670 16344 12406
rect 17236 12238 17264 13126
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16684 3058 16712 4422
rect 17236 4078 17264 12174
rect 18524 8294 18552 13806
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 3618 17356 4014
rect 17512 3738 17540 4082
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 16960 3590 17356 3618
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 3194 16804 3470
rect 16960 3466 16988 3590
rect 17972 3534 18000 3878
rect 17960 3528 18012 3534
rect 17498 3496 17554 3505
rect 16948 3460 17000 3466
rect 17960 3470 18012 3476
rect 17498 3431 17554 3440
rect 16948 3402 17000 3408
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 800 15516 2314
rect 16132 800 16160 2382
rect 17512 1714 17540 3431
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17604 3126 17632 3334
rect 18248 3194 18276 4082
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 18340 2990 18368 3674
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 17420 1686 17540 1714
rect 17420 800 17448 1686
rect 18708 800 18736 22510
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19064 21956 19116 21962
rect 19064 21898 19116 21904
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18984 19514 19012 20470
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 19076 19310 19104 21898
rect 19352 21690 19380 22374
rect 19444 22030 19472 23072
rect 20076 23054 20128 23060
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19890 22128 19946 22137
rect 19890 22063 19892 22072
rect 19944 22063 19946 22072
rect 19892 22034 19944 22040
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19996 21690 20024 22510
rect 20088 22166 20116 23054
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20088 21554 20116 21966
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19352 20942 19380 21082
rect 19444 20942 19472 21490
rect 20074 21448 20130 21457
rect 20074 21383 20130 21392
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19168 19378 19196 20538
rect 19260 20210 19288 20810
rect 19352 20330 19380 20878
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19260 20182 19380 20210
rect 19352 19446 19380 20182
rect 19444 19922 19472 20742
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19904 19922 19932 20198
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19430 19816 19486 19825
rect 19996 19786 20024 19858
rect 19430 19751 19486 19760
rect 19984 19780 20036 19786
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19444 18850 19472 19751
rect 19984 19722 20036 19728
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19260 18822 19472 18850
rect 19260 18170 19288 18822
rect 19536 18766 19564 19246
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19352 18290 19380 18634
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19444 18358 19472 18566
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19338 18184 19394 18193
rect 19260 18142 19338 18170
rect 19338 18119 19394 18128
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17678 19288 18022
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19076 16114 19104 17478
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18892 15094 18920 16050
rect 18880 15088 18932 15094
rect 18880 15030 18932 15036
rect 19076 14822 19104 16050
rect 19168 15978 19196 17070
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 13938 19104 14758
rect 19260 14482 19288 16118
rect 19996 16046 20024 18566
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19352 15570 19380 15846
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19444 15450 19472 15846
rect 19996 15502 20024 15982
rect 19352 15434 19472 15450
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19340 15428 19472 15434
rect 19392 15422 19472 15428
rect 19340 15370 19392 15376
rect 19352 14822 19380 15370
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15094 19472 15302
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19996 14550 20024 15438
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19982 14376 20038 14385
rect 19982 14311 20038 14320
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19628 13530 19656 13806
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19260 3534 19288 3878
rect 19352 3738 19380 7890
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 3058 18828 3334
rect 19352 3194 19380 3470
rect 19444 3194 19472 4082
rect 19996 3602 20024 14311
rect 20088 4758 20116 21383
rect 20180 7954 20208 38218
rect 20260 37256 20312 37262
rect 20260 37198 20312 37204
rect 20272 34746 20300 37198
rect 20352 35080 20404 35086
rect 20352 35022 20404 35028
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 20260 34400 20312 34406
rect 20260 34342 20312 34348
rect 20272 34202 20300 34342
rect 20260 34196 20312 34202
rect 20260 34138 20312 34144
rect 20260 32768 20312 32774
rect 20260 32710 20312 32716
rect 20272 32502 20300 32710
rect 20260 32496 20312 32502
rect 20260 32438 20312 32444
rect 20260 31272 20312 31278
rect 20260 31214 20312 31220
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20180 4078 20208 7754
rect 20272 7562 20300 31214
rect 20364 29306 20392 35022
rect 20352 29300 20404 29306
rect 20352 29242 20404 29248
rect 20364 28422 20392 29242
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 20364 26518 20392 28358
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20364 26314 20392 26454
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20364 7698 20392 25842
rect 20456 7818 20484 38966
rect 22100 38888 22152 38894
rect 22100 38830 22152 38836
rect 20536 38752 20588 38758
rect 20536 38694 20588 38700
rect 20548 35894 20576 38694
rect 22112 38418 22140 38830
rect 22100 38412 22152 38418
rect 22100 38354 22152 38360
rect 21364 38276 21416 38282
rect 21364 38218 21416 38224
rect 21376 37670 21404 38218
rect 21364 37664 21416 37670
rect 21364 37606 21416 37612
rect 21180 36576 21232 36582
rect 21180 36518 21232 36524
rect 21192 36106 21220 36518
rect 21180 36100 21232 36106
rect 21180 36042 21232 36048
rect 21376 35894 21404 37606
rect 21916 37120 21968 37126
rect 21916 37062 21968 37068
rect 21928 36106 21956 37062
rect 22112 36258 22140 38354
rect 22112 36242 22232 36258
rect 22112 36236 22244 36242
rect 22112 36230 22192 36236
rect 22192 36178 22244 36184
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 20548 35866 20668 35894
rect 21376 35866 21496 35894
rect 20536 34740 20588 34746
rect 20536 34682 20588 34688
rect 20548 33998 20576 34682
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20548 33522 20576 33934
rect 20536 33516 20588 33522
rect 20536 33458 20588 33464
rect 20548 32570 20576 33458
rect 20536 32564 20588 32570
rect 20536 32506 20588 32512
rect 20536 32360 20588 32366
rect 20536 32302 20588 32308
rect 20548 30938 20576 32302
rect 20536 30932 20588 30938
rect 20536 30874 20588 30880
rect 20640 30258 20668 35866
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21100 33998 21128 34478
rect 20996 33992 21048 33998
rect 20996 33934 21048 33940
rect 21088 33992 21140 33998
rect 21088 33934 21140 33940
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20824 30258 20852 30534
rect 20916 30394 20944 30534
rect 20904 30388 20956 30394
rect 20904 30330 20956 30336
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 21008 30190 21036 33934
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 21284 32366 21312 32710
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21088 32224 21140 32230
rect 21088 32166 21140 32172
rect 21100 31822 21128 32166
rect 21284 31890 21312 32302
rect 21272 31884 21324 31890
rect 21272 31826 21324 31832
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21088 30796 21140 30802
rect 21088 30738 21140 30744
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20812 29096 20864 29102
rect 20812 29038 20864 29044
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20732 28762 20760 28902
rect 20720 28756 20772 28762
rect 20720 28698 20772 28704
rect 20824 28694 20852 29038
rect 20812 28688 20864 28694
rect 20812 28630 20864 28636
rect 20916 28014 20944 29106
rect 20904 28008 20956 28014
rect 20904 27950 20956 27956
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20732 26994 20760 27814
rect 21008 27470 21036 29242
rect 21100 29170 21128 30738
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 21192 30258 21220 30670
rect 21180 30252 21232 30258
rect 21180 30194 21232 30200
rect 21192 29510 21220 30194
rect 21272 30048 21324 30054
rect 21272 29990 21324 29996
rect 21284 29714 21312 29990
rect 21272 29708 21324 29714
rect 21272 29650 21324 29656
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 21192 29102 21220 29446
rect 21180 29096 21232 29102
rect 21180 29038 21232 29044
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20996 27464 21048 27470
rect 20996 27406 21048 27412
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20824 26042 20852 27406
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 20904 26444 20956 26450
rect 20904 26386 20956 26392
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20628 25968 20680 25974
rect 20628 25910 20680 25916
rect 20536 24336 20588 24342
rect 20536 24278 20588 24284
rect 20548 23254 20576 24278
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 20640 22234 20668 25910
rect 20916 25906 20944 26386
rect 20996 26308 21048 26314
rect 20996 26250 21048 26256
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20732 24750 20760 25842
rect 21008 24750 21036 26250
rect 21100 25226 21128 27338
rect 21192 26858 21220 29038
rect 21272 28688 21324 28694
rect 21272 28630 21324 28636
rect 21284 27334 21312 28630
rect 21364 28620 21416 28626
rect 21364 28562 21416 28568
rect 21376 27606 21404 28562
rect 21364 27600 21416 27606
rect 21364 27542 21416 27548
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 21284 27062 21312 27270
rect 21272 27056 21324 27062
rect 21272 26998 21324 27004
rect 21180 26852 21232 26858
rect 21180 26794 21232 26800
rect 21364 26852 21416 26858
rect 21364 26794 21416 26800
rect 21180 26512 21232 26518
rect 21180 26454 21232 26460
rect 21192 25906 21220 26454
rect 21376 26450 21404 26794
rect 21364 26444 21416 26450
rect 21364 26386 21416 26392
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21284 25770 21312 26250
rect 21272 25764 21324 25770
rect 21272 25706 21324 25712
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 21088 25220 21140 25226
rect 21088 25162 21140 25168
rect 21284 24954 21312 25230
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 20810 23760 20866 23769
rect 20810 23695 20866 23704
rect 20824 23662 20852 23695
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20640 22030 20668 22170
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20548 21706 20576 21830
rect 20548 21678 20668 21706
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20548 20398 20576 21422
rect 20640 21418 20668 21678
rect 20628 21412 20680 21418
rect 20628 21354 20680 21360
rect 20640 21146 20668 21354
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20732 21026 20760 22986
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21284 22234 21312 22510
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 20996 22024 21048 22030
rect 20902 21992 20958 22001
rect 20996 21966 21048 21972
rect 20902 21927 20904 21936
rect 20956 21927 20958 21936
rect 20904 21898 20956 21904
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20824 21554 20852 21830
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20640 20998 20760 21026
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20640 20244 20668 20998
rect 20718 20904 20774 20913
rect 20718 20839 20720 20848
rect 20772 20839 20774 20848
rect 20720 20810 20772 20816
rect 20824 20466 20852 21490
rect 21008 21486 21036 21966
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21008 21146 21036 21422
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 20996 20868 21048 20874
rect 21100 20856 21128 22034
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21192 21622 21220 21898
rect 21284 21690 21312 22170
rect 21376 22166 21404 23054
rect 21364 22160 21416 22166
rect 21364 22102 21416 22108
rect 21468 22094 21496 35866
rect 21548 35760 21600 35766
rect 21548 35702 21600 35708
rect 21560 28150 21588 35702
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21640 35556 21692 35562
rect 21640 35498 21692 35504
rect 21652 35290 21680 35498
rect 21836 35290 21864 35634
rect 21640 35284 21692 35290
rect 21640 35226 21692 35232
rect 21824 35284 21876 35290
rect 21824 35226 21876 35232
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 22112 34202 22140 35022
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22204 34066 22232 36178
rect 22296 35698 22324 47126
rect 25148 45830 25176 49200
rect 25792 46442 25820 49200
rect 25780 46436 25832 46442
rect 25780 46378 25832 46384
rect 25228 46368 25280 46374
rect 25228 46310 25280 46316
rect 25240 45966 25268 46310
rect 26240 46028 26292 46034
rect 26240 45970 26292 45976
rect 25228 45960 25280 45966
rect 25228 45902 25280 45908
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25504 45892 25556 45898
rect 25504 45834 25556 45840
rect 25136 45824 25188 45830
rect 25136 45766 25188 45772
rect 25424 45626 25452 45834
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 22652 39500 22704 39506
rect 22652 39442 22704 39448
rect 22468 39432 22520 39438
rect 22468 39374 22520 39380
rect 22376 38888 22428 38894
rect 22376 38830 22428 38836
rect 22388 38554 22416 38830
rect 22376 38548 22428 38554
rect 22376 38490 22428 38496
rect 22376 36576 22428 36582
rect 22376 36518 22428 36524
rect 22388 35698 22416 36518
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22480 35578 22508 39374
rect 22664 39030 22692 39442
rect 25516 39438 25544 45834
rect 26252 45830 26280 45970
rect 26240 45824 26292 45830
rect 26240 45766 26292 45772
rect 26712 45554 26740 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 28368 46986 28396 49200
rect 29656 47054 29684 49200
rect 30196 47184 30248 47190
rect 30196 47126 30248 47132
rect 28448 47048 28500 47054
rect 28448 46990 28500 46996
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 28356 46980 28408 46986
rect 28356 46922 28408 46928
rect 27620 46504 27672 46510
rect 27620 46446 27672 46452
rect 27632 46170 27660 46446
rect 27620 46164 27672 46170
rect 27620 46106 27672 46112
rect 26528 45526 26740 45554
rect 26056 45484 26108 45490
rect 26056 45426 26108 45432
rect 25504 39432 25556 39438
rect 25504 39374 25556 39380
rect 23480 39296 23532 39302
rect 23480 39238 23532 39244
rect 25320 39296 25372 39302
rect 25320 39238 25372 39244
rect 22652 39024 22704 39030
rect 22836 39024 22888 39030
rect 22704 38984 22784 39012
rect 22652 38966 22704 38972
rect 22388 35550 22508 35578
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22192 34060 22244 34066
rect 22192 34002 22244 34008
rect 22008 33992 22060 33998
rect 22060 33952 22140 33980
rect 22008 33934 22060 33940
rect 22008 33516 22060 33522
rect 22008 33458 22060 33464
rect 21824 33312 21876 33318
rect 21824 33254 21876 33260
rect 21836 32978 21864 33254
rect 22020 33114 22048 33458
rect 22008 33108 22060 33114
rect 22008 33050 22060 33056
rect 21824 32972 21876 32978
rect 21824 32914 21876 32920
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 21928 32026 21956 32370
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 21928 31346 21956 31962
rect 22112 31754 22140 33952
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 22204 33114 22232 33254
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 21916 31340 21968 31346
rect 21916 31282 21968 31288
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21836 30734 21864 31078
rect 21928 30734 21956 31282
rect 22112 31278 22140 31690
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 22008 30660 22060 30666
rect 22008 30602 22060 30608
rect 21914 29608 21970 29617
rect 22020 29594 22048 30602
rect 21970 29566 22048 29594
rect 21914 29543 21970 29552
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 21744 28762 21772 29106
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21732 28552 21784 28558
rect 21732 28494 21784 28500
rect 21548 28144 21600 28150
rect 21548 28086 21600 28092
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21560 26518 21588 26726
rect 21744 26518 21772 28494
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 21836 28082 21864 28358
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21928 27470 21956 29543
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 21928 27282 21956 27406
rect 22020 27402 22048 28018
rect 22008 27396 22060 27402
rect 22008 27338 22060 27344
rect 21928 27254 22048 27282
rect 21916 27056 21968 27062
rect 21916 26998 21968 27004
rect 21548 26512 21600 26518
rect 21548 26454 21600 26460
rect 21732 26512 21784 26518
rect 21732 26454 21784 26460
rect 21560 26382 21588 26454
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21560 25838 21588 26318
rect 21744 26314 21772 26454
rect 21732 26308 21784 26314
rect 21732 26250 21784 26256
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 21548 25832 21600 25838
rect 21548 25774 21600 25780
rect 21548 25424 21600 25430
rect 21548 25366 21600 25372
rect 21560 25294 21588 25366
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21560 24818 21588 25230
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21836 24426 21864 26250
rect 21928 25430 21956 26998
rect 21916 25424 21968 25430
rect 21916 25366 21968 25372
rect 21928 24614 21956 25366
rect 22020 25294 22048 27254
rect 22112 26926 22140 28426
rect 22192 28008 22244 28014
rect 22192 27950 22244 27956
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22112 24750 22140 25094
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21836 24398 21956 24426
rect 21824 23316 21876 23322
rect 21928 23304 21956 24398
rect 22008 23316 22060 23322
rect 21928 23276 22008 23304
rect 21824 23258 21876 23264
rect 22008 23258 22060 23264
rect 21836 22642 21864 23258
rect 22020 22778 22048 23258
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21730 22128 21786 22137
rect 21468 22066 21680 22094
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 21284 20913 21312 21626
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21468 21010 21496 21286
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21364 20936 21416 20942
rect 21048 20828 21128 20856
rect 21270 20904 21326 20913
rect 21364 20878 21416 20884
rect 21270 20839 21326 20848
rect 20996 20810 21048 20816
rect 21100 20754 21128 20828
rect 21376 20754 21404 20878
rect 21100 20726 21404 20754
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20548 20216 20668 20244
rect 20548 17762 20576 20216
rect 20824 20074 20852 20402
rect 20640 20046 20852 20074
rect 20640 19718 20668 20046
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 18222 20668 19654
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20548 17734 20668 17762
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20548 17270 20576 17546
rect 20640 17354 20668 17734
rect 20640 17326 20760 17354
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20640 16114 20668 17138
rect 20732 16182 20760 17326
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20640 15026 20668 15846
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20824 14906 20852 18702
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 20640 14878 20852 14906
rect 20640 14074 20668 14878
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20364 7670 20576 7698
rect 20272 7534 20392 7562
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19996 3058 20024 3334
rect 20088 3058 20116 3878
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20180 3194 20208 3470
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19352 800 19380 2926
rect 20272 2446 20300 3334
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 870 20208 898
rect 19996 800 20024 870
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20180 762 20208 870
rect 20364 762 20392 7534
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20456 2650 20484 4082
rect 20548 2650 20576 7670
rect 20640 4078 20668 14010
rect 20732 8090 20760 14418
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20916 4282 20944 4558
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 3058 20760 3878
rect 20824 3194 20852 4082
rect 21192 3670 21220 4082
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20916 2854 20944 3130
rect 21284 2990 21312 18158
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21560 16998 21588 17546
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21560 15570 21588 16390
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21652 14278 21680 22066
rect 21730 22063 21786 22072
rect 21744 21690 21772 22063
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21836 20602 21864 22578
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 22020 20534 22048 21286
rect 22112 21010 22140 21966
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21928 19786 21956 20198
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 21916 19780 21968 19786
rect 21916 19722 21968 19728
rect 22020 19446 22048 19790
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21836 18290 21864 18702
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21836 17678 21864 18226
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21916 17604 21968 17610
rect 21916 17546 21968 17552
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21836 17270 21864 17478
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21836 16726 21864 17206
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21928 16250 21956 17546
rect 22112 17066 22140 18158
rect 22100 17060 22152 17066
rect 22100 17002 22152 17008
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16590 22048 16934
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22020 15026 22048 16050
rect 22112 15978 22140 16594
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 13938 21680 14214
rect 22112 14074 22140 14282
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21376 3670 21404 13806
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 22020 12442 22048 12718
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21732 4004 21784 4010
rect 21732 3946 21784 3952
rect 21916 4004 21968 4010
rect 21916 3946 21968 3952
rect 21744 3738 21772 3946
rect 21732 3732 21784 3738
rect 21732 3674 21784 3680
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21928 3058 21956 3946
rect 22204 3942 22232 27950
rect 22296 22094 22324 32914
rect 22388 26874 22416 35550
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22480 27010 22508 34886
rect 22572 34542 22600 35226
rect 22664 35086 22692 35566
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22560 34536 22612 34542
rect 22560 34478 22612 34484
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22572 33998 22600 34342
rect 22756 33998 22784 38984
rect 22836 38966 22888 38972
rect 22848 38010 22876 38966
rect 23492 38350 23520 39238
rect 25332 39098 25360 39238
rect 25320 39092 25372 39098
rect 25320 39034 25372 39040
rect 25504 38956 25556 38962
rect 25504 38898 25556 38904
rect 24400 38888 24452 38894
rect 24400 38830 24452 38836
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23664 38208 23716 38214
rect 23664 38150 23716 38156
rect 22836 38004 22888 38010
rect 22836 37946 22888 37952
rect 23676 37942 23704 38150
rect 23664 37936 23716 37942
rect 23664 37878 23716 37884
rect 24412 37874 24440 38830
rect 24584 38276 24636 38282
rect 24584 38218 24636 38224
rect 25412 38276 25464 38282
rect 25412 38218 25464 38224
rect 24492 38208 24544 38214
rect 24492 38150 24544 38156
rect 24400 37868 24452 37874
rect 24400 37810 24452 37816
rect 24412 37398 24440 37810
rect 24504 37806 24532 38150
rect 24596 38010 24624 38218
rect 25424 38010 25452 38218
rect 24584 38004 24636 38010
rect 24584 37946 24636 37952
rect 25412 38004 25464 38010
rect 25412 37946 25464 37952
rect 24860 37868 24912 37874
rect 24860 37810 24912 37816
rect 24492 37800 24544 37806
rect 24492 37742 24544 37748
rect 24400 37392 24452 37398
rect 24400 37334 24452 37340
rect 23388 36236 23440 36242
rect 23388 36178 23440 36184
rect 22928 36100 22980 36106
rect 22928 36042 22980 36048
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22560 33992 22612 33998
rect 22560 33934 22612 33940
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 22560 33312 22612 33318
rect 22560 33254 22612 33260
rect 22572 32910 22600 33254
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22848 28082 22876 35634
rect 22940 34610 22968 36042
rect 23400 35290 23428 36178
rect 23572 36032 23624 36038
rect 23572 35974 23624 35980
rect 23584 35698 23612 35974
rect 23572 35692 23624 35698
rect 23572 35634 23624 35640
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23480 35148 23532 35154
rect 23480 35090 23532 35096
rect 22928 34604 22980 34610
rect 22928 34546 22980 34552
rect 23204 34400 23256 34406
rect 23204 34342 23256 34348
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 22928 32904 22980 32910
rect 22928 32846 22980 32852
rect 22940 32570 22968 32846
rect 22928 32564 22980 32570
rect 22928 32506 22980 32512
rect 23032 28558 23060 33934
rect 23216 32366 23244 34342
rect 23296 34060 23348 34066
rect 23296 34002 23348 34008
rect 23308 33658 23336 34002
rect 23296 33652 23348 33658
rect 23296 33594 23348 33600
rect 23492 32570 23520 35090
rect 23584 35018 23612 35634
rect 23572 35012 23624 35018
rect 23572 34954 23624 34960
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23204 32360 23256 32366
rect 23204 32302 23256 32308
rect 23400 31822 23428 32370
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23296 31748 23348 31754
rect 23296 31690 23348 31696
rect 23204 31680 23256 31686
rect 23204 31622 23256 31628
rect 23112 31340 23164 31346
rect 23112 31282 23164 31288
rect 23124 28762 23152 31282
rect 23216 30734 23244 31622
rect 23308 31210 23336 31690
rect 23296 31204 23348 31210
rect 23296 31146 23348 31152
rect 23480 31136 23532 31142
rect 23480 31078 23532 31084
rect 23492 30802 23520 31078
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23216 29753 23244 30126
rect 23202 29744 23258 29753
rect 23202 29679 23258 29688
rect 23216 29646 23244 29679
rect 23204 29640 23256 29646
rect 23388 29640 23440 29646
rect 23204 29582 23256 29588
rect 23308 29600 23388 29628
rect 23112 28756 23164 28762
rect 23112 28698 23164 28704
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 23032 27606 23060 28494
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 22480 26994 22600 27010
rect 22468 26988 22600 26994
rect 22520 26982 22600 26988
rect 22468 26930 22520 26936
rect 22388 26846 22508 26874
rect 22296 22066 22416 22094
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22296 21146 22324 21422
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22296 19514 22324 19722
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22388 18902 22416 22066
rect 22480 22001 22508 26846
rect 22572 26450 22600 26982
rect 22560 26444 22612 26450
rect 22560 26386 22612 26392
rect 22848 25430 22876 27406
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 25498 23060 26182
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 22836 25424 22888 25430
rect 22836 25366 22888 25372
rect 23124 25294 23152 28698
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23204 24812 23256 24818
rect 23204 24754 23256 24760
rect 23216 24410 23244 24754
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23204 24404 23256 24410
rect 23204 24346 23256 24352
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22572 23050 22600 23258
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22466 21992 22522 22001
rect 22466 21927 22522 21936
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22572 21622 22600 21830
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 22376 18896 22428 18902
rect 22376 18838 22428 18844
rect 22664 18086 22692 23258
rect 22848 23118 22876 24142
rect 23124 23730 23152 24346
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 23308 23633 23336 29600
rect 23584 29628 23612 33798
rect 23664 33448 23716 33454
rect 23664 33390 23716 33396
rect 23676 32842 23704 33390
rect 23664 32836 23716 32842
rect 23664 32778 23716 32784
rect 23676 30326 23704 32778
rect 23860 30920 23888 34138
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 23940 33448 23992 33454
rect 23940 33390 23992 33396
rect 23952 32910 23980 33390
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 23952 31958 23980 32846
rect 24136 32434 24164 33458
rect 24504 33386 24532 37742
rect 24872 37126 24900 37810
rect 24952 37732 25004 37738
rect 24952 37674 25004 37680
rect 24860 37120 24912 37126
rect 24860 37062 24912 37068
rect 24964 36922 24992 37674
rect 25516 37262 25544 38898
rect 25964 38344 26016 38350
rect 25964 38286 26016 38292
rect 25976 37874 26004 38286
rect 25964 37868 26016 37874
rect 25964 37810 26016 37816
rect 25780 37392 25832 37398
rect 25780 37334 25832 37340
rect 25504 37256 25556 37262
rect 25504 37198 25556 37204
rect 25596 37256 25648 37262
rect 25596 37198 25648 37204
rect 25412 37120 25464 37126
rect 25412 37062 25464 37068
rect 24952 36916 25004 36922
rect 24952 36858 25004 36864
rect 25228 36848 25280 36854
rect 25228 36790 25280 36796
rect 24676 36780 24728 36786
rect 24676 36722 24728 36728
rect 24688 36310 24716 36722
rect 24860 36644 24912 36650
rect 24860 36586 24912 36592
rect 24872 36310 24900 36586
rect 24676 36304 24728 36310
rect 24676 36246 24728 36252
rect 24860 36304 24912 36310
rect 24860 36246 24912 36252
rect 25240 36242 25268 36790
rect 25228 36236 25280 36242
rect 25228 36178 25280 36184
rect 25424 36174 25452 37062
rect 25412 36168 25464 36174
rect 25412 36110 25464 36116
rect 25504 36100 25556 36106
rect 25504 36042 25556 36048
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 24676 35488 24728 35494
rect 24676 35430 24728 35436
rect 24584 35284 24636 35290
rect 24584 35226 24636 35232
rect 24596 35057 24624 35226
rect 24688 35193 24716 35430
rect 24780 35290 24808 35566
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 25516 35222 25544 36042
rect 25608 35698 25636 37198
rect 25792 36922 25820 37334
rect 25872 37188 25924 37194
rect 25872 37130 25924 37136
rect 25688 36916 25740 36922
rect 25688 36858 25740 36864
rect 25780 36916 25832 36922
rect 25780 36858 25832 36864
rect 25700 36718 25728 36858
rect 25688 36712 25740 36718
rect 25688 36654 25740 36660
rect 25700 36258 25728 36654
rect 25700 36230 25820 36258
rect 25688 36100 25740 36106
rect 25688 36042 25740 36048
rect 25596 35692 25648 35698
rect 25596 35634 25648 35640
rect 25700 35630 25728 36042
rect 25688 35624 25740 35630
rect 25688 35566 25740 35572
rect 25792 35494 25820 36230
rect 25884 36038 25912 37130
rect 25964 36712 26016 36718
rect 25964 36654 26016 36660
rect 25976 36310 26004 36654
rect 25964 36304 26016 36310
rect 25964 36246 26016 36252
rect 25872 36032 25924 36038
rect 25872 35974 25924 35980
rect 25884 35562 25912 35974
rect 25872 35556 25924 35562
rect 25872 35498 25924 35504
rect 25780 35488 25832 35494
rect 25780 35430 25832 35436
rect 25504 35216 25556 35222
rect 24674 35184 24730 35193
rect 25504 35158 25556 35164
rect 24674 35119 24730 35128
rect 24582 35048 24638 35057
rect 24582 34983 24584 34992
rect 24636 34983 24638 34992
rect 24584 34954 24636 34960
rect 24584 34604 24636 34610
rect 24584 34546 24636 34552
rect 24400 33380 24452 33386
rect 24400 33322 24452 33328
rect 24492 33380 24544 33386
rect 24492 33322 24544 33328
rect 24412 33114 24440 33322
rect 24400 33108 24452 33114
rect 24400 33050 24452 33056
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 23940 31952 23992 31958
rect 23940 31894 23992 31900
rect 23952 31346 23980 31894
rect 24136 31822 24164 32370
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 24412 31890 24440 32166
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 24124 31816 24176 31822
rect 24124 31758 24176 31764
rect 24136 31346 24164 31758
rect 24596 31482 24624 34546
rect 25136 34536 25188 34542
rect 25136 34478 25188 34484
rect 25148 33930 25176 34478
rect 25228 34196 25280 34202
rect 25228 34138 25280 34144
rect 24676 33924 24728 33930
rect 24676 33866 24728 33872
rect 25136 33924 25188 33930
rect 25136 33866 25188 33872
rect 24688 32978 24716 33866
rect 25044 33584 25096 33590
rect 25044 33526 25096 33532
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24964 32978 24992 33254
rect 24676 32972 24728 32978
rect 24676 32914 24728 32920
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 25056 32570 25084 33526
rect 25240 33522 25268 34138
rect 25320 33856 25372 33862
rect 25320 33798 25372 33804
rect 25332 33522 25360 33798
rect 25228 33516 25280 33522
rect 25228 33458 25280 33464
rect 25320 33516 25372 33522
rect 25320 33458 25372 33464
rect 25240 33046 25268 33458
rect 25228 33040 25280 33046
rect 25228 32982 25280 32988
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24768 32020 24820 32026
rect 24768 31962 24820 31968
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 23940 31340 23992 31346
rect 23940 31282 23992 31288
rect 24124 31340 24176 31346
rect 24124 31282 24176 31288
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 23940 30932 23992 30938
rect 23860 30892 23940 30920
rect 23940 30874 23992 30880
rect 23848 30728 23900 30734
rect 23848 30670 23900 30676
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 23768 29714 23796 30534
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23664 29640 23716 29646
rect 23584 29600 23664 29628
rect 23388 29582 23440 29588
rect 23664 29582 23716 29588
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23584 29238 23612 29446
rect 23572 29232 23624 29238
rect 23572 29174 23624 29180
rect 23676 29102 23704 29582
rect 23860 29510 23888 30670
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23952 28490 23980 30874
rect 24596 30297 24624 31282
rect 24780 30802 24808 31962
rect 24872 31890 24900 32370
rect 24860 31884 24912 31890
rect 24860 31826 24912 31832
rect 24872 31414 24900 31826
rect 24860 31408 24912 31414
rect 24860 31350 24912 31356
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 24582 30288 24638 30297
rect 24582 30223 24638 30232
rect 24216 30048 24268 30054
rect 24216 29990 24268 29996
rect 24492 30048 24544 30054
rect 24492 29990 24544 29996
rect 24228 28966 24256 29990
rect 24504 29646 24532 29990
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24216 28960 24268 28966
rect 24216 28902 24268 28908
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23400 28082 23428 28358
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23400 27470 23428 28018
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23664 27396 23716 27402
rect 23664 27338 23716 27344
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23388 27056 23440 27062
rect 23388 26998 23440 27004
rect 23400 26450 23428 26998
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23584 25838 23612 27270
rect 23676 26926 23704 27338
rect 24124 26988 24176 26994
rect 24124 26930 24176 26936
rect 23664 26920 23716 26926
rect 23664 26862 23716 26868
rect 23676 26314 23704 26862
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23664 26308 23716 26314
rect 23664 26250 23716 26256
rect 23676 25838 23704 26250
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23860 25786 23888 26726
rect 24136 26518 24164 26930
rect 24400 26852 24452 26858
rect 24400 26794 24452 26800
rect 24124 26512 24176 26518
rect 24124 26454 24176 26460
rect 24412 26382 24440 26794
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24492 25968 24544 25974
rect 24492 25910 24544 25916
rect 23860 25770 24072 25786
rect 23860 25764 24084 25770
rect 23860 25758 24032 25764
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23492 24954 23520 25638
rect 23860 25294 23888 25758
rect 24032 25706 24084 25712
rect 24504 25498 24532 25910
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 23848 25288 23900 25294
rect 23848 25230 23900 25236
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 24412 24206 24440 25230
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24412 23866 24440 24142
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 23294 23624 23350 23633
rect 23294 23559 23350 23568
rect 23492 23118 23520 23802
rect 24412 23730 24440 23802
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24596 23526 24624 30223
rect 24872 29730 24900 31350
rect 25056 30954 25084 32506
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25240 32026 25268 32302
rect 25228 32020 25280 32026
rect 25228 31962 25280 31968
rect 25134 31648 25190 31657
rect 25134 31583 25190 31592
rect 24964 30926 25084 30954
rect 24964 30326 24992 30926
rect 25148 30326 25176 31583
rect 25320 30932 25372 30938
rect 25320 30874 25372 30880
rect 25228 30592 25280 30598
rect 25228 30534 25280 30540
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 25136 30320 25188 30326
rect 25136 30262 25188 30268
rect 25240 30258 25268 30534
rect 25332 30258 25360 30874
rect 26068 30818 26096 45426
rect 26424 43784 26476 43790
rect 26424 43726 26476 43732
rect 26148 38208 26200 38214
rect 26148 38150 26200 38156
rect 26160 37466 26188 38150
rect 26148 37460 26200 37466
rect 26148 37402 26200 37408
rect 26160 36786 26188 37402
rect 26240 36848 26292 36854
rect 26240 36790 26292 36796
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 26252 36174 26280 36790
rect 26436 36378 26464 43726
rect 26528 41414 26556 45526
rect 26528 41386 26740 41414
rect 26424 36372 26476 36378
rect 26424 36314 26476 36320
rect 26240 36168 26292 36174
rect 26240 36110 26292 36116
rect 26148 31408 26200 31414
rect 26148 31350 26200 31356
rect 26160 30938 26188 31350
rect 26252 31142 26280 36110
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26344 34678 26372 35022
rect 26332 34672 26384 34678
rect 26332 34614 26384 34620
rect 26332 32224 26384 32230
rect 26332 32166 26384 32172
rect 26344 31890 26372 32166
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 26240 31136 26292 31142
rect 26240 31078 26292 31084
rect 26148 30932 26200 30938
rect 26148 30874 26200 30880
rect 26068 30790 26188 30818
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 25596 30660 25648 30666
rect 25596 30602 25648 30608
rect 25228 30252 25280 30258
rect 25228 30194 25280 30200
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 24780 29714 24900 29730
rect 24768 29708 24900 29714
rect 24820 29702 24900 29708
rect 24768 29650 24820 29656
rect 24766 29608 24822 29617
rect 24766 29543 24768 29552
rect 24820 29543 24822 29552
rect 24768 29514 24820 29520
rect 24872 29306 24900 29702
rect 25608 29646 25636 30602
rect 26068 29714 26096 30670
rect 26056 29708 26108 29714
rect 26056 29650 26108 29656
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24676 28960 24728 28966
rect 24676 28902 24728 28908
rect 24688 28558 24716 28902
rect 24964 28626 24992 29446
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24688 24954 24716 28494
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 25362 24900 25638
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24676 24948 24728 24954
rect 24676 24890 24728 24896
rect 25044 24948 25096 24954
rect 25044 24890 25096 24896
rect 24688 24750 24716 24890
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24688 24274 24716 24686
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 22940 22710 22968 22918
rect 22928 22704 22980 22710
rect 22928 22646 22980 22652
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 23124 20602 23152 22442
rect 23308 21962 23336 22510
rect 23296 21956 23348 21962
rect 23296 21898 23348 21904
rect 23308 21486 23336 21898
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23124 18834 23152 20538
rect 23216 20466 23244 20878
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23308 20466 23336 20742
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23216 20346 23244 20402
rect 23216 20318 23336 20346
rect 23308 19990 23336 20318
rect 23296 19984 23348 19990
rect 23296 19926 23348 19932
rect 23400 19854 23428 22918
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23676 21554 23704 21830
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24136 20534 24164 21422
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 24596 19786 24624 23462
rect 24584 19780 24636 19786
rect 24584 19722 24636 19728
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 23308 18630 23336 19314
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22664 17202 22692 18022
rect 23308 17882 23336 18566
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23204 17672 23256 17678
rect 23308 17660 23336 17818
rect 23256 17632 23336 17660
rect 23204 17614 23256 17620
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23216 17202 23244 17478
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22296 16232 22324 16730
rect 23308 16658 23336 17632
rect 23400 17542 23428 18158
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23492 17270 23520 18022
rect 23676 17678 23704 18770
rect 23940 18352 23992 18358
rect 23940 18294 23992 18300
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23860 17746 23888 18226
rect 23952 18222 23980 18294
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23296 16652 23348 16658
rect 23296 16594 23348 16600
rect 23676 16522 23704 17614
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 23664 16516 23716 16522
rect 23664 16458 23716 16464
rect 22388 16402 22416 16458
rect 22388 16374 22508 16402
rect 22376 16244 22428 16250
rect 22296 16204 22376 16232
rect 22376 16186 22428 16192
rect 22284 15428 22336 15434
rect 22284 15370 22336 15376
rect 22296 15162 22324 15370
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22388 12918 22416 16186
rect 22480 16182 22508 16374
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22480 15366 22508 16118
rect 23768 16046 23796 17546
rect 23952 17542 23980 18158
rect 24032 17808 24084 17814
rect 24032 17750 24084 17756
rect 24044 17626 24072 17750
rect 24228 17626 24256 18226
rect 24504 18222 24532 18770
rect 24596 18766 24624 19722
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24780 18290 24808 18566
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24492 18216 24544 18222
rect 24492 18158 24544 18164
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24688 17814 24716 18022
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 24044 17598 24256 17626
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 24044 17134 24072 17598
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 24780 16538 24808 18226
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24872 17270 24900 18022
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24688 16510 24808 16538
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23860 16114 23888 16390
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24596 15706 24624 15982
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24688 15502 24716 16510
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24780 15706 24808 16118
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 14482 22508 15302
rect 24688 15026 24716 15438
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 23400 6866 23428 14418
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 24860 4480 24912 4486
rect 24860 4422 24912 4428
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22112 2990 22140 3878
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 22204 2650 22232 3470
rect 22296 3466 22324 4082
rect 23400 3534 23428 4422
rect 24872 3738 24900 4422
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 23664 3596 23716 3602
rect 23664 3538 23716 3544
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 20640 800 20668 2314
rect 21928 800 21956 2314
rect 22572 800 22600 2926
rect 23676 2650 23704 3538
rect 24584 3460 24636 3466
rect 24584 3402 24636 3408
rect 24596 3058 24624 3402
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24780 2990 24808 3334
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 25056 2650 25084 24890
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23216 800 23244 2382
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 24504 800 24532 2314
rect 25148 800 25176 2926
rect 25240 2310 25268 29582
rect 25608 29170 25636 29582
rect 25688 29504 25740 29510
rect 25688 29446 25740 29452
rect 25700 29238 25728 29446
rect 25688 29232 25740 29238
rect 25688 29174 25740 29180
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25964 28960 26016 28966
rect 25964 28902 26016 28908
rect 25976 28490 26004 28902
rect 26068 28762 26096 29650
rect 26056 28756 26108 28762
rect 26056 28698 26108 28704
rect 26160 28642 26188 30790
rect 26252 29510 26280 31078
rect 26240 29504 26292 29510
rect 26240 29446 26292 29452
rect 26068 28614 26188 28642
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 25424 24274 25452 25094
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25516 23118 25544 28018
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 25596 26852 25648 26858
rect 25596 26794 25648 26800
rect 25608 25294 25636 26794
rect 25700 26450 25728 26930
rect 25780 26920 25832 26926
rect 25780 26862 25832 26868
rect 25688 26444 25740 26450
rect 25688 26386 25740 26392
rect 25792 25906 25820 26862
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25872 25356 25924 25362
rect 25872 25298 25924 25304
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 25792 24954 25820 25230
rect 25780 24948 25832 24954
rect 25780 24890 25832 24896
rect 25884 23322 25912 25298
rect 26068 24410 26096 28614
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26148 26376 26200 26382
rect 26252 26364 26280 26726
rect 26200 26336 26280 26364
rect 26148 26318 26200 26324
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 26252 25838 26280 26182
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 26252 25430 26280 25774
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26252 24682 26280 25094
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26056 24404 26108 24410
rect 26056 24346 26108 24352
rect 25964 24132 26016 24138
rect 25964 24074 26016 24080
rect 25976 23866 26004 24074
rect 25964 23860 26016 23866
rect 25964 23802 26016 23808
rect 25872 23316 25924 23322
rect 25872 23258 25924 23264
rect 25504 23112 25556 23118
rect 25504 23054 25556 23060
rect 25964 22432 26016 22438
rect 25964 22374 26016 22380
rect 25976 22098 26004 22374
rect 25964 22092 26016 22098
rect 25964 22034 26016 22040
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 25504 21888 25556 21894
rect 25504 21830 25556 21836
rect 25516 21622 25544 21830
rect 25504 21616 25556 21622
rect 25504 21558 25556 21564
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25332 21146 25360 21422
rect 26344 21418 26372 21898
rect 26332 21412 26384 21418
rect 26332 21354 26384 21360
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 26252 20942 26280 21286
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26344 19514 26372 19790
rect 26332 19508 26384 19514
rect 26332 19450 26384 19456
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25608 18834 25636 19246
rect 25596 18828 25648 18834
rect 25596 18770 25648 18776
rect 25504 18352 25556 18358
rect 25504 18294 25556 18300
rect 25516 17678 25544 18294
rect 25608 17882 25636 18770
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25700 18154 25728 18226
rect 25688 18148 25740 18154
rect 25688 18090 25740 18096
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25700 17678 25728 18090
rect 25976 18086 26004 18702
rect 26160 18358 26188 19314
rect 26148 18352 26200 18358
rect 26148 18294 26200 18300
rect 26436 18290 26464 36314
rect 26712 31754 26740 41386
rect 26976 38412 27028 38418
rect 26976 38354 27028 38360
rect 26988 37874 27016 38354
rect 27988 38208 28040 38214
rect 27988 38150 28040 38156
rect 28264 38208 28316 38214
rect 28264 38150 28316 38156
rect 28000 37942 28028 38150
rect 27988 37936 28040 37942
rect 27988 37878 28040 37884
rect 26976 37868 27028 37874
rect 26976 37810 27028 37816
rect 26988 37330 27016 37810
rect 27252 37800 27304 37806
rect 27252 37742 27304 37748
rect 26976 37324 27028 37330
rect 26976 37266 27028 37272
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26804 36378 26832 37198
rect 27264 36922 27292 37742
rect 28276 37670 28304 38150
rect 28264 37664 28316 37670
rect 28264 37606 28316 37612
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 27252 36916 27304 36922
rect 27252 36858 27304 36864
rect 27988 36916 28040 36922
rect 27988 36858 28040 36864
rect 27252 36780 27304 36786
rect 27252 36722 27304 36728
rect 27528 36780 27580 36786
rect 27528 36722 27580 36728
rect 26792 36372 26844 36378
rect 26792 36314 26844 36320
rect 26884 36100 26936 36106
rect 26884 36042 26936 36048
rect 26712 31726 26832 31754
rect 26700 31340 26752 31346
rect 26700 31282 26752 31288
rect 26712 29578 26740 31282
rect 26700 29572 26752 29578
rect 26700 29514 26752 29520
rect 26712 29345 26740 29514
rect 26698 29336 26754 29345
rect 26698 29271 26754 29280
rect 26516 27600 26568 27606
rect 26516 27542 26568 27548
rect 26528 26518 26556 27542
rect 26516 26512 26568 26518
rect 26516 26454 26568 26460
rect 26516 26376 26568 26382
rect 26516 26318 26568 26324
rect 26528 25906 26556 26318
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26528 24954 26556 25842
rect 26608 25288 26660 25294
rect 26608 25230 26660 25236
rect 26516 24948 26568 24954
rect 26516 24890 26568 24896
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26424 18284 26476 18290
rect 26424 18226 26476 18232
rect 25964 18080 26016 18086
rect 25964 18022 26016 18028
rect 26528 17678 26556 19314
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25516 15706 25544 15846
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 26620 5098 26648 25230
rect 26804 23798 26832 31726
rect 26896 30054 26924 36042
rect 26976 35760 27028 35766
rect 26976 35702 27028 35708
rect 26988 34746 27016 35702
rect 27160 35624 27212 35630
rect 27160 35566 27212 35572
rect 27172 35086 27200 35566
rect 27264 35290 27292 36722
rect 27436 36032 27488 36038
rect 27436 35974 27488 35980
rect 27448 35698 27476 35974
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 27448 35136 27476 35634
rect 27356 35108 27476 35136
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 26976 34740 27028 34746
rect 26976 34682 27028 34688
rect 27172 34542 27200 35022
rect 27356 35018 27384 35108
rect 27344 35012 27396 35018
rect 27344 34954 27396 34960
rect 27436 35012 27488 35018
rect 27436 34954 27488 34960
rect 27448 34610 27476 34954
rect 27436 34604 27488 34610
rect 27436 34546 27488 34552
rect 27160 34536 27212 34542
rect 27160 34478 27212 34484
rect 27540 34474 27568 36722
rect 27712 36644 27764 36650
rect 27712 36586 27764 36592
rect 27724 36378 27752 36586
rect 27896 36576 27948 36582
rect 27896 36518 27948 36524
rect 27712 36372 27764 36378
rect 27712 36314 27764 36320
rect 27908 35170 27936 36518
rect 28000 36174 28028 36858
rect 28080 36304 28132 36310
rect 28080 36246 28132 36252
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 28092 35290 28120 36246
rect 28172 35760 28224 35766
rect 28172 35702 28224 35708
rect 28080 35284 28132 35290
rect 28080 35226 28132 35232
rect 28078 35184 28134 35193
rect 27804 35148 27856 35154
rect 27908 35142 28028 35170
rect 27804 35090 27856 35096
rect 27712 34944 27764 34950
rect 27712 34886 27764 34892
rect 27724 34542 27752 34886
rect 27712 34536 27764 34542
rect 27712 34478 27764 34484
rect 27528 34468 27580 34474
rect 27528 34410 27580 34416
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27264 32978 27292 33866
rect 27344 33856 27396 33862
rect 27344 33798 27396 33804
rect 27356 33522 27384 33798
rect 27344 33516 27396 33522
rect 27344 33458 27396 33464
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27160 32768 27212 32774
rect 27160 32710 27212 32716
rect 27172 32434 27200 32710
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 27080 31482 27108 32370
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27068 31476 27120 31482
rect 27068 31418 27120 31424
rect 27172 31346 27200 32166
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27068 31136 27120 31142
rect 27068 31078 27120 31084
rect 27080 30802 27108 31078
rect 27068 30796 27120 30802
rect 27068 30738 27120 30744
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 26884 30048 26936 30054
rect 26884 29990 26936 29996
rect 26896 27130 26924 29990
rect 26976 29504 27028 29510
rect 26976 29446 27028 29452
rect 26988 29209 27016 29446
rect 26974 29200 27030 29209
rect 26974 29135 27030 29144
rect 26988 28762 27016 29135
rect 26976 28756 27028 28762
rect 26976 28698 27028 28704
rect 27080 28558 27108 30194
rect 27264 29510 27292 32914
rect 27436 32768 27488 32774
rect 27436 32710 27488 32716
rect 27344 31884 27396 31890
rect 27344 31826 27396 31832
rect 27356 31686 27384 31826
rect 27344 31680 27396 31686
rect 27344 31622 27396 31628
rect 27344 31340 27396 31346
rect 27344 31282 27396 31288
rect 27252 29504 27304 29510
rect 27252 29446 27304 29452
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 26976 28484 27028 28490
rect 26976 28426 27028 28432
rect 26988 28082 27016 28426
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 26884 27124 26936 27130
rect 26884 27066 26936 27072
rect 27080 26790 27108 28018
rect 27264 27470 27292 29446
rect 27252 27464 27304 27470
rect 27252 27406 27304 27412
rect 27068 26784 27120 26790
rect 27068 26726 27120 26732
rect 27264 26382 27292 27406
rect 27068 26376 27120 26382
rect 27252 26376 27304 26382
rect 27120 26336 27200 26364
rect 27068 26318 27120 26324
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26896 25294 26924 25638
rect 26988 25294 27016 26250
rect 27172 25906 27200 26336
rect 27252 26318 27304 26324
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 26792 23792 26844 23798
rect 26792 23734 26844 23740
rect 26988 23730 27016 24754
rect 27172 24410 27200 25842
rect 27356 24614 27384 31282
rect 27448 30938 27476 32710
rect 27620 32292 27672 32298
rect 27620 32234 27672 32240
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27436 30932 27488 30938
rect 27436 30874 27488 30880
rect 27540 30734 27568 31826
rect 27632 31346 27660 32234
rect 27816 31657 27844 35090
rect 27896 35080 27948 35086
rect 27896 35022 27948 35028
rect 27802 31648 27858 31657
rect 27802 31583 27858 31592
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27528 30728 27580 30734
rect 27528 30670 27580 30676
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 27528 30184 27580 30190
rect 27528 30126 27580 30132
rect 27540 30054 27568 30126
rect 27528 30048 27580 30054
rect 27528 29990 27580 29996
rect 27528 29776 27580 29782
rect 27724 29730 27752 30670
rect 27580 29724 27752 29730
rect 27528 29718 27752 29724
rect 27540 29702 27752 29718
rect 27434 29608 27490 29617
rect 27434 29543 27436 29552
rect 27488 29543 27490 29552
rect 27436 29514 27488 29520
rect 27710 29336 27766 29345
rect 27710 29271 27712 29280
rect 27764 29271 27766 29280
rect 27712 29242 27764 29248
rect 27436 29232 27488 29238
rect 27436 29174 27488 29180
rect 27448 27878 27476 29174
rect 27620 29028 27672 29034
rect 27620 28970 27672 28976
rect 27632 28762 27660 28970
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 27528 28552 27580 28558
rect 27528 28494 27580 28500
rect 27540 28218 27568 28494
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 27436 27872 27488 27878
rect 27436 27814 27488 27820
rect 27448 25838 27476 27814
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 27540 26450 27568 27066
rect 27528 26444 27580 26450
rect 27528 26386 27580 26392
rect 27436 25832 27488 25838
rect 27436 25774 27488 25780
rect 27540 25226 27568 26386
rect 27724 25906 27752 29242
rect 27802 29200 27858 29209
rect 27802 29135 27804 29144
rect 27856 29135 27858 29144
rect 27804 29106 27856 29112
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 27528 25220 27580 25226
rect 27528 25162 27580 25168
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 27160 23588 27212 23594
rect 27160 23530 27212 23536
rect 27068 22432 27120 22438
rect 27068 22374 27120 22380
rect 26700 22092 26752 22098
rect 26700 22034 26752 22040
rect 26712 21894 26740 22034
rect 27080 21962 27108 22374
rect 27068 21956 27120 21962
rect 27068 21898 27120 21904
rect 27172 21894 27200 23530
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27356 22098 27384 22578
rect 27344 22092 27396 22098
rect 27344 22034 27396 22040
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27172 21554 27200 21830
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27264 19922 27292 19994
rect 27344 19984 27396 19990
rect 27344 19926 27396 19932
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 27356 19854 27384 19926
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26804 18834 26832 19110
rect 27080 18834 27108 19654
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 27264 18358 27292 18566
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26988 17882 27016 18158
rect 26976 17876 27028 17882
rect 26976 17818 27028 17824
rect 26884 17536 26936 17542
rect 26884 17478 26936 17484
rect 26896 17338 26924 17478
rect 26884 17332 26936 17338
rect 26884 17274 26936 17280
rect 27712 17060 27764 17066
rect 27712 17002 27764 17008
rect 27724 16590 27752 17002
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27172 16114 27200 16526
rect 27264 16114 27292 16526
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27252 16108 27304 16114
rect 27252 16050 27304 16056
rect 26608 5092 26660 5098
rect 26608 5034 26660 5040
rect 26240 4752 26292 4758
rect 26240 4694 26292 4700
rect 26252 4554 26280 4694
rect 26240 4548 26292 4554
rect 26240 4490 26292 4496
rect 26976 4548 27028 4554
rect 26976 4490 27028 4496
rect 26240 3460 26292 3466
rect 26240 3402 26292 3408
rect 26252 2650 26280 3402
rect 26988 3058 27016 4490
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 26436 2446 26464 2926
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 26528 1306 26556 2382
rect 26436 1278 26556 1306
rect 26436 800 26464 1278
rect 27080 800 27108 2994
rect 27264 2514 27292 16050
rect 27724 4554 27752 16526
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27816 16114 27844 16390
rect 27804 16108 27856 16114
rect 27804 16050 27856 16056
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 27724 3602 27752 4490
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27252 2508 27304 2514
rect 27252 2450 27304 2456
rect 27908 2446 27936 35022
rect 28000 33114 28028 35142
rect 28078 35119 28134 35128
rect 28092 34542 28120 35119
rect 28184 34678 28212 35702
rect 28368 35698 28396 37062
rect 28356 35692 28408 35698
rect 28356 35634 28408 35640
rect 28264 35556 28316 35562
rect 28264 35498 28316 35504
rect 28276 35086 28304 35498
rect 28368 35086 28396 35634
rect 28264 35080 28316 35086
rect 28264 35022 28316 35028
rect 28356 35080 28408 35086
rect 28356 35022 28408 35028
rect 28172 34672 28224 34678
rect 28172 34614 28224 34620
rect 28080 34536 28132 34542
rect 28080 34478 28132 34484
rect 28184 34218 28212 34614
rect 28092 34190 28212 34218
rect 27988 33108 28040 33114
rect 27988 33050 28040 33056
rect 27988 32836 28040 32842
rect 27988 32778 28040 32784
rect 28000 31890 28028 32778
rect 27988 31884 28040 31890
rect 27988 31826 28040 31832
rect 28092 30734 28120 34190
rect 28276 33930 28304 35022
rect 28264 33924 28316 33930
rect 28264 33866 28316 33872
rect 28356 33108 28408 33114
rect 28356 33050 28408 33056
rect 28172 32904 28224 32910
rect 28172 32846 28224 32852
rect 28184 32434 28212 32846
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 28264 32292 28316 32298
rect 28264 32234 28316 32240
rect 28276 31822 28304 32234
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28276 30734 28304 31758
rect 28080 30728 28132 30734
rect 28080 30670 28132 30676
rect 28264 30728 28316 30734
rect 28264 30670 28316 30676
rect 28170 30288 28226 30297
rect 28170 30223 28172 30232
rect 28224 30223 28226 30232
rect 28172 30194 28224 30200
rect 28080 29844 28132 29850
rect 28080 29786 28132 29792
rect 27986 29744 28042 29753
rect 27986 29679 27988 29688
rect 28040 29679 28042 29688
rect 27988 29650 28040 29656
rect 28092 29646 28120 29786
rect 28184 29646 28212 30194
rect 28368 30138 28396 33050
rect 28460 31754 28488 46990
rect 29184 38344 29236 38350
rect 29184 38286 29236 38292
rect 29196 37874 29224 38286
rect 29184 37868 29236 37874
rect 29184 37810 29236 37816
rect 28724 37664 28776 37670
rect 28724 37606 28776 37612
rect 29276 37664 29328 37670
rect 29276 37606 29328 37612
rect 28736 36922 28764 37606
rect 29288 37194 29316 37606
rect 29276 37188 29328 37194
rect 29276 37130 29328 37136
rect 28724 36916 28776 36922
rect 28724 36858 28776 36864
rect 29000 36712 29052 36718
rect 29000 36654 29052 36660
rect 29828 36712 29880 36718
rect 29828 36654 29880 36660
rect 28540 36100 28592 36106
rect 28540 36042 28592 36048
rect 28552 35834 28580 36042
rect 28540 35828 28592 35834
rect 28540 35770 28592 35776
rect 28540 35284 28592 35290
rect 28540 35226 28592 35232
rect 28908 35284 28960 35290
rect 28908 35226 28960 35232
rect 28552 32042 28580 35226
rect 28724 35216 28776 35222
rect 28724 35158 28776 35164
rect 28632 35080 28684 35086
rect 28736 35057 28764 35158
rect 28632 35022 28684 35028
rect 28722 35048 28778 35057
rect 28644 34066 28672 35022
rect 28722 34983 28778 34992
rect 28920 34746 28948 35226
rect 28908 34740 28960 34746
rect 28908 34682 28960 34688
rect 28816 34604 28868 34610
rect 28816 34546 28868 34552
rect 28828 34474 28856 34546
rect 28816 34468 28868 34474
rect 28816 34410 28868 34416
rect 28828 34202 28856 34410
rect 28816 34196 28868 34202
rect 28816 34138 28868 34144
rect 28632 34060 28684 34066
rect 28632 34002 28684 34008
rect 28724 33856 28776 33862
rect 28724 33798 28776 33804
rect 28736 32842 28764 33798
rect 28828 32910 28856 34138
rect 28908 33924 28960 33930
rect 28908 33866 28960 33872
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 28724 32836 28776 32842
rect 28724 32778 28776 32784
rect 28552 32014 28856 32042
rect 28460 31726 28580 31754
rect 28446 30288 28502 30297
rect 28446 30223 28502 30232
rect 28460 30190 28488 30223
rect 28276 30110 28396 30138
rect 28448 30184 28500 30190
rect 28448 30126 28500 30132
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 28172 29640 28224 29646
rect 28172 29582 28224 29588
rect 28092 29306 28120 29582
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 28276 28082 28304 30110
rect 28356 30048 28408 30054
rect 28356 29990 28408 29996
rect 28368 29170 28396 29990
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28264 28076 28316 28082
rect 28264 28018 28316 28024
rect 28080 28008 28132 28014
rect 28080 27950 28132 27956
rect 28092 24818 28120 27950
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 28184 25770 28212 26930
rect 28264 26308 28316 26314
rect 28316 26268 28396 26296
rect 28264 26250 28316 26256
rect 28172 25764 28224 25770
rect 28172 25706 28224 25712
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28368 24750 28396 26268
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28276 22710 28304 23054
rect 28264 22704 28316 22710
rect 28264 22646 28316 22652
rect 27988 22568 28040 22574
rect 27988 22510 28040 22516
rect 28000 22166 28028 22510
rect 27988 22160 28040 22166
rect 27988 22102 28040 22108
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28184 21622 28212 21966
rect 28172 21616 28224 21622
rect 28172 21558 28224 21564
rect 28184 21010 28212 21558
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28276 20942 28304 22646
rect 28354 21448 28410 21457
rect 28354 21383 28356 21392
rect 28408 21383 28410 21392
rect 28356 21354 28408 21360
rect 28552 21010 28580 31726
rect 28724 31680 28776 31686
rect 28724 31622 28776 31628
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28644 29850 28672 30670
rect 28736 30258 28764 31622
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28632 29844 28684 29850
rect 28632 29786 28684 29792
rect 28632 28688 28684 28694
rect 28632 28630 28684 28636
rect 28644 28422 28672 28630
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28632 25900 28684 25906
rect 28632 25842 28684 25848
rect 28644 25362 28672 25842
rect 28632 25356 28684 25362
rect 28632 25298 28684 25304
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 28644 23730 28672 24142
rect 28632 23724 28684 23730
rect 28632 23666 28684 23672
rect 28540 21004 28592 21010
rect 28540 20946 28592 20952
rect 28264 20936 28316 20942
rect 28264 20878 28316 20884
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28460 20466 28488 20810
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 28644 20058 28672 23666
rect 28724 22976 28776 22982
rect 28724 22918 28776 22924
rect 28736 22642 28764 22918
rect 28724 22636 28776 22642
rect 28724 22578 28776 22584
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28736 21622 28764 21830
rect 28724 21616 28776 21622
rect 28724 21558 28776 21564
rect 28736 21350 28764 21558
rect 28724 21344 28776 21350
rect 28724 21286 28776 21292
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 28644 19378 28672 19994
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28276 18358 28304 19314
rect 28264 18352 28316 18358
rect 28264 18294 28316 18300
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 28000 16250 28028 17138
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 28092 16658 28120 16934
rect 28080 16652 28132 16658
rect 28080 16594 28132 16600
rect 28276 16250 28304 17138
rect 28552 16794 28580 17138
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 27988 16244 28040 16250
rect 27988 16186 28040 16192
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28552 12434 28580 16730
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 28644 16114 28672 16458
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28736 16046 28764 16390
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28552 12406 28764 12434
rect 28736 4146 28764 12406
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28828 2650 28856 32014
rect 28920 28762 28948 33866
rect 29012 33454 29040 36654
rect 29840 36378 29868 36654
rect 29828 36372 29880 36378
rect 29828 36314 29880 36320
rect 29828 36168 29880 36174
rect 29828 36110 29880 36116
rect 29840 35834 29868 36110
rect 29828 35828 29880 35834
rect 29828 35770 29880 35776
rect 29460 35692 29512 35698
rect 29460 35634 29512 35640
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 29104 35086 29132 35566
rect 29092 35080 29144 35086
rect 29092 35022 29144 35028
rect 29368 34536 29420 34542
rect 29368 34478 29420 34484
rect 29276 33856 29328 33862
rect 29276 33798 29328 33804
rect 29288 33590 29316 33798
rect 29276 33584 29328 33590
rect 29276 33526 29328 33532
rect 29000 33448 29052 33454
rect 29000 33390 29052 33396
rect 29276 33448 29328 33454
rect 29276 33390 29328 33396
rect 29012 33114 29040 33390
rect 29000 33108 29052 33114
rect 29000 33050 29052 33056
rect 29012 32026 29040 33050
rect 29288 33046 29316 33390
rect 29276 33040 29328 33046
rect 29276 32982 29328 32988
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 29000 32020 29052 32026
rect 29000 31962 29052 31968
rect 29012 30802 29040 31962
rect 29104 30870 29132 32370
rect 29380 32366 29408 34478
rect 29368 32360 29420 32366
rect 29368 32302 29420 32308
rect 29472 31657 29500 35634
rect 30104 35080 30156 35086
rect 30104 35022 30156 35028
rect 30116 34610 30144 35022
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 30116 34202 30144 34546
rect 30104 34196 30156 34202
rect 30104 34138 30156 34144
rect 29552 33992 29604 33998
rect 29552 33934 29604 33940
rect 30012 33992 30064 33998
rect 30012 33934 30064 33940
rect 29564 33046 29592 33934
rect 30024 33454 30052 33934
rect 30012 33448 30064 33454
rect 30012 33390 30064 33396
rect 29552 33040 29604 33046
rect 29552 32982 29604 32988
rect 29920 32224 29972 32230
rect 29920 32166 29972 32172
rect 29932 31822 29960 32166
rect 30024 31822 30052 33390
rect 29920 31816 29972 31822
rect 29920 31758 29972 31764
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30208 31754 30236 47126
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49314 41318 50000
rect 40788 49286 41318 49314
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 31576 47048 31628 47054
rect 31576 46990 31628 46996
rect 31588 41414 31616 46990
rect 32036 46640 32088 46646
rect 32036 46582 32088 46588
rect 32232 46594 32260 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 31496 41386 31616 41414
rect 32048 41414 32076 46582
rect 32232 46566 32352 46594
rect 32324 46510 32352 46566
rect 32312 46504 32364 46510
rect 32312 46446 32364 46452
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 38028 45554 38056 49200
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38200 45960 38252 45966
rect 38200 45902 38252 45908
rect 38212 45626 38240 45902
rect 38200 45620 38252 45626
rect 38200 45562 38252 45568
rect 37292 45526 38056 45554
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 32048 41386 32260 41414
rect 31024 37868 31076 37874
rect 31024 37810 31076 37816
rect 31036 37262 31064 37810
rect 31024 37256 31076 37262
rect 31024 37198 31076 37204
rect 30840 37120 30892 37126
rect 30840 37062 30892 37068
rect 30852 36854 30880 37062
rect 30840 36848 30892 36854
rect 30840 36790 30892 36796
rect 31036 36174 31064 37198
rect 31116 36576 31168 36582
rect 31116 36518 31168 36524
rect 31300 36576 31352 36582
rect 31300 36518 31352 36524
rect 30840 36168 30892 36174
rect 30840 36110 30892 36116
rect 31024 36168 31076 36174
rect 31024 36110 31076 36116
rect 30852 35698 30880 36110
rect 30932 35828 30984 35834
rect 30932 35770 30984 35776
rect 30380 35692 30432 35698
rect 30380 35634 30432 35640
rect 30840 35692 30892 35698
rect 30840 35634 30892 35640
rect 30288 34672 30340 34678
rect 30288 34614 30340 34620
rect 30300 34218 30328 34614
rect 30392 34406 30420 35634
rect 30564 35012 30616 35018
rect 30564 34954 30616 34960
rect 30472 34672 30524 34678
rect 30472 34614 30524 34620
rect 30484 34474 30512 34614
rect 30472 34468 30524 34474
rect 30472 34410 30524 34416
rect 30576 34406 30604 34954
rect 30852 34746 30880 35634
rect 30944 35086 30972 35770
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 31036 35086 31064 35430
rect 30932 35080 30984 35086
rect 30932 35022 30984 35028
rect 31024 35080 31076 35086
rect 31024 35022 31076 35028
rect 30840 34740 30892 34746
rect 30840 34682 30892 34688
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 30656 34468 30708 34474
rect 30656 34410 30708 34416
rect 30380 34400 30432 34406
rect 30380 34342 30432 34348
rect 30564 34400 30616 34406
rect 30564 34342 30616 34348
rect 30300 34190 30512 34218
rect 30380 33516 30432 33522
rect 30380 33458 30432 33464
rect 30392 32570 30420 33458
rect 30484 32570 30512 34190
rect 30668 34134 30696 34410
rect 30656 34128 30708 34134
rect 30656 34070 30708 34076
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30380 32564 30432 32570
rect 30380 32506 30432 32512
rect 30472 32564 30524 32570
rect 30472 32506 30524 32512
rect 30576 31754 30604 33798
rect 30668 33318 30696 34070
rect 30852 33998 30880 34546
rect 31036 34542 31064 35022
rect 31024 34536 31076 34542
rect 31024 34478 31076 34484
rect 30840 33992 30892 33998
rect 30840 33934 30892 33940
rect 30656 33312 30708 33318
rect 30656 33254 30708 33260
rect 30668 33046 30696 33254
rect 30656 33040 30708 33046
rect 30656 32982 30708 32988
rect 30656 32836 30708 32842
rect 30656 32778 30708 32784
rect 30748 32836 30800 32842
rect 30748 32778 30800 32784
rect 30208 31726 30328 31754
rect 29458 31648 29514 31657
rect 29380 31606 29458 31634
rect 29092 30864 29144 30870
rect 29092 30806 29144 30812
rect 29000 30796 29052 30802
rect 29000 30738 29052 30744
rect 29104 30260 29132 30806
rect 29276 30320 29328 30326
rect 29274 30288 29276 30297
rect 29328 30288 29330 30297
rect 29092 30254 29144 30260
rect 29092 30196 29144 30202
rect 29184 30252 29236 30258
rect 29274 30223 29330 30232
rect 29184 30194 29236 30200
rect 29196 30138 29224 30194
rect 29196 30110 29316 30138
rect 29184 30048 29236 30054
rect 29184 29990 29236 29996
rect 28908 28756 28960 28762
rect 28908 28698 28960 28704
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 28920 26586 28948 26930
rect 28908 26580 28960 26586
rect 28908 26522 28960 26528
rect 29196 26382 29224 29990
rect 29288 29578 29316 30110
rect 29380 30054 29408 31606
rect 29458 31583 29514 31592
rect 29828 30660 29880 30666
rect 29828 30602 29880 30608
rect 29840 30394 29868 30602
rect 29828 30388 29880 30394
rect 29828 30330 29880 30336
rect 29460 30252 29512 30258
rect 29460 30194 29512 30200
rect 29368 30048 29420 30054
rect 29368 29990 29420 29996
rect 29276 29572 29328 29578
rect 29276 29514 29328 29520
rect 29184 26376 29236 26382
rect 29184 26318 29236 26324
rect 29288 25430 29316 29514
rect 29368 27396 29420 27402
rect 29368 27338 29420 27344
rect 29276 25424 29328 25430
rect 29276 25366 29328 25372
rect 29092 22568 29144 22574
rect 29092 22510 29144 22516
rect 29000 21956 29052 21962
rect 29000 21898 29052 21904
rect 29012 21570 29040 21898
rect 29104 21894 29132 22510
rect 29184 22024 29236 22030
rect 29184 21966 29236 21972
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 29196 21622 29224 21966
rect 29184 21616 29236 21622
rect 28920 21554 29132 21570
rect 29184 21558 29236 21564
rect 28908 21548 29132 21554
rect 28960 21542 29132 21548
rect 28908 21490 28960 21496
rect 29000 21344 29052 21350
rect 29000 21286 29052 21292
rect 29012 20534 29040 21286
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 29104 20398 29132 21542
rect 29092 20392 29144 20398
rect 29092 20334 29144 20340
rect 28908 19168 28960 19174
rect 28908 19110 28960 19116
rect 28920 18698 28948 19110
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 28908 18692 28960 18698
rect 28908 18634 28960 18640
rect 29012 17134 29040 18906
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 28908 16448 28960 16454
rect 28908 16390 28960 16396
rect 28920 16182 28948 16390
rect 28908 16176 28960 16182
rect 28908 16118 28960 16124
rect 29196 16114 29224 16934
rect 29184 16108 29236 16114
rect 29184 16050 29236 16056
rect 29380 3058 29408 27338
rect 29472 22094 29500 30194
rect 30104 30048 30156 30054
rect 30104 29990 30156 29996
rect 29734 29608 29790 29617
rect 29734 29543 29790 29552
rect 29748 29102 29776 29543
rect 30012 29164 30064 29170
rect 30012 29106 30064 29112
rect 29736 29096 29788 29102
rect 30024 29073 30052 29106
rect 29736 29038 29788 29044
rect 30010 29064 30066 29073
rect 30010 28999 30066 29008
rect 29552 28960 29604 28966
rect 29552 28902 29604 28908
rect 29644 28960 29696 28966
rect 29644 28902 29696 28908
rect 29564 28150 29592 28902
rect 29656 28694 29684 28902
rect 29644 28688 29696 28694
rect 29644 28630 29696 28636
rect 30116 28558 30144 29990
rect 30104 28552 30156 28558
rect 30104 28494 30156 28500
rect 29828 28416 29880 28422
rect 29828 28358 29880 28364
rect 29552 28144 29604 28150
rect 29552 28086 29604 28092
rect 29552 28008 29604 28014
rect 29552 27950 29604 27956
rect 29564 27606 29592 27950
rect 29552 27600 29604 27606
rect 29552 27542 29604 27548
rect 29840 27470 29868 28358
rect 29828 27464 29880 27470
rect 29828 27406 29880 27412
rect 29552 26308 29604 26314
rect 29552 26250 29604 26256
rect 29564 25974 29592 26250
rect 29552 25968 29604 25974
rect 29552 25910 29604 25916
rect 29564 25702 29592 25910
rect 29920 25900 29972 25906
rect 29920 25842 29972 25848
rect 29552 25696 29604 25702
rect 29552 25638 29604 25644
rect 29564 25294 29592 25638
rect 29552 25288 29604 25294
rect 29552 25230 29604 25236
rect 29644 24812 29696 24818
rect 29644 24754 29696 24760
rect 29656 24410 29684 24754
rect 29644 24404 29696 24410
rect 29644 24346 29696 24352
rect 29644 22704 29696 22710
rect 29644 22646 29696 22652
rect 29656 22098 29684 22646
rect 29472 22066 29592 22094
rect 29460 22024 29512 22030
rect 29460 21966 29512 21972
rect 29472 20942 29500 21966
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29460 17128 29512 17134
rect 29460 17070 29512 17076
rect 29472 16046 29500 17070
rect 29460 16040 29512 16046
rect 29460 15982 29512 15988
rect 29564 12434 29592 22066
rect 29644 22092 29696 22098
rect 29644 22034 29696 22040
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 29748 21457 29776 21490
rect 29734 21448 29790 21457
rect 29734 21383 29790 21392
rect 29736 20800 29788 20806
rect 29736 20742 29788 20748
rect 29748 20534 29776 20742
rect 29736 20528 29788 20534
rect 29736 20470 29788 20476
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 29840 16250 29868 16526
rect 29828 16244 29880 16250
rect 29828 16186 29880 16192
rect 29472 12406 29592 12434
rect 29472 3942 29500 12406
rect 29932 8838 29960 25842
rect 30196 23112 30248 23118
rect 30196 23054 30248 23060
rect 30208 22438 30236 23054
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30012 22092 30064 22098
rect 30012 22034 30064 22040
rect 30024 18766 30052 22034
rect 30300 21622 30328 31726
rect 30484 31726 30604 31754
rect 30484 30326 30512 31726
rect 30564 31204 30616 31210
rect 30668 31192 30696 32778
rect 30760 32502 30788 32778
rect 30748 32496 30800 32502
rect 30748 32438 30800 32444
rect 30616 31164 30696 31192
rect 30564 31146 30616 31152
rect 30472 30320 30524 30326
rect 30472 30262 30524 30268
rect 30484 29714 30512 30262
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30576 29646 30604 31146
rect 30852 30802 30880 33934
rect 31024 32768 31076 32774
rect 31024 32710 31076 32716
rect 31036 32570 31064 32710
rect 31024 32564 31076 32570
rect 31024 32506 31076 32512
rect 30932 32496 30984 32502
rect 30932 32438 30984 32444
rect 30840 30796 30892 30802
rect 30840 30738 30892 30744
rect 30944 30410 30972 32438
rect 31128 32434 31156 36518
rect 31312 36242 31340 36518
rect 31300 36236 31352 36242
rect 31300 36178 31352 36184
rect 31312 35766 31340 36178
rect 31300 35760 31352 35766
rect 31300 35702 31352 35708
rect 31208 34740 31260 34746
rect 31208 34682 31260 34688
rect 31220 32722 31248 34682
rect 31392 34060 31444 34066
rect 31392 34002 31444 34008
rect 31300 33856 31352 33862
rect 31300 33798 31352 33804
rect 31312 32910 31340 33798
rect 31404 33046 31432 34002
rect 31392 33040 31444 33046
rect 31392 32982 31444 32988
rect 31300 32904 31352 32910
rect 31300 32846 31352 32852
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31404 32722 31432 32846
rect 31220 32694 31432 32722
rect 31496 32434 31524 41386
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 32036 35488 32088 35494
rect 32036 35430 32088 35436
rect 31852 35284 31904 35290
rect 31852 35226 31904 35232
rect 31864 35086 31892 35226
rect 31944 35216 31996 35222
rect 31944 35158 31996 35164
rect 31668 35080 31720 35086
rect 31668 35022 31720 35028
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 31576 32904 31628 32910
rect 31576 32846 31628 32852
rect 31588 32570 31616 32846
rect 31576 32564 31628 32570
rect 31576 32506 31628 32512
rect 31116 32428 31168 32434
rect 31116 32370 31168 32376
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31128 31754 31156 32370
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31128 31726 31248 31754
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 31116 31136 31168 31142
rect 31116 31078 31168 31084
rect 31036 30870 31064 31078
rect 31024 30864 31076 30870
rect 31024 30806 31076 30812
rect 31128 30666 31156 31078
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 30760 30382 30972 30410
rect 30760 29782 30788 30382
rect 30932 30252 30984 30258
rect 30932 30194 30984 30200
rect 30840 30048 30892 30054
rect 30840 29990 30892 29996
rect 30748 29776 30800 29782
rect 30748 29718 30800 29724
rect 30564 29640 30616 29646
rect 30564 29582 30616 29588
rect 30760 29306 30788 29718
rect 30852 29714 30880 29990
rect 30944 29782 30972 30194
rect 30932 29776 30984 29782
rect 30932 29718 30984 29724
rect 30840 29708 30892 29714
rect 30840 29650 30892 29656
rect 30748 29300 30800 29306
rect 30748 29242 30800 29248
rect 30748 29164 30800 29170
rect 30748 29106 30800 29112
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30392 28014 30420 28494
rect 30656 28484 30708 28490
rect 30656 28426 30708 28432
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30668 27062 30696 28426
rect 30760 28064 30788 29106
rect 30944 28558 30972 29718
rect 30932 28552 30984 28558
rect 30932 28494 30984 28500
rect 30944 28150 30972 28494
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 30932 28144 30984 28150
rect 30932 28086 30984 28092
rect 30840 28076 30892 28082
rect 30760 28036 30840 28064
rect 30840 28018 30892 28024
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 30392 25888 30420 26386
rect 30852 26314 30880 28018
rect 31036 27606 31064 28358
rect 31024 27600 31076 27606
rect 31024 27542 31076 27548
rect 31220 27402 31248 31726
rect 31496 31278 31524 31758
rect 31484 31272 31536 31278
rect 31484 31214 31536 31220
rect 31392 30252 31444 30258
rect 31392 30194 31444 30200
rect 31404 29170 31432 30194
rect 31496 29646 31524 31214
rect 31576 30660 31628 30666
rect 31576 30602 31628 30608
rect 31484 29640 31536 29646
rect 31484 29582 31536 29588
rect 31496 29510 31524 29582
rect 31484 29504 31536 29510
rect 31484 29446 31536 29452
rect 31588 29306 31616 30602
rect 31576 29300 31628 29306
rect 31576 29242 31628 29248
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31404 28626 31432 29106
rect 31392 28620 31444 28626
rect 31392 28562 31444 28568
rect 31680 28558 31708 35022
rect 31760 30932 31812 30938
rect 31760 30874 31812 30880
rect 31772 29306 31800 30874
rect 31864 29730 31892 35022
rect 31956 30802 31984 35158
rect 32048 35154 32076 35430
rect 32036 35148 32088 35154
rect 32036 35090 32088 35096
rect 32140 33114 32168 35566
rect 32128 33108 32180 33114
rect 32128 33050 32180 33056
rect 32036 33040 32088 33046
rect 32036 32982 32088 32988
rect 32048 32842 32076 32982
rect 32036 32836 32088 32842
rect 32036 32778 32088 32784
rect 32140 32434 32168 33050
rect 32128 32428 32180 32434
rect 32128 32370 32180 32376
rect 31944 30796 31996 30802
rect 31944 30738 31996 30744
rect 32036 30728 32088 30734
rect 32036 30670 32088 30676
rect 32048 30258 32076 30670
rect 32036 30252 32088 30258
rect 32036 30194 32088 30200
rect 32036 30048 32088 30054
rect 32036 29990 32088 29996
rect 31864 29702 31984 29730
rect 31760 29300 31812 29306
rect 31760 29242 31812 29248
rect 31956 28762 31984 29702
rect 32048 29578 32076 29990
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 32036 29572 32088 29578
rect 32036 29514 32088 29520
rect 31944 28756 31996 28762
rect 31944 28698 31996 28704
rect 31668 28552 31720 28558
rect 31668 28494 31720 28500
rect 31944 28552 31996 28558
rect 31944 28494 31996 28500
rect 31576 28484 31628 28490
rect 31576 28426 31628 28432
rect 31588 28082 31616 28426
rect 31576 28076 31628 28082
rect 31576 28018 31628 28024
rect 31956 27674 31984 28494
rect 32048 28218 32076 29514
rect 32140 29170 32168 29582
rect 32128 29164 32180 29170
rect 32128 29106 32180 29112
rect 32140 28626 32168 29106
rect 32128 28620 32180 28626
rect 32128 28562 32180 28568
rect 32232 28234 32260 41386
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 33140 36032 33192 36038
rect 33140 35974 33192 35980
rect 33152 35766 33180 35974
rect 33140 35760 33192 35766
rect 33140 35702 33192 35708
rect 32496 35624 32548 35630
rect 32496 35566 32548 35572
rect 32508 35290 32536 35566
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 32496 35284 32548 35290
rect 32496 35226 32548 35232
rect 32864 35148 32916 35154
rect 32864 35090 32916 35096
rect 32312 35080 32364 35086
rect 32312 35022 32364 35028
rect 32324 29617 32352 35022
rect 32588 32904 32640 32910
rect 32588 32846 32640 32852
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32416 32502 32444 32778
rect 32496 32768 32548 32774
rect 32496 32710 32548 32716
rect 32404 32496 32456 32502
rect 32404 32438 32456 32444
rect 32508 30938 32536 32710
rect 32600 32026 32628 32846
rect 32772 32224 32824 32230
rect 32772 32166 32824 32172
rect 32588 32020 32640 32026
rect 32588 31962 32640 31968
rect 32784 31822 32812 32166
rect 32588 31816 32640 31822
rect 32588 31758 32640 31764
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 32600 30954 32628 31758
rect 32496 30932 32548 30938
rect 32600 30926 32720 30954
rect 32496 30874 32548 30880
rect 32588 30796 32640 30802
rect 32588 30738 32640 30744
rect 32404 30184 32456 30190
rect 32404 30126 32456 30132
rect 32310 29608 32366 29617
rect 32310 29543 32366 29552
rect 32416 29510 32444 30126
rect 32496 29844 32548 29850
rect 32496 29786 32548 29792
rect 32508 29594 32536 29786
rect 32600 29714 32628 30738
rect 32692 30666 32720 30926
rect 32680 30660 32732 30666
rect 32680 30602 32732 30608
rect 32588 29708 32640 29714
rect 32588 29650 32640 29656
rect 32692 29594 32720 30602
rect 32772 30252 32824 30258
rect 32772 30194 32824 30200
rect 32508 29566 32720 29594
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32496 29504 32548 29510
rect 32496 29446 32548 29452
rect 32416 29170 32444 29446
rect 32508 29306 32536 29446
rect 32496 29300 32548 29306
rect 32496 29242 32548 29248
rect 32404 29164 32456 29170
rect 32404 29106 32456 29112
rect 32416 28762 32444 29106
rect 32404 28756 32456 28762
rect 32404 28698 32456 28704
rect 32036 28212 32088 28218
rect 32232 28206 32444 28234
rect 32036 28154 32088 28160
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32128 27872 32180 27878
rect 32128 27814 32180 27820
rect 31944 27668 31996 27674
rect 31944 27610 31996 27616
rect 32140 27470 32168 27814
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 32128 27464 32180 27470
rect 32128 27406 32180 27412
rect 31208 27396 31260 27402
rect 31208 27338 31260 27344
rect 31668 27396 31720 27402
rect 31668 27338 31720 27344
rect 31116 26988 31168 26994
rect 31116 26930 31168 26936
rect 30840 26308 30892 26314
rect 30840 26250 30892 26256
rect 30852 26042 30880 26250
rect 31128 26042 31156 26930
rect 31208 26784 31260 26790
rect 31208 26726 31260 26732
rect 30840 26036 30892 26042
rect 30840 25978 30892 25984
rect 31116 26036 31168 26042
rect 31116 25978 31168 25984
rect 30472 25900 30524 25906
rect 30392 25860 30472 25888
rect 30392 24750 30420 25860
rect 30472 25842 30524 25848
rect 30852 25158 30880 25978
rect 31116 25288 31168 25294
rect 31116 25230 31168 25236
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30392 24410 30420 24550
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30668 24342 30696 24550
rect 30656 24336 30708 24342
rect 30656 24278 30708 24284
rect 30288 21616 30340 21622
rect 30288 21558 30340 21564
rect 31128 21146 31156 25230
rect 31220 24818 31248 26726
rect 31680 26364 31708 27338
rect 31760 26376 31812 26382
rect 31680 26336 31760 26364
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31404 25362 31432 25842
rect 31680 25770 31708 26336
rect 31760 26318 31812 26324
rect 31956 26314 31984 27406
rect 32220 26988 32272 26994
rect 32220 26930 32272 26936
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 31944 26308 31996 26314
rect 31944 26250 31996 26256
rect 31668 25764 31720 25770
rect 31668 25706 31720 25712
rect 31392 25356 31444 25362
rect 31392 25298 31444 25304
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31312 24886 31340 25094
rect 31300 24880 31352 24886
rect 31300 24822 31352 24828
rect 31208 24812 31260 24818
rect 31208 24754 31260 24760
rect 31576 22092 31628 22098
rect 31576 22034 31628 22040
rect 31588 21622 31616 22034
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31116 21140 31168 21146
rect 31116 21082 31168 21088
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30024 18358 30052 18702
rect 30116 18358 30144 18702
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 30012 18352 30064 18358
rect 30012 18294 30064 18300
rect 30104 18352 30156 18358
rect 30104 18294 30156 18300
rect 30024 17066 30052 18294
rect 30208 18204 30236 18566
rect 30288 18216 30340 18222
rect 30208 18176 30288 18204
rect 30208 17678 30236 18176
rect 30288 18158 30340 18164
rect 30392 18154 30420 20878
rect 31024 20868 31076 20874
rect 31024 20810 31076 20816
rect 31036 20058 31064 20810
rect 31024 20052 31076 20058
rect 31024 19994 31076 20000
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 31300 19848 31352 19854
rect 31300 19790 31352 19796
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30300 17338 30328 17682
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30012 17060 30064 17066
rect 30012 17002 30064 17008
rect 30484 13938 30512 19790
rect 31312 19514 31340 19790
rect 31300 19508 31352 19514
rect 31300 19450 31352 19456
rect 31944 19508 31996 19514
rect 31944 19450 31996 19456
rect 31208 19372 31260 19378
rect 31208 19314 31260 19320
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 31128 17746 31156 18702
rect 31220 18358 31248 19314
rect 31208 18352 31260 18358
rect 31208 18294 31260 18300
rect 31956 18222 31984 19450
rect 31944 18216 31996 18222
rect 31944 18158 31996 18164
rect 31116 17740 31168 17746
rect 31116 17682 31168 17688
rect 30656 17060 30708 17066
rect 30656 17002 30708 17008
rect 30668 16658 30696 17002
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30472 13932 30524 13938
rect 30472 13874 30524 13880
rect 32048 12646 32076 26318
rect 32128 26308 32180 26314
rect 32128 26250 32180 26256
rect 32140 25906 32168 26250
rect 32232 26042 32260 26930
rect 32220 26036 32272 26042
rect 32220 25978 32272 25984
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 32220 25764 32272 25770
rect 32220 25706 32272 25712
rect 32232 25430 32260 25706
rect 32220 25424 32272 25430
rect 32220 25366 32272 25372
rect 32324 25362 32352 28018
rect 32312 25356 32364 25362
rect 32312 25298 32364 25304
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32128 24744 32180 24750
rect 32128 24686 32180 24692
rect 32140 24614 32168 24686
rect 32232 24614 32260 24754
rect 32128 24608 32180 24614
rect 32128 24550 32180 24556
rect 32220 24608 32272 24614
rect 32220 24550 32272 24556
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 32140 23866 32168 24142
rect 32128 23860 32180 23866
rect 32128 23802 32180 23808
rect 32232 23746 32260 24550
rect 32324 24274 32352 25298
rect 32416 24818 32444 28206
rect 32508 25770 32536 29242
rect 32692 28558 32720 29566
rect 32680 28552 32732 28558
rect 32680 28494 32732 28500
rect 32588 28416 32640 28422
rect 32588 28358 32640 28364
rect 32600 28150 32628 28358
rect 32588 28144 32640 28150
rect 32588 28086 32640 28092
rect 32784 26586 32812 30194
rect 32680 26580 32732 26586
rect 32680 26522 32732 26528
rect 32772 26580 32824 26586
rect 32772 26522 32824 26528
rect 32588 26444 32640 26450
rect 32588 26386 32640 26392
rect 32600 25906 32628 26386
rect 32692 25906 32720 26522
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 32680 25900 32732 25906
rect 32680 25842 32732 25848
rect 32496 25764 32548 25770
rect 32496 25706 32548 25712
rect 32600 25226 32628 25842
rect 32588 25220 32640 25226
rect 32588 25162 32640 25168
rect 32404 24812 32456 24818
rect 32404 24754 32456 24760
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32312 24268 32364 24274
rect 32312 24210 32364 24216
rect 32140 23718 32260 23746
rect 32508 23730 32536 24754
rect 32600 24410 32628 25162
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 32496 23724 32548 23730
rect 32140 20466 32168 23718
rect 32496 23666 32548 23672
rect 32220 23044 32272 23050
rect 32220 22986 32272 22992
rect 32232 22778 32260 22986
rect 32220 22772 32272 22778
rect 32220 22714 32272 22720
rect 32404 21956 32456 21962
rect 32404 21898 32456 21904
rect 32416 21690 32444 21898
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32404 21344 32456 21350
rect 32404 21286 32456 21292
rect 32128 20460 32180 20466
rect 32128 20402 32180 20408
rect 32140 19378 32168 20402
rect 32220 20256 32272 20262
rect 32220 20198 32272 20204
rect 32232 19718 32260 20198
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32220 19168 32272 19174
rect 32220 19110 32272 19116
rect 32232 18834 32260 19110
rect 32220 18828 32272 18834
rect 32220 18770 32272 18776
rect 32312 18828 32364 18834
rect 32312 18770 32364 18776
rect 32324 18358 32352 18770
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32036 12640 32088 12646
rect 32036 12582 32088 12588
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 32220 4072 32272 4078
rect 32220 4014 32272 4020
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 30932 3664 30984 3670
rect 30932 3606 30984 3612
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28368 800 28396 2382
rect 29656 800 29684 2382
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 29748 2038 29776 2246
rect 29736 2032 29788 2038
rect 29736 1974 29788 1980
rect 30944 800 30972 3606
rect 32232 800 32260 4014
rect 32416 2378 32444 21286
rect 32772 3596 32824 3602
rect 32772 3538 32824 3544
rect 32784 3194 32812 3538
rect 32772 3188 32824 3194
rect 32772 3130 32824 3136
rect 32404 2372 32456 2378
rect 32404 2314 32456 2320
rect 32876 1970 32904 35090
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 33416 32496 33468 32502
rect 33416 32438 33468 32444
rect 33428 32026 33456 32438
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 33416 32020 33468 32026
rect 33416 31962 33468 31968
rect 34612 31816 34664 31822
rect 34612 31758 34664 31764
rect 33048 30796 33100 30802
rect 33048 30738 33100 30744
rect 33060 30054 33088 30738
rect 33692 30728 33744 30734
rect 33692 30670 33744 30676
rect 33704 30258 33732 30670
rect 34520 30660 34572 30666
rect 34520 30602 34572 30608
rect 33876 30592 33928 30598
rect 33876 30534 33928 30540
rect 33416 30252 33468 30258
rect 33416 30194 33468 30200
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33692 30252 33744 30258
rect 33692 30194 33744 30200
rect 33048 30048 33100 30054
rect 33048 29990 33100 29996
rect 32956 29640 33008 29646
rect 32956 29582 33008 29588
rect 32968 29306 32996 29582
rect 32956 29300 33008 29306
rect 32956 29242 33008 29248
rect 33060 29170 33088 29990
rect 33428 29850 33456 30194
rect 33416 29844 33468 29850
rect 33416 29786 33468 29792
rect 33520 29646 33548 30194
rect 33888 29782 33916 30534
rect 34532 30326 34560 30602
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 34624 30258 34652 31758
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35992 30660 36044 30666
rect 35992 30602 36044 30608
rect 36004 30326 36032 30602
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 33968 30252 34020 30258
rect 33968 30194 34020 30200
rect 34612 30252 34664 30258
rect 34612 30194 34664 30200
rect 33876 29776 33928 29782
rect 33876 29718 33928 29724
rect 33508 29640 33560 29646
rect 33508 29582 33560 29588
rect 33600 29640 33652 29646
rect 33876 29640 33928 29646
rect 33600 29582 33652 29588
rect 33874 29608 33876 29617
rect 33980 29628 34008 30194
rect 34152 30184 34204 30190
rect 34152 30126 34204 30132
rect 33928 29608 34008 29628
rect 33930 29600 34008 29608
rect 33612 29306 33640 29582
rect 33874 29543 33930 29552
rect 33600 29300 33652 29306
rect 33600 29242 33652 29248
rect 33784 29300 33836 29306
rect 33784 29242 33836 29248
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 33508 28960 33560 28966
rect 33508 28902 33560 28908
rect 32956 28620 33008 28626
rect 32956 28562 33008 28568
rect 32968 28218 32996 28562
rect 32956 28212 33008 28218
rect 32956 28154 33008 28160
rect 33520 26586 33548 28902
rect 33600 28144 33652 28150
rect 33600 28086 33652 28092
rect 33612 27606 33640 28086
rect 33600 27600 33652 27606
rect 33600 27542 33652 27548
rect 33508 26580 33560 26586
rect 33508 26522 33560 26528
rect 33692 26444 33744 26450
rect 33692 26386 33744 26392
rect 33048 26308 33100 26314
rect 33048 26250 33100 26256
rect 33060 25974 33088 26250
rect 33048 25968 33100 25974
rect 33048 25910 33100 25916
rect 33060 25838 33088 25910
rect 33704 25906 33732 26386
rect 33796 26382 33824 29242
rect 33968 26512 34020 26518
rect 33968 26454 34020 26460
rect 33784 26376 33836 26382
rect 33784 26318 33836 26324
rect 33980 25906 34008 26454
rect 33692 25900 33744 25906
rect 33692 25842 33744 25848
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 33324 25696 33376 25702
rect 33324 25638 33376 25644
rect 33336 25362 33364 25638
rect 33704 25498 33732 25842
rect 33692 25492 33744 25498
rect 33692 25434 33744 25440
rect 33324 25356 33376 25362
rect 33324 25298 33376 25304
rect 33140 25220 33192 25226
rect 33140 25162 33192 25168
rect 33152 24818 33180 25162
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 33152 22642 33180 23054
rect 33784 22976 33836 22982
rect 33784 22918 33836 22924
rect 33796 22710 33824 22918
rect 33784 22704 33836 22710
rect 33784 22646 33836 22652
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33152 20942 33180 22578
rect 34164 22094 34192 30126
rect 34244 29504 34296 29510
rect 34244 29446 34296 29452
rect 34256 29238 34284 29446
rect 34244 29232 34296 29238
rect 34244 29174 34296 29180
rect 34624 29073 34652 30194
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34610 29064 34666 29073
rect 34610 28999 34666 29008
rect 34624 28558 34652 28999
rect 34808 28762 34836 29174
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 34612 28552 34664 28558
rect 34612 28494 34664 28500
rect 34624 27470 34652 28494
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34612 27464 34664 27470
rect 34612 27406 34664 27412
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35164 25220 35216 25226
rect 35164 25162 35216 25168
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34808 24886 34836 25094
rect 34796 24880 34848 24886
rect 34796 24822 34848 24828
rect 34808 24614 34836 24822
rect 35176 24818 35204 25162
rect 35164 24812 35216 24818
rect 35164 24754 35216 24760
rect 35176 24698 35204 24754
rect 35176 24670 35388 24698
rect 34796 24608 34848 24614
rect 34796 24550 34848 24556
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 35360 24274 35388 24670
rect 35348 24268 35400 24274
rect 35348 24210 35400 24216
rect 34612 24200 34664 24206
rect 34612 24142 34664 24148
rect 34520 24132 34572 24138
rect 34520 24074 34572 24080
rect 34532 23866 34560 24074
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34164 22066 34284 22094
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33980 21690 34008 21966
rect 34060 21956 34112 21962
rect 34060 21898 34112 21904
rect 33968 21684 34020 21690
rect 33968 21626 34020 21632
rect 33600 21344 33652 21350
rect 33600 21286 33652 21292
rect 33612 21078 33640 21286
rect 33600 21072 33652 21078
rect 33600 21014 33652 21020
rect 34072 21010 34100 21898
rect 34060 21004 34112 21010
rect 34060 20946 34112 20952
rect 33140 20936 33192 20942
rect 33140 20878 33192 20884
rect 33232 20800 33284 20806
rect 33232 20742 33284 20748
rect 33244 20534 33272 20742
rect 33232 20528 33284 20534
rect 33232 20470 33284 20476
rect 34060 19440 34112 19446
rect 34060 19382 34112 19388
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 33520 18358 33548 18702
rect 33508 18352 33560 18358
rect 33508 18294 33560 18300
rect 34072 18222 34100 19382
rect 34060 18216 34112 18222
rect 34060 18158 34112 18164
rect 33140 18080 33192 18086
rect 33140 18022 33192 18028
rect 33152 17746 33180 18022
rect 33140 17740 33192 17746
rect 33140 17682 33192 17688
rect 34072 17610 34100 18158
rect 34060 17604 34112 17610
rect 34060 17546 34112 17552
rect 34072 17338 34100 17546
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 32956 3664 33008 3670
rect 32956 3606 33008 3612
rect 32968 3058 32996 3606
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33152 3126 33180 3334
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 32956 3052 33008 3058
rect 32956 2994 33008 3000
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33140 2848 33192 2854
rect 33140 2790 33192 2796
rect 33152 2650 33180 2790
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 32864 1964 32916 1970
rect 32864 1906 32916 1912
rect 33520 800 33548 2926
rect 34256 2514 34284 22066
rect 34428 20392 34480 20398
rect 34428 20334 34480 20340
rect 34440 3398 34468 20334
rect 34624 18698 34652 24142
rect 35360 23730 35388 24210
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35360 23118 35388 23666
rect 35992 23588 36044 23594
rect 35992 23530 36044 23536
rect 35716 23316 35768 23322
rect 35716 23258 35768 23264
rect 35728 23186 35756 23258
rect 35716 23180 35768 23186
rect 35716 23122 35768 23128
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35072 21616 35124 21622
rect 34808 21564 35072 21570
rect 34808 21558 35124 21564
rect 34808 21554 35112 21558
rect 34796 21548 35112 21554
rect 34848 21542 35112 21548
rect 34796 21490 34848 21496
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35348 19236 35400 19242
rect 35348 19178 35400 19184
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35360 18970 35388 19178
rect 35348 18964 35400 18970
rect 35348 18906 35400 18912
rect 34612 18692 34664 18698
rect 34612 18634 34664 18640
rect 34796 18624 34848 18630
rect 34796 18566 34848 18572
rect 34808 18290 34836 18566
rect 34796 18284 34848 18290
rect 34796 18226 34848 18232
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 35360 17678 35388 18906
rect 35532 18760 35584 18766
rect 35532 18702 35584 18708
rect 35544 18154 35572 18702
rect 35532 18148 35584 18154
rect 35532 18090 35584 18096
rect 35544 17746 35572 18090
rect 35532 17740 35584 17746
rect 35532 17682 35584 17688
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 35072 17604 35124 17610
rect 35072 17546 35124 17552
rect 35084 17270 35112 17546
rect 35072 17264 35124 17270
rect 35072 17206 35124 17212
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35728 3466 35756 23122
rect 35808 21956 35860 21962
rect 35808 21898 35860 21904
rect 35820 21486 35848 21898
rect 35808 21480 35860 21486
rect 35808 21422 35860 21428
rect 36004 16590 36032 23530
rect 37292 22778 37320 45526
rect 38212 38214 38240 45562
rect 39960 45554 39988 49200
rect 40132 47184 40184 47190
rect 40132 47126 40184 47132
rect 39960 45526 40080 45554
rect 38660 44872 38712 44878
rect 38660 44814 38712 44820
rect 38568 44328 38620 44334
rect 38568 44270 38620 44276
rect 38580 43654 38608 44270
rect 38568 43648 38620 43654
rect 38568 43590 38620 43596
rect 38672 39574 38700 44814
rect 38752 44736 38804 44742
rect 38752 44678 38804 44684
rect 38764 44470 38792 44678
rect 38752 44464 38804 44470
rect 38752 44406 38804 44412
rect 40052 44334 40080 45526
rect 40040 44328 40092 44334
rect 40040 44270 40092 44276
rect 39672 40928 39724 40934
rect 39672 40870 39724 40876
rect 38660 39568 38712 39574
rect 38660 39510 38712 39516
rect 38200 38208 38252 38214
rect 38200 38150 38252 38156
rect 39684 23730 39712 40870
rect 40040 24608 40092 24614
rect 40040 24550 40092 24556
rect 40052 24274 40080 24550
rect 40040 24268 40092 24274
rect 40040 24210 40092 24216
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 39672 23724 39724 23730
rect 39672 23666 39724 23672
rect 39396 23656 39448 23662
rect 39396 23598 39448 23604
rect 37280 22772 37332 22778
rect 37280 22714 37332 22720
rect 36360 21616 36412 21622
rect 36360 21558 36412 21564
rect 38384 21616 38436 21622
rect 38384 21558 38436 21564
rect 35992 16584 36044 16590
rect 35992 16526 36044 16532
rect 35716 3460 35768 3466
rect 35716 3402 35768 3408
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 36372 2650 36400 21558
rect 37004 21412 37056 21418
rect 37004 21354 37056 21360
rect 37016 20874 37044 21354
rect 38396 21350 38424 21558
rect 38384 21344 38436 21350
rect 38384 21286 38436 21292
rect 37004 20868 37056 20874
rect 37004 20810 37056 20816
rect 36544 16584 36596 16590
rect 36544 16526 36596 16532
rect 36556 16250 36584 16526
rect 36544 16244 36596 16250
rect 36544 16186 36596 16192
rect 36556 12434 36584 16186
rect 36464 12406 36584 12434
rect 36464 3602 36492 12406
rect 37740 6724 37792 6730
rect 37740 6666 37792 6672
rect 37752 6458 37780 6666
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 37740 6316 37792 6322
rect 37740 6258 37792 6264
rect 37752 5370 37780 6258
rect 38396 6254 38424 21286
rect 39408 6866 39436 23598
rect 39856 23112 39908 23118
rect 39856 23054 39908 23060
rect 39488 23044 39540 23050
rect 39488 22986 39540 22992
rect 39500 22778 39528 22986
rect 39580 22976 39632 22982
rect 39580 22918 39632 22924
rect 39488 22772 39540 22778
rect 39488 22714 39540 22720
rect 39592 22642 39620 22918
rect 39580 22636 39632 22642
rect 39580 22578 39632 22584
rect 39868 22234 39896 23054
rect 40052 22642 40080 24074
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 40144 22234 40172 47126
rect 40224 47048 40276 47054
rect 40224 46990 40276 46996
rect 40236 29714 40264 46990
rect 40788 45554 40816 49286
rect 41206 49200 41318 49286
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49314 44538 50000
rect 44426 49286 44864 49314
rect 44426 49200 44538 49286
rect 41328 46368 41380 46374
rect 41328 46310 41380 46316
rect 41420 46368 41472 46374
rect 41420 46310 41472 46316
rect 41340 46034 41368 46310
rect 41432 46102 41460 46310
rect 41420 46096 41472 46102
rect 41420 46038 41472 46044
rect 41892 46034 41920 49200
rect 42536 46442 42564 49200
rect 43180 47122 43208 49200
rect 43168 47116 43220 47122
rect 43168 47058 43220 47064
rect 42800 46980 42852 46986
rect 42800 46922 42852 46928
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 42432 46164 42484 46170
rect 42432 46106 42484 46112
rect 41328 46028 41380 46034
rect 41328 45970 41380 45976
rect 41880 46028 41932 46034
rect 41880 45970 41932 45976
rect 41512 45892 41564 45898
rect 41512 45834 41564 45840
rect 41524 45626 41552 45834
rect 41512 45620 41564 45626
rect 41512 45562 41564 45568
rect 40512 45526 40816 45554
rect 40224 29708 40276 29714
rect 40224 29650 40276 29656
rect 40316 24268 40368 24274
rect 40316 24210 40368 24216
rect 40328 23798 40356 24210
rect 40316 23792 40368 23798
rect 40316 23734 40368 23740
rect 40512 23186 40540 45526
rect 42444 45490 42472 46106
rect 42628 45626 42656 46446
rect 42616 45620 42668 45626
rect 42616 45562 42668 45568
rect 41328 45484 41380 45490
rect 41328 45426 41380 45432
rect 42432 45484 42484 45490
rect 42432 45426 42484 45432
rect 41340 44334 41368 45426
rect 41328 44328 41380 44334
rect 41328 44270 41380 44276
rect 41340 38554 41368 44270
rect 42444 41138 42472 45426
rect 42812 45082 42840 46922
rect 43824 45966 43852 49200
rect 44836 47462 44864 49286
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 44824 47456 44876 47462
rect 44824 47398 44876 47404
rect 45112 47410 45140 49200
rect 45468 47456 45520 47462
rect 45112 47382 45416 47410
rect 45468 47398 45520 47404
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 46980 45152 46986
rect 45100 46922 45152 46928
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 44180 45892 44232 45898
rect 44180 45834 44232 45840
rect 42892 45484 42944 45490
rect 42892 45426 42944 45432
rect 42800 45076 42852 45082
rect 42800 45018 42852 45024
rect 42904 44878 42932 45426
rect 43260 45280 43312 45286
rect 43260 45222 43312 45228
rect 42892 44872 42944 44878
rect 42892 44814 42944 44820
rect 42432 41132 42484 41138
rect 42432 41074 42484 41080
rect 41328 38548 41380 38554
rect 41328 38490 41380 38496
rect 42444 26234 42472 41074
rect 42524 27668 42576 27674
rect 42524 27610 42576 27616
rect 42352 26206 42472 26234
rect 41052 24132 41104 24138
rect 41052 24074 41104 24080
rect 41064 23866 41092 24074
rect 41052 23860 41104 23866
rect 41052 23802 41104 23808
rect 42352 23322 42380 26206
rect 42340 23316 42392 23322
rect 42340 23258 42392 23264
rect 40500 23180 40552 23186
rect 40500 23122 40552 23128
rect 42432 23112 42484 23118
rect 42432 23054 42484 23060
rect 42444 22642 42472 23054
rect 42432 22636 42484 22642
rect 42432 22578 42484 22584
rect 40224 22568 40276 22574
rect 40224 22510 40276 22516
rect 40236 22234 40264 22510
rect 42536 22506 42564 27610
rect 42904 26234 42932 44814
rect 42812 26206 42932 26234
rect 42616 23724 42668 23730
rect 42616 23666 42668 23672
rect 42628 22506 42656 23666
rect 42524 22500 42576 22506
rect 42524 22442 42576 22448
rect 42616 22500 42668 22506
rect 42616 22442 42668 22448
rect 39856 22228 39908 22234
rect 39856 22170 39908 22176
rect 40132 22228 40184 22234
rect 40132 22170 40184 22176
rect 40224 22228 40276 22234
rect 40224 22170 40276 22176
rect 40038 22128 40094 22137
rect 40038 22063 40094 22072
rect 40052 22030 40080 22063
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 39948 21548 40000 21554
rect 40052 21536 40080 21966
rect 40144 21554 40172 22170
rect 42708 21684 42760 21690
rect 42708 21626 42760 21632
rect 42720 21593 42748 21626
rect 42706 21584 42762 21593
rect 40000 21508 40080 21536
rect 40132 21548 40184 21554
rect 39948 21490 40000 21496
rect 42706 21519 42762 21528
rect 40132 21490 40184 21496
rect 40132 21344 40184 21350
rect 40132 21286 40184 21292
rect 39396 6860 39448 6866
rect 39396 6802 39448 6808
rect 39408 6390 39436 6802
rect 38476 6384 38528 6390
rect 38476 6326 38528 6332
rect 39396 6384 39448 6390
rect 39396 6326 39448 6332
rect 38384 6248 38436 6254
rect 38384 6190 38436 6196
rect 37740 5364 37792 5370
rect 37740 5306 37792 5312
rect 37372 5024 37424 5030
rect 37372 4966 37424 4972
rect 36544 3936 36596 3942
rect 36544 3878 36596 3884
rect 36556 3670 36584 3878
rect 36544 3664 36596 3670
rect 36544 3606 36596 3612
rect 36452 3596 36504 3602
rect 36452 3538 36504 3544
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 37384 2582 37412 4966
rect 38396 4486 38424 6190
rect 38488 5234 38516 6326
rect 39212 6248 39264 6254
rect 39212 6190 39264 6196
rect 38476 5228 38528 5234
rect 38476 5170 38528 5176
rect 38384 4480 38436 4486
rect 38384 4422 38436 4428
rect 37372 2576 37424 2582
rect 37372 2518 37424 2524
rect 34244 2508 34296 2514
rect 34244 2450 34296 2456
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 36096 800 36124 2314
rect 38028 800 38056 2314
rect 38488 2310 38516 5170
rect 39120 5024 39172 5030
rect 39120 4966 39172 4972
rect 39132 4622 39160 4966
rect 39120 4616 39172 4622
rect 39120 4558 39172 4564
rect 38660 4480 38712 4486
rect 38660 4422 38712 4428
rect 38672 4146 38700 4422
rect 38660 4140 38712 4146
rect 38660 4082 38712 4088
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 39132 3194 39160 3470
rect 39120 3188 39172 3194
rect 39120 3130 39172 3136
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 39132 2650 39160 2994
rect 39224 2990 39252 6190
rect 39672 5228 39724 5234
rect 39672 5170 39724 5176
rect 39488 4276 39540 4282
rect 39488 4218 39540 4224
rect 39500 4010 39528 4218
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 39488 4004 39540 4010
rect 39488 3946 39540 3952
rect 39592 3942 39620 4014
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 39684 3738 39712 5170
rect 40144 4622 40172 21286
rect 42812 17678 42840 26206
rect 43272 23730 43300 45222
rect 44192 33386 44220 45834
rect 44456 45416 44508 45422
rect 44456 45358 44508 45364
rect 44468 44402 44496 45358
rect 44456 44396 44508 44402
rect 44456 44338 44508 44344
rect 45112 44266 45140 46922
rect 45204 46594 45232 46990
rect 45204 46566 45324 46594
rect 45192 46504 45244 46510
rect 45192 46446 45244 46452
rect 45100 44260 45152 44266
rect 45100 44202 45152 44208
rect 45204 43994 45232 46446
rect 45192 43988 45244 43994
rect 45192 43930 45244 43936
rect 45296 43314 45324 46566
rect 45388 45422 45416 47382
rect 45376 45416 45428 45422
rect 45376 45358 45428 45364
rect 45480 44878 45508 47398
rect 45560 46504 45612 46510
rect 45560 46446 45612 46452
rect 45468 44872 45520 44878
rect 45468 44814 45520 44820
rect 45572 44538 45600 46446
rect 45756 45966 45784 49200
rect 46400 47444 46428 49200
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46400 47416 46612 47444
rect 46386 47016 46442 47025
rect 46386 46951 46442 46960
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45744 45620 45796 45626
rect 45744 45562 45796 45568
rect 45652 44804 45704 44810
rect 45652 44746 45704 44752
rect 45560 44532 45612 44538
rect 45560 44474 45612 44480
rect 45284 43308 45336 43314
rect 45284 43250 45336 43256
rect 44180 33380 44232 33386
rect 44180 33322 44232 33328
rect 45664 27538 45692 44746
rect 45756 44402 45784 45562
rect 45928 44940 45980 44946
rect 45928 44882 45980 44888
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45940 43858 45968 44882
rect 46296 44872 46348 44878
rect 46296 44814 46348 44820
rect 46308 44470 46336 44814
rect 46296 44464 46348 44470
rect 46296 44406 46348 44412
rect 46204 44396 46256 44402
rect 46204 44338 46256 44344
rect 45928 43852 45980 43858
rect 45928 43794 45980 43800
rect 46216 33114 46244 44338
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 46204 33108 46256 33114
rect 46204 33050 46256 33056
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46308 31890 46336 32846
rect 46296 31884 46348 31890
rect 46296 31826 46348 31832
rect 46400 31090 46428 46951
rect 46480 46028 46532 46034
rect 46480 45970 46532 45976
rect 46492 43314 46520 45970
rect 46584 45558 46612 47416
rect 46860 46510 46888 47631
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 48044 47184 48096 47190
rect 48044 47126 48096 47132
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47216 46368 47268 46374
rect 47216 46310 47268 46316
rect 47308 46368 47360 46374
rect 47964 46345 47992 46514
rect 47308 46310 47360 46316
rect 47950 46336 48006 46345
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 46572 45552 46624 45558
rect 46572 45494 46624 45500
rect 47228 45490 47256 46310
rect 47216 45484 47268 45490
rect 47216 45426 47268 45432
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 46952 43858 46980 44134
rect 46940 43852 46992 43858
rect 46940 43794 46992 43800
rect 46480 43308 46532 43314
rect 46480 43250 46532 43256
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 46570 39536 46626 39545
rect 46570 39471 46626 39480
rect 46480 33108 46532 33114
rect 46480 33050 46532 33056
rect 46492 32434 46520 33050
rect 46480 32428 46532 32434
rect 46480 32370 46532 32376
rect 46480 32224 46532 32230
rect 46480 32166 46532 32172
rect 46492 31890 46520 32166
rect 46480 31884 46532 31890
rect 46480 31826 46532 31832
rect 46584 31090 46612 39471
rect 46940 38344 46992 38350
rect 46940 38286 46992 38292
rect 46952 37126 46980 38286
rect 46940 37120 46992 37126
rect 46940 37062 46992 37068
rect 47320 35894 47348 46310
rect 47950 46271 48006 46280
rect 47676 45892 47728 45898
rect 47676 45834 47728 45840
rect 47688 45558 47716 45834
rect 47676 45552 47728 45558
rect 47676 45494 47728 45500
rect 47492 45484 47544 45490
rect 47492 45426 47544 45432
rect 47504 37874 47532 45426
rect 47676 44804 47728 44810
rect 47676 44746 47728 44752
rect 47584 44736 47636 44742
rect 47584 44678 47636 44684
rect 47596 42226 47624 44678
rect 47688 44538 47716 44746
rect 47676 44532 47728 44538
rect 47676 44474 47728 44480
rect 47768 43104 47820 43110
rect 47768 43046 47820 43052
rect 47780 42770 47808 43046
rect 47768 42764 47820 42770
rect 47768 42706 47820 42712
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47584 42220 47636 42226
rect 47584 42162 47636 42168
rect 47492 37868 47544 37874
rect 47492 37810 47544 37816
rect 47320 35866 47440 35894
rect 47124 35488 47176 35494
rect 47124 35430 47176 35436
rect 47136 34066 47164 35430
rect 47216 34400 47268 34406
rect 47216 34342 47268 34348
rect 47124 34060 47176 34066
rect 47124 34002 47176 34008
rect 47228 33930 47256 34342
rect 47216 33924 47268 33930
rect 47216 33866 47268 33872
rect 46848 33516 46900 33522
rect 46848 33458 46900 33464
rect 47308 33516 47360 33522
rect 47308 33458 47360 33464
rect 46860 33425 46888 33458
rect 46846 33416 46902 33425
rect 46846 33351 46902 33360
rect 46940 33312 46992 33318
rect 46940 33254 46992 33260
rect 46848 32768 46900 32774
rect 46848 32710 46900 32716
rect 46860 32065 46888 32710
rect 46952 32570 46980 33254
rect 46940 32564 46992 32570
rect 46940 32506 46992 32512
rect 46846 32056 46902 32065
rect 46846 31991 46902 32000
rect 46662 31376 46718 31385
rect 46662 31311 46718 31320
rect 46032 31062 46428 31090
rect 46492 31062 46612 31090
rect 45836 28076 45888 28082
rect 45836 28018 45888 28024
rect 45652 27532 45704 27538
rect 45652 27474 45704 27480
rect 45650 26616 45706 26625
rect 45650 26551 45706 26560
rect 45008 24812 45060 24818
rect 45008 24754 45060 24760
rect 44364 24744 44416 24750
rect 44364 24686 44416 24692
rect 44376 24274 44404 24686
rect 44364 24268 44416 24274
rect 44364 24210 44416 24216
rect 45020 24206 45048 24754
rect 45100 24744 45152 24750
rect 45100 24686 45152 24692
rect 45376 24744 45428 24750
rect 45376 24686 45428 24692
rect 45008 24200 45060 24206
rect 45008 24142 45060 24148
rect 43260 23724 43312 23730
rect 43260 23666 43312 23672
rect 43904 23724 43956 23730
rect 43904 23666 43956 23672
rect 44088 23724 44140 23730
rect 44088 23666 44140 23672
rect 43272 22438 43300 23666
rect 43812 23520 43864 23526
rect 43812 23462 43864 23468
rect 43628 23180 43680 23186
rect 43628 23122 43680 23128
rect 43640 22642 43668 23122
rect 43824 23118 43852 23462
rect 43812 23112 43864 23118
rect 43812 23054 43864 23060
rect 43916 22642 43944 23666
rect 43996 22704 44048 22710
rect 44100 22658 44128 23666
rect 44048 22652 44128 22658
rect 43996 22646 44128 22652
rect 43536 22636 43588 22642
rect 43536 22578 43588 22584
rect 43628 22636 43680 22642
rect 43628 22578 43680 22584
rect 43904 22636 43956 22642
rect 44008 22630 44128 22646
rect 43904 22578 43956 22584
rect 43260 22432 43312 22438
rect 43260 22374 43312 22380
rect 43168 22160 43220 22166
rect 43168 22102 43220 22108
rect 43180 22030 43208 22102
rect 43272 22030 43300 22374
rect 43548 22234 43576 22578
rect 43536 22228 43588 22234
rect 43536 22170 43588 22176
rect 43640 22114 43668 22578
rect 43916 22166 43944 22578
rect 44100 22506 44128 22630
rect 44272 22636 44324 22642
rect 44272 22578 44324 22584
rect 44088 22500 44140 22506
rect 44088 22442 44140 22448
rect 44284 22438 44312 22578
rect 44272 22432 44324 22438
rect 44272 22374 44324 22380
rect 44456 22228 44508 22234
rect 44456 22170 44508 22176
rect 43548 22094 43668 22114
rect 43904 22160 43956 22166
rect 43904 22102 43956 22108
rect 43548 22066 43760 22094
rect 43168 22024 43220 22030
rect 43168 21966 43220 21972
rect 43260 22024 43312 22030
rect 43260 21966 43312 21972
rect 42892 21548 42944 21554
rect 42892 21490 42944 21496
rect 42904 19854 42932 21490
rect 42984 20868 43036 20874
rect 42984 20810 43036 20816
rect 42996 20058 43024 20810
rect 43076 20800 43128 20806
rect 43076 20742 43128 20748
rect 43088 20466 43116 20742
rect 43076 20460 43128 20466
rect 43076 20402 43128 20408
rect 42984 20052 43036 20058
rect 42984 19994 43036 20000
rect 42892 19848 42944 19854
rect 42892 19790 42944 19796
rect 43076 19848 43128 19854
rect 43076 19790 43128 19796
rect 42800 17672 42852 17678
rect 42800 17614 42852 17620
rect 41420 17128 41472 17134
rect 41420 17070 41472 17076
rect 40132 4616 40184 4622
rect 40132 4558 40184 4564
rect 40868 4616 40920 4622
rect 40868 4558 40920 4564
rect 39948 4548 40000 4554
rect 39948 4490 40000 4496
rect 39672 3732 39724 3738
rect 39672 3674 39724 3680
rect 39960 3534 39988 4490
rect 40144 3738 40172 4558
rect 40224 4480 40276 4486
rect 40224 4422 40276 4428
rect 40236 4214 40264 4422
rect 40224 4208 40276 4214
rect 40224 4150 40276 4156
rect 40880 3738 40908 4558
rect 41052 4480 41104 4486
rect 41052 4422 41104 4428
rect 40132 3732 40184 3738
rect 40132 3674 40184 3680
rect 40868 3732 40920 3738
rect 40868 3674 40920 3680
rect 41064 3602 41092 4422
rect 41432 4078 41460 17070
rect 42800 17060 42852 17066
rect 42800 17002 42852 17008
rect 42812 15026 42840 17002
rect 42800 15020 42852 15026
rect 42800 14962 42852 14968
rect 42892 4208 42944 4214
rect 42892 4150 42944 4156
rect 41420 4072 41472 4078
rect 41420 4014 41472 4020
rect 41512 4072 41564 4078
rect 41512 4014 41564 4020
rect 41432 3602 41460 4014
rect 41052 3596 41104 3602
rect 41052 3538 41104 3544
rect 41420 3596 41472 3602
rect 41420 3538 41472 3544
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 40592 3528 40644 3534
rect 40592 3470 40644 3476
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 39960 3058 39988 3470
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 40604 2990 40632 3470
rect 40880 3194 40908 3470
rect 40868 3188 40920 3194
rect 40868 3130 40920 3136
rect 39212 2984 39264 2990
rect 39212 2926 39264 2932
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 41432 2922 41460 3538
rect 41524 3058 41552 4014
rect 42800 3460 42852 3466
rect 42800 3402 42852 3408
rect 42432 3392 42484 3398
rect 42432 3334 42484 3340
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 41696 2984 41748 2990
rect 41696 2926 41748 2932
rect 41420 2916 41472 2922
rect 41420 2858 41472 2864
rect 41708 2650 41736 2926
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 41696 2644 41748 2650
rect 41696 2586 41748 2592
rect 39948 2440 40000 2446
rect 39948 2382 40000 2388
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 39396 2372 39448 2378
rect 39396 2314 39448 2320
rect 38476 2304 38528 2310
rect 38476 2246 38528 2252
rect 39408 1170 39436 2314
rect 39316 1142 39436 1170
rect 39316 800 39344 1142
rect 39960 800 39988 2382
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 41248 800 41276 2382
rect 41788 2304 41840 2310
rect 41788 2246 41840 2252
rect 41800 1970 41828 2246
rect 41788 1964 41840 1970
rect 41788 1906 41840 1912
rect 42444 1850 42472 3334
rect 42812 3058 42840 3402
rect 42800 3052 42852 3058
rect 42800 2994 42852 3000
rect 42524 2644 42576 2650
rect 42524 2586 42576 2592
rect 42536 2038 42564 2586
rect 42904 2514 42932 4150
rect 42984 3392 43036 3398
rect 42984 3334 43036 3340
rect 42996 3126 43024 3334
rect 42984 3120 43036 3126
rect 42984 3062 43036 3068
rect 43088 2582 43116 19790
rect 43180 12434 43208 21966
rect 43260 21548 43312 21554
rect 43260 21490 43312 21496
rect 43536 21548 43588 21554
rect 43536 21490 43588 21496
rect 43272 21457 43300 21490
rect 43258 21448 43314 21457
rect 43258 21383 43314 21392
rect 43260 21004 43312 21010
rect 43260 20946 43312 20952
rect 43352 21004 43404 21010
rect 43352 20946 43404 20952
rect 43272 20534 43300 20946
rect 43260 20528 43312 20534
rect 43260 20470 43312 20476
rect 43364 20058 43392 20946
rect 43444 20936 43496 20942
rect 43444 20878 43496 20884
rect 43456 20806 43484 20878
rect 43444 20800 43496 20806
rect 43444 20742 43496 20748
rect 43548 20505 43576 21490
rect 43628 21344 43680 21350
rect 43628 21286 43680 21292
rect 43640 21010 43668 21286
rect 43732 21078 43760 22066
rect 43904 21956 43956 21962
rect 43904 21898 43956 21904
rect 43996 21956 44048 21962
rect 43996 21898 44048 21904
rect 43916 21486 43944 21898
rect 43904 21480 43956 21486
rect 43904 21422 43956 21428
rect 43720 21072 43772 21078
rect 43720 21014 43772 21020
rect 43628 21004 43680 21010
rect 43628 20946 43680 20952
rect 43916 20942 43944 21422
rect 43904 20936 43956 20942
rect 43824 20884 43904 20890
rect 43824 20878 43956 20884
rect 43824 20862 43944 20878
rect 44008 20874 44036 21898
rect 44272 21888 44324 21894
rect 44272 21830 44324 21836
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 43996 20868 44048 20874
rect 43534 20496 43590 20505
rect 43444 20460 43496 20466
rect 43534 20431 43590 20440
rect 43444 20402 43496 20408
rect 43352 20052 43404 20058
rect 43352 19994 43404 20000
rect 43364 19378 43392 19994
rect 43456 19514 43484 20402
rect 43548 19854 43576 20431
rect 43824 19854 43852 20862
rect 43996 20810 44048 20816
rect 43904 20392 43956 20398
rect 43904 20334 43956 20340
rect 43916 19922 43944 20334
rect 43904 19916 43956 19922
rect 43904 19858 43956 19864
rect 43536 19848 43588 19854
rect 43536 19790 43588 19796
rect 43812 19848 43864 19854
rect 43812 19790 43864 19796
rect 43444 19508 43496 19514
rect 43444 19450 43496 19456
rect 43352 19372 43404 19378
rect 43352 19314 43404 19320
rect 43916 18358 43944 19858
rect 44008 19854 44036 20810
rect 44088 20800 44140 20806
rect 44088 20742 44140 20748
rect 43996 19848 44048 19854
rect 43996 19790 44048 19796
rect 43904 18352 43956 18358
rect 43904 18294 43956 18300
rect 43536 18216 43588 18222
rect 43536 18158 43588 18164
rect 43548 17882 43576 18158
rect 43536 17876 43588 17882
rect 43536 17818 43588 17824
rect 43536 17672 43588 17678
rect 43536 17614 43588 17620
rect 43548 15502 43576 17614
rect 43720 17196 43772 17202
rect 43720 17138 43772 17144
rect 43732 16658 43760 17138
rect 43720 16652 43772 16658
rect 43720 16594 43772 16600
rect 43536 15496 43588 15502
rect 43536 15438 43588 15444
rect 43812 15360 43864 15366
rect 43812 15302 43864 15308
rect 43824 15094 43852 15302
rect 43812 15088 43864 15094
rect 43812 15030 43864 15036
rect 43180 12406 43484 12434
rect 43456 6914 43484 12406
rect 43272 6886 43484 6914
rect 43272 4690 43300 6886
rect 44008 6458 44036 19790
rect 44100 19378 44128 20742
rect 44192 19990 44220 21490
rect 44180 19984 44232 19990
rect 44180 19926 44232 19932
rect 44088 19372 44140 19378
rect 44088 19314 44140 19320
rect 44192 17882 44220 19926
rect 44284 19378 44312 21830
rect 44468 21672 44496 22170
rect 44376 21644 44496 21672
rect 45112 22114 45140 24686
rect 45388 24410 45416 24686
rect 45376 24404 45428 24410
rect 45376 24346 45428 24352
rect 45664 24342 45692 26551
rect 45652 24336 45704 24342
rect 45652 24278 45704 24284
rect 45848 24206 45876 28018
rect 45836 24200 45888 24206
rect 45836 24142 45888 24148
rect 45744 23724 45796 23730
rect 45744 23666 45796 23672
rect 45652 23588 45704 23594
rect 45652 23530 45704 23536
rect 45560 23044 45612 23050
rect 45560 22986 45612 22992
rect 45376 22976 45428 22982
rect 45376 22918 45428 22924
rect 45388 22710 45416 22918
rect 45376 22704 45428 22710
rect 45376 22646 45428 22652
rect 45572 22574 45600 22986
rect 45560 22568 45612 22574
rect 45560 22510 45612 22516
rect 45112 22086 45324 22114
rect 44376 21457 44404 21644
rect 45112 21622 45140 22086
rect 45296 22030 45324 22086
rect 45192 22024 45244 22030
rect 45192 21966 45244 21972
rect 45284 22024 45336 22030
rect 45664 21978 45692 23530
rect 45756 23225 45784 23666
rect 45742 23216 45798 23225
rect 45742 23151 45798 23160
rect 45284 21966 45336 21972
rect 45204 21622 45232 21966
rect 45572 21962 45692 21978
rect 45560 21956 45692 21962
rect 45612 21950 45692 21956
rect 45560 21898 45612 21904
rect 45468 21888 45520 21894
rect 45468 21830 45520 21836
rect 45100 21616 45152 21622
rect 44454 21584 44510 21593
rect 45100 21558 45152 21564
rect 45192 21616 45244 21622
rect 45192 21558 45244 21564
rect 44454 21519 44510 21528
rect 44548 21548 44600 21554
rect 44468 21486 44496 21519
rect 44548 21490 44600 21496
rect 44456 21480 44508 21486
rect 44362 21448 44418 21457
rect 44456 21422 44508 21428
rect 44362 21383 44418 21392
rect 44376 20466 44404 21383
rect 44364 20460 44416 20466
rect 44364 20402 44416 20408
rect 44560 19514 44588 21490
rect 45480 21350 45508 21830
rect 45848 21706 45876 24142
rect 45928 23248 45980 23254
rect 45928 23190 45980 23196
rect 45572 21678 45876 21706
rect 45468 21344 45520 21350
rect 45468 21286 45520 21292
rect 45480 20942 45508 21286
rect 45468 20936 45520 20942
rect 45468 20878 45520 20884
rect 44730 20496 44786 20505
rect 44730 20431 44732 20440
rect 44784 20431 44786 20440
rect 44732 20402 44784 20408
rect 44548 19508 44600 19514
rect 44548 19450 44600 19456
rect 44272 19372 44324 19378
rect 44272 19314 44324 19320
rect 45192 18216 45244 18222
rect 45192 18158 45244 18164
rect 44180 17876 44232 17882
rect 44180 17818 44232 17824
rect 44916 17672 44968 17678
rect 44916 17614 44968 17620
rect 44364 17536 44416 17542
rect 44364 17478 44416 17484
rect 44376 17202 44404 17478
rect 44928 17338 44956 17614
rect 45008 17536 45060 17542
rect 45008 17478 45060 17484
rect 45020 17338 45048 17478
rect 44916 17332 44968 17338
rect 44916 17274 44968 17280
rect 45008 17332 45060 17338
rect 45008 17274 45060 17280
rect 44456 17264 44508 17270
rect 44456 17206 44508 17212
rect 44364 17196 44416 17202
rect 44364 17138 44416 17144
rect 44468 16114 44496 17206
rect 44456 16108 44508 16114
rect 44456 16050 44508 16056
rect 45204 6914 45232 18158
rect 45572 16046 45600 21678
rect 45836 20800 45888 20806
rect 45836 20742 45888 20748
rect 45848 20466 45876 20742
rect 45836 20460 45888 20466
rect 45836 20402 45888 20408
rect 45744 20392 45796 20398
rect 45744 20334 45796 20340
rect 45756 19922 45784 20334
rect 45744 19916 45796 19922
rect 45744 19858 45796 19864
rect 45836 18760 45888 18766
rect 45836 18702 45888 18708
rect 45652 18624 45704 18630
rect 45652 18566 45704 18572
rect 45664 17134 45692 18566
rect 45848 18465 45876 18702
rect 45834 18456 45890 18465
rect 45834 18391 45890 18400
rect 45744 17740 45796 17746
rect 45744 17682 45796 17688
rect 45652 17128 45704 17134
rect 45652 17070 45704 17076
rect 45664 16726 45692 17070
rect 45756 16794 45784 17682
rect 45744 16788 45796 16794
rect 45744 16730 45796 16736
rect 45652 16720 45704 16726
rect 45652 16662 45704 16668
rect 45560 16040 45612 16046
rect 45560 15982 45612 15988
rect 45558 15736 45614 15745
rect 45558 15671 45560 15680
rect 45612 15671 45614 15680
rect 45560 15642 45612 15648
rect 45284 14952 45336 14958
rect 45284 14894 45336 14900
rect 45112 6886 45232 6914
rect 43996 6452 44048 6458
rect 43996 6394 44048 6400
rect 43260 4684 43312 4690
rect 43260 4626 43312 4632
rect 43272 4214 43300 4626
rect 44088 4548 44140 4554
rect 44088 4490 44140 4496
rect 43260 4208 43312 4214
rect 43260 4150 43312 4156
rect 44100 3942 44128 4490
rect 44456 4140 44508 4146
rect 44456 4082 44508 4088
rect 44088 3936 44140 3942
rect 44088 3878 44140 3884
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 43076 2576 43128 2582
rect 43076 2518 43128 2524
rect 42892 2508 42944 2514
rect 42892 2450 42944 2456
rect 42524 2032 42576 2038
rect 42524 1974 42576 1980
rect 42444 1822 42564 1850
rect 42536 800 42564 1822
rect 43180 800 43208 2926
rect 44468 2650 44496 4082
rect 45112 3194 45140 6886
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 45100 3188 45152 3194
rect 45100 3130 45152 3136
rect 45204 3058 45232 3470
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45296 2938 45324 14894
rect 45940 12238 45968 23190
rect 46032 21418 46060 31062
rect 46112 30660 46164 30666
rect 46112 30602 46164 30608
rect 46124 21690 46152 30602
rect 46202 28656 46258 28665
rect 46202 28591 46258 28600
rect 46216 27674 46244 28591
rect 46204 27668 46256 27674
rect 46204 27610 46256 27616
rect 46388 26376 46440 26382
rect 46388 26318 46440 26324
rect 46296 25696 46348 25702
rect 46296 25638 46348 25644
rect 46308 25362 46336 25638
rect 46296 25356 46348 25362
rect 46296 25298 46348 25304
rect 46296 24200 46348 24206
rect 46296 24142 46348 24148
rect 46204 23656 46256 23662
rect 46204 23598 46256 23604
rect 46216 22545 46244 23598
rect 46308 22982 46336 24142
rect 46400 23254 46428 26318
rect 46492 24274 46520 31062
rect 46676 26234 46704 31311
rect 47320 30666 47348 33458
rect 47308 30660 47360 30666
rect 47308 30602 47360 30608
rect 46848 30184 46900 30190
rect 46848 30126 46900 30132
rect 46860 30025 46888 30126
rect 46846 30016 46902 30025
rect 46846 29951 46902 29960
rect 47216 29708 47268 29714
rect 47216 29650 47268 29656
rect 46940 28552 46992 28558
rect 46940 28494 46992 28500
rect 46952 27606 46980 28494
rect 46940 27600 46992 27606
rect 46940 27542 46992 27548
rect 46584 26206 46704 26234
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46388 23248 46440 23254
rect 46388 23190 46440 23196
rect 46296 22976 46348 22982
rect 46296 22918 46348 22924
rect 46202 22536 46258 22545
rect 46202 22471 46258 22480
rect 46202 21856 46258 21865
rect 46202 21791 46258 21800
rect 46112 21684 46164 21690
rect 46112 21626 46164 21632
rect 46216 21554 46244 21791
rect 46204 21548 46256 21554
rect 46204 21490 46256 21496
rect 46480 21480 46532 21486
rect 46480 21422 46532 21428
rect 46020 21412 46072 21418
rect 46020 21354 46072 21360
rect 46492 21146 46520 21422
rect 46480 21140 46532 21146
rect 46480 21082 46532 21088
rect 46480 20868 46532 20874
rect 46480 20810 46532 20816
rect 46492 20602 46520 20810
rect 46480 20596 46532 20602
rect 46480 20538 46532 20544
rect 46584 19786 46612 26206
rect 46754 25936 46810 25945
rect 46754 25871 46810 25880
rect 46768 24750 46796 25871
rect 46756 24744 46808 24750
rect 46756 24686 46808 24692
rect 46848 24676 46900 24682
rect 46848 24618 46900 24624
rect 46860 23905 46888 24618
rect 46846 23896 46902 23905
rect 46846 23831 46902 23840
rect 47032 23724 47084 23730
rect 47032 23666 47084 23672
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 46952 22710 46980 23462
rect 46940 22704 46992 22710
rect 46940 22646 46992 22652
rect 46952 21078 46980 22646
rect 47044 21554 47072 23666
rect 47228 22658 47256 29650
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47320 29345 47348 29582
rect 47306 29336 47362 29345
rect 47306 29271 47362 29280
rect 47412 26234 47440 35866
rect 47136 22642 47256 22658
rect 47124 22636 47256 22642
rect 47176 22630 47256 22636
rect 47320 26206 47440 26234
rect 47124 22578 47176 22584
rect 47216 22568 47268 22574
rect 47216 22510 47268 22516
rect 47228 22094 47256 22510
rect 47136 22066 47256 22094
rect 47136 21962 47164 22066
rect 47124 21956 47176 21962
rect 47124 21898 47176 21904
rect 47032 21548 47084 21554
rect 47032 21490 47084 21496
rect 46940 21072 46992 21078
rect 46940 21014 46992 21020
rect 46940 19916 46992 19922
rect 46940 19858 46992 19864
rect 46572 19780 46624 19786
rect 46572 19722 46624 19728
rect 46020 19508 46072 19514
rect 46020 19450 46072 19456
rect 46032 18290 46060 19450
rect 46388 19440 46440 19446
rect 46388 19382 46440 19388
rect 46400 18290 46428 19382
rect 46756 19372 46808 19378
rect 46756 19314 46808 19320
rect 46768 18290 46796 19314
rect 46020 18284 46072 18290
rect 46020 18226 46072 18232
rect 46388 18284 46440 18290
rect 46388 18226 46440 18232
rect 46756 18284 46808 18290
rect 46756 18226 46808 18232
rect 46296 18080 46348 18086
rect 46296 18022 46348 18028
rect 46308 17270 46336 18022
rect 46400 17814 46428 18226
rect 46768 18154 46796 18226
rect 46952 18170 46980 19858
rect 47044 19394 47072 21490
rect 47136 19922 47164 21898
rect 47216 21140 47268 21146
rect 47216 21082 47268 21088
rect 47124 19916 47176 19922
rect 47124 19858 47176 19864
rect 47044 19366 47164 19394
rect 47032 19236 47084 19242
rect 47032 19178 47084 19184
rect 47044 18290 47072 19178
rect 47032 18284 47084 18290
rect 47032 18226 47084 18232
rect 46756 18148 46808 18154
rect 46952 18142 47072 18170
rect 46756 18090 46808 18096
rect 46388 17808 46440 17814
rect 46388 17750 46440 17756
rect 46296 17264 46348 17270
rect 46296 17206 46348 17212
rect 46664 17196 46716 17202
rect 46664 17138 46716 17144
rect 46676 17082 46704 17138
rect 46584 17054 46704 17082
rect 46584 16454 46612 17054
rect 46572 16448 46624 16454
rect 46572 16390 46624 16396
rect 46112 16040 46164 16046
rect 46112 15982 46164 15988
rect 45928 12232 45980 12238
rect 45928 12174 45980 12180
rect 45652 7948 45704 7954
rect 45652 7890 45704 7896
rect 45664 4078 45692 7890
rect 46124 6914 46152 15982
rect 46480 12096 46532 12102
rect 46480 12038 46532 12044
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46492 11218 46520 12038
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46480 11212 46532 11218
rect 46480 11154 46532 11160
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46584 7818 46612 16390
rect 46204 7812 46256 7818
rect 46204 7754 46256 7760
rect 46572 7812 46624 7818
rect 46572 7754 46624 7760
rect 46216 7410 46244 7754
rect 46204 7404 46256 7410
rect 46204 7346 46256 7352
rect 46216 7290 46244 7346
rect 46216 7262 46336 7290
rect 46124 6886 46244 6914
rect 45652 4072 45704 4078
rect 45652 4014 45704 4020
rect 46216 3505 46244 6886
rect 46308 4758 46336 7262
rect 46296 4752 46348 4758
rect 46296 4694 46348 4700
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 46388 4208 46440 4214
rect 46388 4150 46440 4156
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3602 46336 3878
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46202 3496 46258 3505
rect 46202 3431 46258 3440
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45112 2910 45324 2938
rect 44456 2644 44508 2650
rect 44456 2586 44508 2592
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 45112 800 45140 2910
rect 46400 800 46428 4150
rect 46492 3602 46520 4422
rect 46664 4208 46716 4214
rect 46664 4150 46716 4156
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 20180 734 20392 762
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46676 82 46704 4150
rect 46768 2514 46796 18090
rect 46848 17740 46900 17746
rect 46848 17682 46900 17688
rect 46860 15026 46888 17682
rect 46940 17604 46992 17610
rect 46940 17546 46992 17552
rect 46952 16250 46980 17546
rect 47044 17134 47072 18142
rect 47032 17128 47084 17134
rect 47032 17070 47084 17076
rect 46940 16244 46992 16250
rect 46940 16186 46992 16192
rect 47136 16114 47164 19366
rect 47124 16108 47176 16114
rect 47124 16050 47176 16056
rect 47124 15972 47176 15978
rect 47124 15914 47176 15920
rect 46848 15020 46900 15026
rect 46848 14962 46900 14968
rect 47136 14414 47164 15914
rect 47124 14408 47176 14414
rect 47124 14350 47176 14356
rect 46848 8492 46900 8498
rect 46848 8434 46900 8440
rect 46860 8378 46888 8434
rect 46860 8350 46980 8378
rect 46848 8288 46900 8294
rect 46846 8256 46848 8265
rect 46900 8256 46902 8265
rect 46846 8191 46902 8200
rect 46952 8106 46980 8350
rect 47124 8288 47176 8294
rect 47124 8230 47176 8236
rect 46860 8078 46980 8106
rect 46860 6905 46888 8078
rect 47136 7954 47164 8230
rect 47124 7948 47176 7954
rect 47124 7890 47176 7896
rect 46846 6896 46902 6905
rect 46846 6831 46902 6840
rect 47228 6798 47256 21082
rect 47320 19514 47348 26206
rect 47504 23798 47532 37810
rect 47596 24818 47624 42162
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 40730 47716 41618
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47676 38956 47728 38962
rect 47676 38898 47728 38904
rect 47688 38865 47716 38898
rect 47860 38888 47912 38894
rect 47674 38856 47730 38865
rect 47860 38830 47912 38836
rect 47674 38791 47730 38800
rect 47676 37664 47728 37670
rect 47676 37606 47728 37612
rect 47688 37194 47716 37606
rect 47676 37188 47728 37194
rect 47676 37130 47728 37136
rect 47872 35894 47900 38830
rect 47872 35866 47992 35894
rect 47860 34944 47912 34950
rect 47860 34886 47912 34892
rect 47768 34604 47820 34610
rect 47768 34546 47820 34552
rect 47676 34060 47728 34066
rect 47676 34002 47728 34008
rect 47688 30802 47716 34002
rect 47780 33658 47808 34546
rect 47768 33652 47820 33658
rect 47768 33594 47820 33600
rect 47872 33318 47900 34886
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 47964 31090 47992 35866
rect 48056 32026 48084 47126
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48148 37330 48176 38111
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 48136 35692 48188 35698
rect 48136 35634 48188 35640
rect 48148 34785 48176 35634
rect 48228 35080 48280 35086
rect 48228 35022 48280 35028
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48240 34105 48268 35022
rect 48226 34096 48282 34105
rect 48226 34031 48282 34040
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48044 32020 48096 32026
rect 48044 31962 48096 31968
rect 48148 31890 48176 32671
rect 48136 31884 48188 31890
rect 48136 31826 48188 31832
rect 47780 31062 47992 31090
rect 47676 30796 47728 30802
rect 47676 30738 47728 30744
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27538 47716 27814
rect 47676 27532 47728 27538
rect 47676 27474 47728 27480
rect 47676 25220 47728 25226
rect 47676 25162 47728 25168
rect 47688 24818 47716 25162
rect 47584 24812 47636 24818
rect 47584 24754 47636 24760
rect 47676 24812 47728 24818
rect 47676 24754 47728 24760
rect 47492 23792 47544 23798
rect 47492 23734 47544 23740
rect 47596 22794 47624 24754
rect 47780 24070 47808 31062
rect 48044 30796 48096 30802
rect 48044 30738 48096 30744
rect 47952 30660 48004 30666
rect 47952 30602 48004 30608
rect 47768 24064 47820 24070
rect 47768 24006 47820 24012
rect 47676 23520 47728 23526
rect 47676 23462 47728 23468
rect 47688 23186 47716 23462
rect 47676 23180 47728 23186
rect 47676 23122 47728 23128
rect 47768 23044 47820 23050
rect 47768 22986 47820 22992
rect 47504 22766 47624 22794
rect 47676 22772 47728 22778
rect 47504 22506 47532 22766
rect 47676 22714 47728 22720
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47492 22500 47544 22506
rect 47492 22442 47544 22448
rect 47400 22092 47452 22098
rect 47400 22034 47452 22040
rect 47412 20466 47440 22034
rect 47400 20460 47452 20466
rect 47400 20402 47452 20408
rect 47308 19508 47360 19514
rect 47308 19450 47360 19456
rect 47412 19446 47440 20402
rect 47400 19440 47452 19446
rect 47400 19382 47452 19388
rect 47504 18306 47532 22442
rect 47596 21706 47624 22578
rect 47688 22098 47716 22714
rect 47676 22092 47728 22098
rect 47676 22034 47728 22040
rect 47596 21678 47716 21706
rect 47780 21690 47808 22986
rect 47860 22636 47912 22642
rect 47860 22578 47912 22584
rect 47688 21622 47716 21678
rect 47768 21684 47820 21690
rect 47768 21626 47820 21632
rect 47676 21616 47728 21622
rect 47676 21558 47728 21564
rect 47584 21548 47636 21554
rect 47584 21490 47636 21496
rect 47596 21078 47624 21490
rect 47584 21072 47636 21078
rect 47584 21014 47636 21020
rect 47688 20262 47716 21558
rect 47872 21486 47900 22578
rect 47860 21480 47912 21486
rect 47860 21422 47912 21428
rect 47872 21146 47900 21422
rect 47860 21140 47912 21146
rect 47860 21082 47912 21088
rect 47860 21004 47912 21010
rect 47860 20946 47912 20952
rect 47676 20256 47728 20262
rect 47676 20198 47728 20204
rect 47872 20058 47900 20946
rect 47860 20052 47912 20058
rect 47860 19994 47912 20000
rect 47768 19168 47820 19174
rect 47768 19110 47820 19116
rect 47780 18834 47808 19110
rect 47768 18828 47820 18834
rect 47768 18770 47820 18776
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47688 18426 47716 18634
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47504 18290 47624 18306
rect 47504 18284 47636 18290
rect 47504 18278 47584 18284
rect 47584 18226 47636 18232
rect 47492 16652 47544 16658
rect 47492 16594 47544 16600
rect 47400 16108 47452 16114
rect 47400 16050 47452 16056
rect 47308 14272 47360 14278
rect 47308 14214 47360 14220
rect 47320 13258 47348 14214
rect 47308 13252 47360 13258
rect 47308 13194 47360 13200
rect 47412 10674 47440 16050
rect 47504 15706 47532 16594
rect 47492 15700 47544 15706
rect 47492 15642 47544 15648
rect 47596 12434 47624 18226
rect 47860 18216 47912 18222
rect 47860 18158 47912 18164
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47688 16250 47716 16458
rect 47676 16244 47728 16250
rect 47676 16186 47728 16192
rect 47768 13728 47820 13734
rect 47768 13670 47820 13676
rect 47780 13394 47808 13670
rect 47768 13388 47820 13394
rect 47768 13330 47820 13336
rect 47504 12406 47624 12434
rect 47400 10668 47452 10674
rect 47400 10610 47452 10616
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47320 6866 47348 7511
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 47216 6792 47268 6798
rect 47216 6734 47268 6740
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46860 4185 46888 4558
rect 46846 4176 46902 4185
rect 46846 4111 46902 4120
rect 47412 3466 47440 10610
rect 47504 4690 47532 12406
rect 47676 10464 47728 10470
rect 47676 10406 47728 10412
rect 47688 10130 47716 10406
rect 47676 10124 47728 10130
rect 47676 10066 47728 10072
rect 47872 10010 47900 18158
rect 47688 9982 47900 10010
rect 47584 7812 47636 7818
rect 47584 7754 47636 7760
rect 47596 7546 47624 7754
rect 47584 7540 47636 7546
rect 47584 7482 47636 7488
rect 47492 4684 47544 4690
rect 47492 4626 47544 4632
rect 47400 3460 47452 3466
rect 47400 3402 47452 3408
rect 47688 3194 47716 9982
rect 47858 9616 47914 9625
rect 47858 9551 47860 9560
rect 47912 9551 47914 9560
rect 47860 9522 47912 9528
rect 47964 9450 47992 30602
rect 48056 22234 48084 30738
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48226 25256 48282 25265
rect 48136 25220 48188 25226
rect 48226 25191 48282 25200
rect 48136 25162 48188 25168
rect 48148 24585 48176 25162
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48240 23186 48268 25191
rect 48228 23180 48280 23186
rect 48228 23122 48280 23128
rect 48136 22432 48188 22438
rect 48136 22374 48188 22380
rect 48044 22228 48096 22234
rect 48044 22170 48096 22176
rect 48148 22137 48176 22374
rect 48134 22128 48190 22137
rect 48134 22063 48190 22072
rect 48044 22024 48096 22030
rect 48044 21966 48096 21972
rect 48056 20602 48084 21966
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48044 20596 48096 20602
rect 48044 20538 48096 20544
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 48148 17105 48176 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 48148 16425 48176 16458
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 48148 12345 48176 13194
rect 48134 12336 48190 12345
rect 48134 12271 48190 12280
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 47952 9444 48004 9450
rect 47952 9386 48004 9392
rect 47766 8936 47822 8945
rect 47766 8871 47768 8880
rect 47820 8871 47822 8880
rect 47768 8842 47820 8848
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 47964 6225 47992 6258
rect 47950 6216 48006 6225
rect 47950 6151 48006 6160
rect 47952 5228 48004 5234
rect 47952 5170 48004 5176
rect 47860 3936 47912 3942
rect 47860 3878 47912 3884
rect 47872 3670 47900 3878
rect 47860 3664 47912 3670
rect 47860 3606 47912 3612
rect 47964 3505 47992 5170
rect 47950 3496 48006 3505
rect 47950 3431 48006 3440
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 47676 3188 47728 3194
rect 47676 3130 47728 3136
rect 48320 3052 48372 3058
rect 48320 2994 48372 3000
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 46756 2508 46808 2514
rect 46756 2450 46808 2456
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 46756 2372 46808 2378
rect 46756 2314 46808 2320
rect 46768 1465 46796 2314
rect 46754 1456 46810 1465
rect 46754 1391 46810 1400
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 46754 96 46810 105
rect 46676 54 46754 82
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48056 785 48084 2382
rect 48332 800 48360 2994
rect 48976 800 49004 3402
rect 48042 776 48098 785
rect 48042 711 48098 720
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1858 47640 1914 47696
rect 3514 46960 3570 47016
rect 1398 42880 1454 42936
rect 1398 33360 1454 33416
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1582 35400 1638 35456
rect 1582 32680 1638 32736
rect 2778 46280 2834 46336
rect 1398 17720 1454 17776
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 1858 23160 1914 23216
rect 1858 16360 1914 16416
rect 1398 12280 1454 12336
rect 2778 36760 2834 36816
rect 2778 32000 2834 32056
rect 3422 44920 3478 44976
rect 3330 31320 3386 31376
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3698 43560 3754 43616
rect 3606 28600 3662 28656
rect 3882 39480 3938 39536
rect 2962 19760 3018 19816
rect 2226 19080 2282 19136
rect 3422 18420 3478 18456
rect 3422 18400 3424 18420
rect 3424 18400 3476 18420
rect 3476 18400 3478 18420
rect 3422 17040 3478 17096
rect 2778 15000 2834 15056
rect 3422 13640 3478 13696
rect 2962 10240 3018 10296
rect 3330 6860 3386 6896
rect 3330 6840 3332 6860
rect 3332 6840 3384 6860
rect 3384 6840 3386 6860
rect 3514 7520 3570 7576
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3514 3440 3570 3496
rect 3422 1400 3478 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 20074 24112 20130 24168
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19522 23704 19578 23760
rect 19338 23568 19394 23624
rect 17498 3440 17554 3496
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19890 22092 19946 22128
rect 19890 22072 19892 22092
rect 19892 22072 19944 22092
rect 19944 22072 19946 22092
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 20074 21392 20130 21448
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19430 19760 19486 19816
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19338 18128 19394 18184
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19982 14320 20038 14376
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20810 23704 20866 23760
rect 20902 21956 20958 21992
rect 20902 21936 20904 21956
rect 20904 21936 20956 21956
rect 20956 21936 20958 21956
rect 20718 20868 20774 20904
rect 20718 20848 20720 20868
rect 20720 20848 20772 20868
rect 20772 20848 20774 20868
rect 21914 29552 21970 29608
rect 21270 20848 21326 20904
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 2870 720 2926 776
rect 21730 22072 21786 22128
rect 23202 29688 23258 29744
rect 22466 21936 22522 21992
rect 24674 35128 24730 35184
rect 24582 35012 24638 35048
rect 24582 34992 24584 35012
rect 24584 34992 24636 35012
rect 24636 34992 24638 35012
rect 24582 30232 24638 30288
rect 23294 23568 23350 23624
rect 25134 31592 25190 31648
rect 24766 29572 24822 29608
rect 24766 29552 24768 29572
rect 24768 29552 24820 29572
rect 24820 29552 24822 29572
rect 26698 29280 26754 29336
rect 26974 29144 27030 29200
rect 27802 31592 27858 31648
rect 27434 29572 27490 29608
rect 27434 29552 27436 29572
rect 27436 29552 27488 29572
rect 27488 29552 27490 29572
rect 27710 29300 27766 29336
rect 27710 29280 27712 29300
rect 27712 29280 27764 29300
rect 27764 29280 27766 29300
rect 27802 29164 27858 29200
rect 27802 29144 27804 29164
rect 27804 29144 27856 29164
rect 27856 29144 27858 29164
rect 28078 35128 28134 35184
rect 28170 30252 28226 30288
rect 28170 30232 28172 30252
rect 28172 30232 28224 30252
rect 28224 30232 28226 30252
rect 27986 29708 28042 29744
rect 27986 29688 27988 29708
rect 27988 29688 28040 29708
rect 28040 29688 28042 29708
rect 28722 34992 28778 35048
rect 28446 30232 28502 30288
rect 28354 21412 28410 21448
rect 28354 21392 28356 21412
rect 28356 21392 28408 21412
rect 28408 21392 28410 21412
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 29274 30268 29276 30288
rect 29276 30268 29328 30288
rect 29328 30268 29330 30288
rect 29274 30232 29330 30268
rect 29458 31592 29514 31648
rect 29734 29552 29790 29608
rect 30010 29008 30066 29064
rect 29734 21392 29790 21448
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 32310 29552 32366 29608
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 33874 29588 33876 29608
rect 33876 29588 33928 29608
rect 33928 29588 33930 29608
rect 33874 29552 33930 29588
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34610 29008 34666 29064
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 40038 22072 40094 22128
rect 42706 21528 42762 21584
rect 46846 47640 46902 47696
rect 46386 46960 46442 47016
rect 46570 39480 46626 39536
rect 47950 46280 48006 46336
rect 46846 33360 46902 33416
rect 46846 32000 46902 32056
rect 46662 31320 46718 31376
rect 45650 26560 45706 26616
rect 43258 21392 43314 21448
rect 43534 20440 43590 20496
rect 45742 23160 45798 23216
rect 44454 21528 44510 21584
rect 44362 21392 44418 21448
rect 44730 20460 44786 20496
rect 44730 20440 44732 20460
rect 44732 20440 44784 20460
rect 44784 20440 44786 20460
rect 45834 18400 45890 18456
rect 45558 15700 45614 15736
rect 45558 15680 45560 15700
rect 45560 15680 45612 15700
rect 45612 15680 45614 15700
rect 46202 28600 46258 28656
rect 46846 29960 46902 30016
rect 46202 22480 46258 22536
rect 46202 21800 46258 21856
rect 46754 25880 46810 25936
rect 46846 23840 46902 23896
rect 47306 29280 47362 29336
rect 46202 3440 46258 3496
rect 46846 8236 46848 8256
rect 46848 8236 46900 8256
rect 46900 8236 46902 8256
rect 46846 8200 46902 8236
rect 46846 6840 46902 6896
rect 47950 40840 48006 40896
rect 47674 38800 47730 38856
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48226 34040 48282 34096
rect 48134 32680 48190 32736
rect 47306 7520 47362 7576
rect 46846 4120 46902 4176
rect 47858 9580 47914 9616
rect 47858 9560 47860 9580
rect 47860 9560 47912 9580
rect 47912 9560 47914 9580
rect 48134 27920 48190 27976
rect 48226 25200 48282 25256
rect 48134 24520 48190 24576
rect 48134 22072 48190 22128
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12280 48190 12336
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 47766 8900 47822 8936
rect 47766 8880 47768 8900
rect 47768 8880 47820 8900
rect 47820 8880 47822 8900
rect 47950 6160 48006 6216
rect 47950 3440 48006 3496
rect 46754 1400 46810 1456
rect 46754 40 46810 96
rect 48042 720 48098 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1853 47698 1919 47701
rect 0 47696 1919 47698
rect 0 47640 1858 47696
rect 1914 47640 1919 47696
rect 0 47638 1919 47640
rect 0 47548 800 47638
rect 1853 47635 1919 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3509 47018 3575 47021
rect 0 47016 3575 47018
rect 0 46960 3514 47016
rect 3570 46960 3575 47016
rect 0 46958 3575 46960
rect 0 46868 800 46958
rect 3509 46955 3575 46958
rect 46381 47018 46447 47021
rect 49200 47018 50000 47108
rect 46381 47016 50000 47018
rect 46381 46960 46386 47016
rect 46442 46960 50000 47016
rect 46381 46958 50000 46960
rect 46381 46955 46447 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3417 44978 3483 44981
rect 0 44976 3483 44978
rect 0 44920 3422 44976
rect 3478 44920 3483 44976
rect 0 44918 3483 44920
rect 0 44828 800 44918
rect 3417 44915 3483 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3693 43618 3759 43621
rect 0 43616 3759 43618
rect 0 43560 3698 43616
rect 3754 43560 3759 43616
rect 0 43558 3759 43560
rect 0 43468 800 43558
rect 3693 43555 3759 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3877 39538 3943 39541
rect 0 39536 3943 39538
rect 0 39480 3882 39536
rect 3938 39480 3943 39536
rect 0 39478 3943 39480
rect 0 39388 800 39478
rect 3877 39475 3943 39478
rect 46565 39538 46631 39541
rect 49200 39538 50000 39628
rect 46565 39536 50000 39538
rect 46565 39480 46570 39536
rect 46626 39480 50000 39536
rect 46565 39478 50000 39480
rect 46565 39475 46631 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47669 38858 47735 38861
rect 49200 38858 50000 38948
rect 47669 38856 50000 38858
rect 47669 38800 47674 38856
rect 47730 38800 50000 38856
rect 47669 38798 50000 38800
rect 47669 38795 47735 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 24669 35186 24735 35189
rect 28073 35186 28139 35189
rect 24669 35184 28139 35186
rect 24669 35128 24674 35184
rect 24730 35128 28078 35184
rect 28134 35128 28139 35184
rect 24669 35126 28139 35128
rect 24669 35123 24735 35126
rect 28073 35123 28139 35126
rect 24577 35050 24643 35053
rect 28717 35050 28783 35053
rect 24577 35048 28783 35050
rect 24577 34992 24582 35048
rect 24638 34992 28722 35048
rect 28778 34992 28783 35048
rect 24577 34990 28783 34992
rect 24577 34987 24643 34990
rect 28717 34987 28783 34990
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48221 34098 48287 34101
rect 49200 34098 50000 34188
rect 48221 34096 50000 34098
rect 48221 34040 48226 34096
rect 48282 34040 50000 34096
rect 48221 34038 50000 34040
rect 48221 34035 48287 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 46841 33418 46907 33421
rect 49200 33418 50000 33508
rect 46841 33416 50000 33418
rect 46841 33360 46846 33416
rect 46902 33360 50000 33416
rect 46841 33358 50000 33360
rect 46841 33355 46907 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 2773 32058 2839 32061
rect 0 32056 2839 32058
rect 0 32000 2778 32056
rect 2834 32000 2839 32056
rect 0 31998 2839 32000
rect 0 31908 800 31998
rect 2773 31995 2839 31998
rect 46841 32058 46907 32061
rect 49200 32058 50000 32148
rect 46841 32056 50000 32058
rect 46841 32000 46846 32056
rect 46902 32000 50000 32056
rect 46841 31998 50000 32000
rect 46841 31995 46907 31998
rect 49200 31908 50000 31998
rect 25129 31650 25195 31653
rect 27797 31650 27863 31653
rect 29453 31650 29519 31653
rect 25129 31648 29519 31650
rect 25129 31592 25134 31648
rect 25190 31592 27802 31648
rect 27858 31592 29458 31648
rect 29514 31592 29519 31648
rect 25129 31590 29519 31592
rect 25129 31587 25195 31590
rect 27797 31587 27863 31590
rect 29453 31587 29519 31590
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3325 31378 3391 31381
rect 0 31376 3391 31378
rect 0 31320 3330 31376
rect 3386 31320 3391 31376
rect 0 31318 3391 31320
rect 0 31228 800 31318
rect 3325 31315 3391 31318
rect 46657 31378 46723 31381
rect 49200 31378 50000 31468
rect 46657 31376 50000 31378
rect 46657 31320 46662 31376
rect 46718 31320 50000 31376
rect 46657 31318 50000 31320
rect 46657 31315 46723 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 24577 30290 24643 30293
rect 28165 30290 28231 30293
rect 24577 30288 28231 30290
rect 24577 30232 24582 30288
rect 24638 30232 28170 30288
rect 28226 30232 28231 30288
rect 24577 30230 28231 30232
rect 24577 30227 24643 30230
rect 28165 30227 28231 30230
rect 28441 30290 28507 30293
rect 29269 30290 29335 30293
rect 28441 30288 29335 30290
rect 28441 30232 28446 30288
rect 28502 30232 29274 30288
rect 29330 30232 29335 30288
rect 28441 30230 29335 30232
rect 28441 30227 28507 30230
rect 29269 30227 29335 30230
rect 0 29868 800 30108
rect 46841 30018 46907 30021
rect 49200 30018 50000 30108
rect 46841 30016 50000 30018
rect 46841 29960 46846 30016
rect 46902 29960 50000 30016
rect 46841 29958 50000 29960
rect 46841 29955 46907 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 23197 29746 23263 29749
rect 27981 29746 28047 29749
rect 23197 29744 28047 29746
rect 23197 29688 23202 29744
rect 23258 29688 27986 29744
rect 28042 29688 28047 29744
rect 23197 29686 28047 29688
rect 23197 29683 23263 29686
rect 27981 29683 28047 29686
rect 21909 29610 21975 29613
rect 24761 29610 24827 29613
rect 27429 29610 27495 29613
rect 21909 29608 27495 29610
rect 21909 29552 21914 29608
rect 21970 29552 24766 29608
rect 24822 29552 27434 29608
rect 27490 29552 27495 29608
rect 21909 29550 27495 29552
rect 21909 29547 21975 29550
rect 24761 29547 24827 29550
rect 27429 29547 27495 29550
rect 29729 29610 29795 29613
rect 32305 29610 32371 29613
rect 33869 29610 33935 29613
rect 29729 29608 33935 29610
rect 29729 29552 29734 29608
rect 29790 29552 32310 29608
rect 32366 29552 33874 29608
rect 33930 29552 33935 29608
rect 29729 29550 33935 29552
rect 29729 29547 29795 29550
rect 32305 29547 32371 29550
rect 33869 29547 33935 29550
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 26693 29338 26759 29341
rect 27705 29338 27771 29341
rect 26693 29336 27771 29338
rect 26693 29280 26698 29336
rect 26754 29280 27710 29336
rect 27766 29280 27771 29336
rect 26693 29278 27771 29280
rect 26693 29275 26759 29278
rect 27705 29275 27771 29278
rect 47301 29338 47367 29341
rect 49200 29338 50000 29428
rect 47301 29336 50000 29338
rect 47301 29280 47306 29336
rect 47362 29280 50000 29336
rect 47301 29278 50000 29280
rect 47301 29275 47367 29278
rect 26969 29202 27035 29205
rect 27797 29202 27863 29205
rect 26969 29200 27863 29202
rect 26969 29144 26974 29200
rect 27030 29144 27802 29200
rect 27858 29144 27863 29200
rect 49200 29188 50000 29278
rect 26969 29142 27863 29144
rect 26969 29139 27035 29142
rect 27797 29139 27863 29142
rect 30005 29066 30071 29069
rect 34605 29066 34671 29069
rect 30005 29064 34671 29066
rect 30005 29008 30010 29064
rect 30066 29008 34610 29064
rect 34666 29008 34671 29064
rect 30005 29006 34671 29008
rect 30005 29003 30071 29006
rect 34605 29003 34671 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3601 28658 3667 28661
rect 0 28656 3667 28658
rect 0 28600 3606 28656
rect 3662 28600 3667 28656
rect 0 28598 3667 28600
rect 0 28508 800 28598
rect 3601 28595 3667 28598
rect 46197 28658 46263 28661
rect 49200 28658 50000 28748
rect 46197 28656 50000 28658
rect 46197 28600 46202 28656
rect 46258 28600 50000 28656
rect 46197 28598 50000 28600
rect 46197 28595 46263 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 45645 26618 45711 26621
rect 49200 26618 50000 26708
rect 45645 26616 50000 26618
rect 45645 26560 45650 26616
rect 45706 26560 50000 26616
rect 45645 26558 50000 26560
rect 45645 26555 45711 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 46749 25938 46815 25941
rect 49200 25938 50000 26028
rect 46749 25936 50000 25938
rect 46749 25880 46754 25936
rect 46810 25880 50000 25936
rect 46749 25878 50000 25880
rect 46749 25875 46815 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 48221 25258 48287 25261
rect 49200 25258 50000 25348
rect 48221 25256 50000 25258
rect 48221 25200 48226 25256
rect 48282 25200 50000 25256
rect 48221 25198 50000 25200
rect 48221 25195 48287 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 20069 24172 20135 24173
rect 20069 24168 20116 24172
rect 20180 24170 20186 24172
rect 20069 24112 20074 24168
rect 20069 24108 20116 24112
rect 20180 24110 20226 24170
rect 20180 24108 20186 24110
rect 20069 24107 20135 24108
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46841 23898 46907 23901
rect 49200 23898 50000 23988
rect 46841 23896 50000 23898
rect 46841 23840 46846 23896
rect 46902 23840 50000 23896
rect 46841 23838 50000 23840
rect 46841 23835 46907 23838
rect 19517 23762 19583 23765
rect 20805 23762 20871 23765
rect 19517 23760 20871 23762
rect 19517 23704 19522 23760
rect 19578 23704 20810 23760
rect 20866 23704 20871 23760
rect 49200 23748 50000 23838
rect 19517 23702 20871 23704
rect 19517 23699 19583 23702
rect 20805 23699 20871 23702
rect 19333 23626 19399 23629
rect 23289 23626 23355 23629
rect 19333 23624 23355 23626
rect 19333 23568 19338 23624
rect 19394 23568 23294 23624
rect 23350 23568 23355 23624
rect 19333 23566 23355 23568
rect 19333 23563 19399 23566
rect 23289 23563 23355 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 45737 23218 45803 23221
rect 49200 23218 50000 23308
rect 45737 23216 50000 23218
rect 45737 23160 45742 23216
rect 45798 23160 50000 23216
rect 45737 23158 50000 23160
rect 45737 23155 45803 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46197 22538 46263 22541
rect 49200 22538 50000 22628
rect 46197 22536 50000 22538
rect 46197 22480 46202 22536
rect 46258 22480 50000 22536
rect 46197 22478 50000 22480
rect 46197 22475 46263 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19374 22068 19380 22132
rect 19444 22130 19450 22132
rect 19885 22130 19951 22133
rect 21725 22130 21791 22133
rect 19444 22128 21791 22130
rect 19444 22072 19890 22128
rect 19946 22072 21730 22128
rect 21786 22072 21791 22128
rect 19444 22070 21791 22072
rect 19444 22068 19450 22070
rect 19885 22067 19951 22070
rect 21725 22067 21791 22070
rect 40033 22130 40099 22133
rect 48129 22130 48195 22133
rect 40033 22128 48195 22130
rect 40033 22072 40038 22128
rect 40094 22072 48134 22128
rect 48190 22072 48195 22128
rect 40033 22070 48195 22072
rect 40033 22067 40099 22070
rect 48129 22067 48195 22070
rect 20897 21994 20963 21997
rect 22461 21994 22527 21997
rect 20897 21992 22527 21994
rect 0 21708 800 21948
rect 20897 21936 20902 21992
rect 20958 21936 22466 21992
rect 22522 21936 22527 21992
rect 20897 21934 22527 21936
rect 20897 21931 20963 21934
rect 22461 21931 22527 21934
rect 46197 21858 46263 21861
rect 49200 21858 50000 21948
rect 46197 21856 50000 21858
rect 46197 21800 46202 21856
rect 46258 21800 50000 21856
rect 46197 21798 50000 21800
rect 46197 21795 46263 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 42701 21586 42767 21589
rect 44449 21586 44515 21589
rect 42701 21584 44515 21586
rect 42701 21528 42706 21584
rect 42762 21528 44454 21584
rect 44510 21528 44515 21584
rect 42701 21526 44515 21528
rect 42701 21523 42767 21526
rect 44449 21523 44515 21526
rect 20069 21452 20135 21453
rect 20069 21450 20116 21452
rect 20024 21448 20116 21450
rect 20024 21392 20074 21448
rect 20024 21390 20116 21392
rect 20069 21388 20116 21390
rect 20180 21388 20186 21452
rect 28349 21450 28415 21453
rect 29729 21450 29795 21453
rect 28349 21448 29795 21450
rect 28349 21392 28354 21448
rect 28410 21392 29734 21448
rect 29790 21392 29795 21448
rect 28349 21390 29795 21392
rect 20069 21387 20135 21388
rect 28349 21387 28415 21390
rect 29729 21387 29795 21390
rect 43253 21450 43319 21453
rect 44357 21450 44423 21453
rect 43253 21448 44423 21450
rect 43253 21392 43258 21448
rect 43314 21392 44362 21448
rect 44418 21392 44423 21448
rect 43253 21390 44423 21392
rect 43253 21387 43319 21390
rect 44357 21387 44423 21390
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 20713 20906 20779 20909
rect 21265 20906 21331 20909
rect 20713 20904 21331 20906
rect 20713 20848 20718 20904
rect 20774 20848 21270 20904
rect 21326 20848 21331 20904
rect 20713 20846 21331 20848
rect 20713 20843 20779 20846
rect 21265 20843 21331 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 43529 20498 43595 20501
rect 44725 20498 44791 20501
rect 43529 20496 44791 20498
rect 43529 20440 43534 20496
rect 43590 20440 44730 20496
rect 44786 20440 44791 20496
rect 43529 20438 44791 20440
rect 43529 20435 43595 20438
rect 44725 20435 44791 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 2957 19818 3023 19821
rect 19425 19820 19491 19821
rect 0 19816 3023 19818
rect 0 19760 2962 19816
rect 3018 19760 3023 19816
rect 0 19758 3023 19760
rect 0 19668 800 19758
rect 2957 19755 3023 19758
rect 19374 19756 19380 19820
rect 19444 19818 19491 19820
rect 19444 19816 19536 19818
rect 19486 19760 19536 19816
rect 19444 19758 19536 19760
rect 19444 19756 19491 19758
rect 19425 19755 19491 19756
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3417 18458 3483 18461
rect 0 18456 3483 18458
rect 0 18400 3422 18456
rect 3478 18400 3483 18456
rect 0 18398 3483 18400
rect 0 18308 800 18398
rect 3417 18395 3483 18398
rect 45829 18458 45895 18461
rect 49200 18458 50000 18548
rect 45829 18456 50000 18458
rect 45829 18400 45834 18456
rect 45890 18400 50000 18456
rect 45829 18398 50000 18400
rect 45829 18395 45895 18398
rect 49200 18308 50000 18398
rect 19333 18188 19399 18189
rect 19333 18184 19380 18188
rect 19444 18186 19450 18188
rect 19333 18128 19338 18184
rect 19333 18124 19380 18128
rect 19444 18126 19490 18186
rect 19444 18124 19450 18126
rect 19333 18123 19399 18124
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3417 17098 3483 17101
rect 0 17096 3483 17098
rect 0 17040 3422 17096
rect 3478 17040 3483 17096
rect 0 17038 3483 17040
rect 0 16948 800 17038
rect 3417 17035 3483 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 19374 14316 19380 14380
rect 19444 14378 19450 14380
rect 19977 14378 20043 14381
rect 19444 14376 20043 14378
rect 19444 14320 19982 14376
rect 20038 14320 20043 14376
rect 19444 14318 20043 14320
rect 19444 14316 19450 14318
rect 19977 14315 20043 14318
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13548 800 13638
rect 3417 13635 3483 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 2957 10298 3023 10301
rect 0 10296 3023 10298
rect 0 10240 2962 10296
rect 3018 10240 3023 10296
rect 0 10238 3023 10240
rect 0 10148 800 10238
rect 2957 10235 3023 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 47853 9618 47919 9621
rect 49200 9618 50000 9708
rect 47853 9616 50000 9618
rect 47853 9560 47858 9616
rect 47914 9560 50000 9616
rect 47853 9558 50000 9560
rect 47853 9555 47919 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 46841 8258 46907 8261
rect 49200 8258 50000 8348
rect 46841 8256 50000 8258
rect 46841 8200 46846 8256
rect 46902 8200 50000 8256
rect 46841 8198 50000 8200
rect 46841 8195 46907 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3509 7578 3575 7581
rect 0 7576 3575 7578
rect 0 7520 3514 7576
rect 3570 7520 3575 7576
rect 0 7518 3575 7520
rect 0 7428 800 7518
rect 3509 7515 3575 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3325 6898 3391 6901
rect 0 6896 3391 6898
rect 0 6840 3330 6896
rect 3386 6840 3391 6896
rect 0 6838 3391 6840
rect 0 6748 800 6838
rect 3325 6835 3391 6838
rect 46841 6898 46907 6901
rect 49200 6898 50000 6988
rect 46841 6896 50000 6898
rect 46841 6840 46846 6896
rect 46902 6840 50000 6896
rect 46841 6838 50000 6840
rect 46841 6835 46907 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 47945 6218 48011 6221
rect 49200 6218 50000 6308
rect 47945 6216 50000 6218
rect 47945 6160 47950 6216
rect 48006 6160 50000 6216
rect 47945 6158 50000 6160
rect 47945 6155 48011 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 49200 4028 50000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 3509 3498 3575 3501
rect 0 3496 3575 3498
rect 0 3440 3514 3496
rect 3570 3440 3575 3496
rect 0 3438 3575 3440
rect 0 3348 800 3438
rect 3509 3435 3575 3438
rect 17493 3498 17559 3501
rect 46197 3498 46263 3501
rect 17493 3496 46263 3498
rect 17493 3440 17498 3496
rect 17554 3440 46202 3496
rect 46258 3440 46263 3496
rect 17493 3438 46263 3440
rect 17493 3435 17559 3438
rect 46197 3435 46263 3438
rect 47945 3498 48011 3501
rect 49200 3498 50000 3588
rect 47945 3496 50000 3498
rect 47945 3440 47950 3496
rect 48006 3440 50000 3496
rect 47945 3438 50000 3440
rect 47945 3435 48011 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2668 800 2908
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1308 800 1398
rect 3417 1395 3483 1398
rect 46749 1458 46815 1461
rect 49200 1458 50000 1548
rect 46749 1456 50000 1458
rect 46749 1400 46754 1456
rect 46810 1400 50000 1456
rect 46749 1398 50000 1400
rect 46749 1395 46815 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 48037 778 48103 781
rect 49200 778 50000 868
rect 48037 776 50000 778
rect 48037 720 48042 776
rect 48098 720 50000 776
rect 48037 718 50000 720
rect 48037 715 48103 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 20116 24168 20180 24172
rect 20116 24112 20130 24168
rect 20130 24112 20180 24168
rect 20116 24108 20180 24112
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19380 22068 19444 22132
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 20116 21448 20180 21452
rect 20116 21392 20130 21448
rect 20130 21392 20180 21448
rect 20116 21388 20180 21392
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19380 19816 19444 19820
rect 19380 19760 19430 19816
rect 19430 19760 19444 19816
rect 19380 19756 19444 19760
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 19380 18184 19444 18188
rect 19380 18128 19394 18184
rect 19394 18128 19444 18184
rect 19380 18124 19444 18128
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19380 14316 19444 14380
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 20115 24172 20181 24173
rect 20115 24108 20116 24172
rect 20180 24108 20181 24172
rect 20115 24107 20181 24108
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19379 22132 19445 22133
rect 19379 22068 19380 22132
rect 19444 22068 19445 22132
rect 19379 22067 19445 22068
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 19382 19821 19442 22067
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 20118 21453 20178 24107
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 20115 21452 20181 21453
rect 20115 21388 20116 21452
rect 20180 21388 20181 21452
rect 20115 21387 20181 21388
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19379 19820 19445 19821
rect 19379 19756 19380 19820
rect 19444 19756 19445 19820
rect 19379 19755 19445 19756
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19379 18188 19445 18189
rect 19379 18124 19380 18188
rect 19444 18124 19445 18188
rect 19379 18123 19445 18124
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 19382 14381 19442 18123
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19379 14380 19445 14381
rect 19379 14316 19380 14380
rect 19444 14316 19445 14380
rect 19379 14315 19445 14316
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35972 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 45908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 33764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 41860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 37168 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_70 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1644511149
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1644511149
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_144
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_185
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_206
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_314
timestamp 1644511149
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_412
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_455
timestamp 1644511149
transform 1 0 42964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_80
timestamp 1644511149
transform 1 0 8464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1644511149
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1644511149
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1644511149
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_176
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1644511149
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1644511149
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1644511149
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_247
timestamp 1644511149
transform 1 0 23828 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_287
timestamp 1644511149
transform 1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_295
timestamp 1644511149
transform 1 0 28244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_307
timestamp 1644511149
transform 1 0 29348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_319
timestamp 1644511149
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1644511149
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_413
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_422
timestamp 1644511149
transform 1 0 39928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_426
timestamp 1644511149
transform 1 0 40296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_435
timestamp 1644511149
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_474
timestamp 1644511149
transform 1 0 44712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_62
timestamp 1644511149
transform 1 0 6808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1644511149
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_94
timestamp 1644511149
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1644511149
transform 1 0 10120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_123
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_131
timestamp 1644511149
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1644511149
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_214
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_222
timestamp 1644511149
transform 1 0 21528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_239
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1644511149
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_260
timestamp 1644511149
transform 1 0 25024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_267
timestamp 1644511149
transform 1 0 25668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_284
timestamp 1644511149
transform 1 0 27232 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_296
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_428
timestamp 1644511149
transform 1 0 40480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1644511149
transform 1 0 42780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_460
timestamp 1644511149
transform 1 0 43424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1644511149
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_87
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1644511149
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_138
timestamp 1644511149
transform 1 0 13800 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_144
timestamp 1644511149
transform 1 0 14352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp 1644511149
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1644511149
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_159
timestamp 1644511149
transform 1 0 15732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1644511149
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1644511149
transform 1 0 17204 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_186
timestamp 1644511149
transform 1 0 18216 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_198
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_203
timestamp 1644511149
transform 1 0 19780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_209
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1644511149
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_408
timestamp 1644511149
transform 1 0 38640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_415
timestamp 1644511149
transform 1 0 39284 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1644511149
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_465
timestamp 1644511149
transform 1 0 43884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_472
timestamp 1644511149
transform 1 0 44528 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_484
timestamp 1644511149
transform 1 0 45632 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_499
timestamp 1644511149
transform 1 0 47012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1644511149
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_155
timestamp 1644511149
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_162
timestamp 1644511149
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_169
timestamp 1644511149
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_176
timestamp 1644511149
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_188
timestamp 1644511149
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1644511149
transform 1 0 21160 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_225
timestamp 1644511149
transform 1 0 21804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1644511149
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_284
timestamp 1644511149
transform 1 0 27232 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_296
timestamp 1644511149
transform 1 0 28336 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1644511149
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_426
timestamp 1644511149
transform 1 0 40296 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_441
timestamp 1644511149
transform 1 0 41676 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_460
timestamp 1644511149
transform 1 0 43424 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_472
timestamp 1644511149
transform 1 0 44528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_399
timestamp 1644511149
transform 1 0 37812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_411
timestamp 1644511149
transform 1 0 38916 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_422
timestamp 1644511149
transform 1 0 39928 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_434
timestamp 1644511149
transform 1 0 41032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1644511149
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_399
timestamp 1644511149
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_403
timestamp 1644511149
transform 1 0 38180 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_394
timestamp 1644511149
transform 1 0 37352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_409
timestamp 1644511149
transform 1 0 38732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp 1644511149
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_489
timestamp 1644511149
transform 1 0 46092 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1644511149
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_481
timestamp 1644511149
transform 1 0 45356 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_495
timestamp 1644511149
transform 1 0 46644 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_505
timestamp 1644511149
transform 1 0 47564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1644511149
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_226
timestamp 1644511149
transform 1 0 21896 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_238
timestamp 1644511149
transform 1 0 23000 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1644511149
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_495
timestamp 1644511149
transform 1 0 46644 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_499
timestamp 1644511149
transform 1 0 47012 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_511
timestamp 1644511149
transform 1 0 48116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_515
timestamp 1644511149
transform 1 0 48484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_246
timestamp 1644511149
transform 1 0 23736 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_258
timestamp 1644511149
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1644511149
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1644511149
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 1644511149
transform 1 0 15916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1644511149
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1644511149
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_200
timestamp 1644511149
transform 1 0 19504 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_212
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_224
timestamp 1644511149
transform 1 0 21712 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_236
timestamp 1644511149
transform 1 0 22816 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_190
timestamp 1644511149
transform 1 0 18584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1644511149
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_242
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_254
timestamp 1644511149
transform 1 0 24472 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_266
timestamp 1644511149
transform 1 0 25576 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1644511149
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_180
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_184
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_218
timestamp 1644511149
transform 1 0 21160 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_224
timestamp 1644511149
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1644511149
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_504
timestamp 1644511149
transform 1 0 47472 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_148
timestamp 1644511149
transform 1 0 14720 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1644511149
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1644511149
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1644511149
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1644511149
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1644511149
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_233
timestamp 1644511149
transform 1 0 22540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1644511149
transform 1 0 23644 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1644511149
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_483
timestamp 1644511149
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_495
timestamp 1644511149
transform 1 0 46644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_508
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1644511149
transform 1 0 16468 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1644511149
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_204
timestamp 1644511149
transform 1 0 19872 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_210
timestamp 1644511149
transform 1 0 20424 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1644511149
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1644511149
transform 1 0 23092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_259
timestamp 1644511149
transform 1 0 24932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_271
timestamp 1644511149
transform 1 0 26036 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_283
timestamp 1644511149
transform 1 0 27140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_295
timestamp 1644511149
transform 1 0 28244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_464
timestamp 1644511149
transform 1 0 43792 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_507
timestamp 1644511149
transform 1 0 47748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1644511149
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_134
timestamp 1644511149
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_146
timestamp 1644511149
transform 1 0 14536 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_155
timestamp 1644511149
transform 1 0 15364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_173
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_180
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_192
timestamp 1644511149
transform 1 0 18768 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_232
timestamp 1644511149
transform 1 0 22448 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1644511149
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_268
timestamp 1644511149
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_286
timestamp 1644511149
transform 1 0 27416 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_294
timestamp 1644511149
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1644511149
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_309
timestamp 1644511149
transform 1 0 29532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_321
timestamp 1644511149
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1644511149
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_467
timestamp 1644511149
transform 1 0 44068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_492
timestamp 1644511149
transform 1 0 46368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_496
timestamp 1644511149
transform 1 0 46736 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_500
timestamp 1644511149
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_105
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 1644511149
transform 1 0 11316 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1644511149
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_150
timestamp 1644511149
transform 1 0 14904 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_162
timestamp 1644511149
transform 1 0 16008 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1644511149
transform 1 0 16744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_175
timestamp 1644511149
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1644511149
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1644511149
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_235
timestamp 1644511149
transform 1 0 22724 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1644511149
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_256
timestamp 1644511149
transform 1 0 24656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_268
timestamp 1644511149
transform 1 0 25760 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_280
timestamp 1644511149
transform 1 0 26864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1644511149
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_293
timestamp 1644511149
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_322
timestamp 1644511149
transform 1 0 30728 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_334
timestamp 1644511149
transform 1 0 31832 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_346
timestamp 1644511149
transform 1 0 32936 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_358
timestamp 1644511149
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_483
timestamp 1644511149
transform 1 0 45540 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_487
timestamp 1644511149
transform 1 0 45908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1644511149
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_154
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_191
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_203
timestamp 1644511149
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_207
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_211
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_232
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_296
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1644511149
transform 1 0 29256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1644511149
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1644511149
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1644511149
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_475
timestamp 1644511149
transform 1 0 44804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_510
timestamp 1644511149
transform 1 0 48024 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_129
timestamp 1644511149
transform 1 0 12972 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1644511149
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_173
timestamp 1644511149
transform 1 0 17020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1644511149
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1644511149
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_259
timestamp 1644511149
transform 1 0 24932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_268
timestamp 1644511149
transform 1 0 25760 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_278
timestamp 1644511149
transform 1 0 26680 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_290
timestamp 1644511149
transform 1 0 27784 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1644511149
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_313
timestamp 1644511149
transform 1 0 29900 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_337
timestamp 1644511149
transform 1 0 32108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1644511149
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_375
timestamp 1644511149
transform 1 0 35604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_379
timestamp 1644511149
transform 1 0 35972 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_391
timestamp 1644511149
transform 1 0 37076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_415
timestamp 1644511149
transform 1 0 39284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_462
timestamp 1644511149
transform 1 0 43608 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_468
timestamp 1644511149
transform 1 0 44160 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_485
timestamp 1644511149
transform 1 0 45724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1644511149
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_142
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_153
timestamp 1644511149
transform 1 0 15180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_175
timestamp 1644511149
transform 1 0 17204 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_187
timestamp 1644511149
transform 1 0 18308 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1644511149
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_198
timestamp 1644511149
transform 1 0 19320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_242
timestamp 1644511149
transform 1 0 23368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_253
timestamp 1644511149
transform 1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_260
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1644511149
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_302
timestamp 1644511149
transform 1 0 28888 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1644511149
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_360
timestamp 1644511149
transform 1 0 34224 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1644511149
transform 1 0 34868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1644511149
transform 1 0 35972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_457
timestamp 1644511149
transform 1 0 43148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_480
timestamp 1644511149
transform 1 0 45264 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_122
timestamp 1644511149
transform 1 0 12328 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_152
timestamp 1644511149
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_176
timestamp 1644511149
transform 1 0 17296 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1644511149
transform 1 0 19688 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_214
timestamp 1644511149
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_257
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_275
timestamp 1644511149
transform 1 0 26404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1644511149
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_316
timestamp 1644511149
transform 1 0 30176 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_324
timestamp 1644511149
transform 1 0 30912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_348
timestamp 1644511149
transform 1 0 33120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1644511149
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_483
timestamp 1644511149
transform 1 0 45540 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1644511149
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_101
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_116
timestamp 1644511149
transform 1 0 11776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_148
timestamp 1644511149
transform 1 0 14720 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_190
timestamp 1644511149
transform 1 0 18584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_197
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_209
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1644511149
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_233
timestamp 1644511149
transform 1 0 22540 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_239
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_251
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_263
timestamp 1644511149
transform 1 0 25300 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1644511149
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_285
timestamp 1644511149
transform 1 0 27324 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_297
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_304
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_316
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_324
timestamp 1644511149
transform 1 0 30912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_352
timestamp 1644511149
transform 1 0 33488 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_364
timestamp 1644511149
transform 1 0 34592 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_376
timestamp 1644511149
transform 1 0 35696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1644511149
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_457
timestamp 1644511149
transform 1 0 43148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_462
timestamp 1644511149
transform 1 0 43608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_466
timestamp 1644511149
transform 1 0 43976 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_470
timestamp 1644511149
transform 1 0 44344 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_482
timestamp 1644511149
transform 1 0 45448 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_490
timestamp 1644511149
transform 1 0 46184 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_499
timestamp 1644511149
transform 1 0 47012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_101
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1644511149
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1644511149
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_147
timestamp 1644511149
transform 1 0 14628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_158
timestamp 1644511149
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_170
timestamp 1644511149
transform 1 0 16744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_280
timestamp 1644511149
transform 1 0 26864 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_292
timestamp 1644511149
transform 1 0 27968 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1644511149
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_324
timestamp 1644511149
transform 1 0 30912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_349
timestamp 1644511149
transform 1 0 33212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_453
timestamp 1644511149
transform 1 0 42780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_467
timestamp 1644511149
transform 1 0 44068 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_504
timestamp 1644511149
transform 1 0 47472 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_511
timestamp 1644511149
transform 1 0 48116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_515
timestamp 1644511149
transform 1 0 48484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_133
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_141
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_172
timestamp 1644511149
transform 1 0 16928 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1644511149
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_204
timestamp 1644511149
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1644511149
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_228
timestamp 1644511149
transform 1 0 22080 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_236
timestamp 1644511149
transform 1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1644511149
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_251
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1644511149
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_340
timestamp 1644511149
transform 1 0 32384 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_365
timestamp 1644511149
transform 1 0 34684 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_377
timestamp 1644511149
transform 1 0 35788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1644511149
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_468
timestamp 1644511149
transform 1 0 44160 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_477
timestamp 1644511149
transform 1 0 44988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_486
timestamp 1644511149
transform 1 0 45816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_511
timestamp 1644511149
transform 1 0 48116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_515
timestamp 1644511149
transform 1 0 48484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_88
timestamp 1644511149
transform 1 0 9200 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_100
timestamp 1644511149
transform 1 0 10304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_106
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_116
timestamp 1644511149
transform 1 0 11776 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_128
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_162
timestamp 1644511149
transform 1 0 16008 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_203
timestamp 1644511149
transform 1 0 19780 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_211
timestamp 1644511149
transform 1 0 20516 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_226
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_230
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 1644511149
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_264
timestamp 1644511149
transform 1 0 25392 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1644511149
transform 1 0 26496 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_288
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_298
timestamp 1644511149
transform 1 0 28520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1644511149
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_312
timestamp 1644511149
transform 1 0 29808 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_320
timestamp 1644511149
transform 1 0 30544 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_344
timestamp 1644511149
transform 1 0 32752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1644511149
transform 1 0 33396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_449
timestamp 1644511149
transform 1 0 42412 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_453
timestamp 1644511149
transform 1 0 42780 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_464
timestamp 1644511149
transform 1 0 43792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_471
timestamp 1644511149
transform 1 0 44436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_481
timestamp 1644511149
transform 1 0 45356 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1644511149
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_77
timestamp 1644511149
transform 1 0 8188 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_99
timestamp 1644511149
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_119
timestamp 1644511149
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_128
timestamp 1644511149
transform 1 0 12880 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_136
timestamp 1644511149
transform 1 0 13616 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_140
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_148
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_154
timestamp 1644511149
transform 1 0 15272 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_160
timestamp 1644511149
transform 1 0 15824 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_191
timestamp 1644511149
transform 1 0 18676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_197
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1644511149
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_229
timestamp 1644511149
transform 1 0 22172 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_250
timestamp 1644511149
transform 1 0 24104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_288
timestamp 1644511149
transform 1 0 27600 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_297
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_312
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_318
timestamp 1644511149
transform 1 0 30360 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1644511149
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_350
timestamp 1644511149
transform 1 0 33304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_355
timestamp 1644511149
transform 1 0 33764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_363
timestamp 1644511149
transform 1 0 34500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_380
timestamp 1644511149
transform 1 0 36064 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_421
timestamp 1644511149
transform 1 0 39836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_427
timestamp 1644511149
transform 1 0 40388 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_439
timestamp 1644511149
transform 1 0 41492 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_460
timestamp 1644511149
transform 1 0 43424 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_481
timestamp 1644511149
transform 1 0 45356 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_489
timestamp 1644511149
transform 1 0 46092 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_111
timestamp 1644511149
transform 1 0 11316 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1644511149
transform 1 0 12420 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1644511149
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_154
timestamp 1644511149
transform 1 0 15272 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_166
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1644511149
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_206
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_222
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_230
timestamp 1644511149
transform 1 0 22264 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1644511149
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_261
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_267
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1644511149
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_312
timestamp 1644511149
transform 1 0 29808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_324
timestamp 1644511149
transform 1 0 30912 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_336
timestamp 1644511149
transform 1 0 32016 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_351
timestamp 1644511149
transform 1 0 33396 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_378
timestamp 1644511149
transform 1 0 35880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_390
timestamp 1644511149
transform 1 0 36984 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_402
timestamp 1644511149
transform 1 0 38088 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_414
timestamp 1644511149
transform 1 0 39192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_429
timestamp 1644511149
transform 1 0 40572 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_436
timestamp 1644511149
transform 1 0 41216 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_448
timestamp 1644511149
transform 1 0 42320 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_456
timestamp 1644511149
transform 1 0 43056 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_460
timestamp 1644511149
transform 1 0 43424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_464
timestamp 1644511149
transform 1 0 43792 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_470
timestamp 1644511149
transform 1 0 44344 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_480
timestamp 1644511149
transform 1 0 45264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_505
timestamp 1644511149
transform 1 0 47564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_98
timestamp 1644511149
transform 1 0 10120 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_118
timestamp 1644511149
transform 1 0 11960 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_128
timestamp 1644511149
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_132
timestamp 1644511149
transform 1 0 13248 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1644511149
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_157
timestamp 1644511149
transform 1 0 15548 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1644511149
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_192
timestamp 1644511149
transform 1 0 18768 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_196
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_228
timestamp 1644511149
transform 1 0 22080 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_240
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_262
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1644511149
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_285
timestamp 1644511149
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_296
timestamp 1644511149
transform 1 0 28336 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_320
timestamp 1644511149
transform 1 0 30544 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_340
timestamp 1644511149
transform 1 0 32384 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_352
timestamp 1644511149
transform 1 0 33488 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_374
timestamp 1644511149
transform 1 0 35512 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1644511149
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_413
timestamp 1644511149
transform 1 0 39100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_419
timestamp 1644511149
transform 1 0 39652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1644511149
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_455
timestamp 1644511149
transform 1 0 42964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_463
timestamp 1644511149
transform 1 0 43700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_470
timestamp 1644511149
transform 1 0 44344 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_478
timestamp 1644511149
transform 1 0 45080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_103
timestamp 1644511149
transform 1 0 10580 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1644511149
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_115
timestamp 1644511149
transform 1 0 11684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_122
timestamp 1644511149
transform 1 0 12328 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_162
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_186
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_214
timestamp 1644511149
transform 1 0 20792 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_226
timestamp 1644511149
transform 1 0 21896 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_234
timestamp 1644511149
transform 1 0 22632 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_239
timestamp 1644511149
transform 1 0 23092 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1644511149
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_269
timestamp 1644511149
transform 1 0 25852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_281
timestamp 1644511149
transform 1 0 26956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_293
timestamp 1644511149
transform 1 0 28060 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_298
timestamp 1644511149
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1644511149
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_315
timestamp 1644511149
transform 1 0 30084 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_337
timestamp 1644511149
transform 1 0 32108 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_349
timestamp 1644511149
transform 1 0 33212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_353
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_378
timestamp 1644511149
transform 1 0 35880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_390
timestamp 1644511149
transform 1 0 36984 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_402
timestamp 1644511149
transform 1 0 38088 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_414
timestamp 1644511149
transform 1 0 39192 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_442
timestamp 1644511149
transform 1 0 41768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_452
timestamp 1644511149
transform 1 0 42688 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_458
timestamp 1644511149
transform 1 0 43240 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1644511149
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_483
timestamp 1644511149
transform 1 0 45540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_487
timestamp 1644511149
transform 1 0 45908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_97
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_102
timestamp 1644511149
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1644511149
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1644511149
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_153
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1644511149
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_195
timestamp 1644511149
transform 1 0 19044 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1644511149
transform 1 0 23460 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_248
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_256
timestamp 1644511149
transform 1 0 24656 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_268
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_340
timestamp 1644511149
transform 1 0 32384 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_352
timestamp 1644511149
transform 1 0 33488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_360
timestamp 1644511149
transform 1 0 34224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_365
timestamp 1644511149
transform 1 0 34684 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_424
timestamp 1644511149
transform 1 0 40112 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_435
timestamp 1644511149
transform 1 0 41124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_457
timestamp 1644511149
transform 1 0 43148 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_463
timestamp 1644511149
transform 1 0 43700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_470
timestamp 1644511149
transform 1 0 44344 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_482
timestamp 1644511149
transform 1 0 45448 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_486
timestamp 1644511149
transform 1 0 45816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_120
timestamp 1644511149
transform 1 0 12144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1644511149
transform 1 0 16744 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_178
timestamp 1644511149
transform 1 0 17480 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_184
timestamp 1644511149
transform 1 0 18032 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_201
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_208
timestamp 1644511149
transform 1 0 20240 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_220
timestamp 1644511149
transform 1 0 21344 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_232
timestamp 1644511149
transform 1 0 22448 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_243
timestamp 1644511149
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1644511149
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_312
timestamp 1644511149
transform 1 0 29808 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_320
timestamp 1644511149
transform 1 0 30544 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_342
timestamp 1644511149
transform 1 0 32568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_354
timestamp 1644511149
transform 1 0 33672 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_390
timestamp 1644511149
transform 1 0 36984 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_402
timestamp 1644511149
transform 1 0 38088 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_414
timestamp 1644511149
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_442
timestamp 1644511149
transform 1 0 41768 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_454
timestamp 1644511149
transform 1 0 42872 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_466
timestamp 1644511149
transform 1 0 43976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_474
timestamp 1644511149
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_480
timestamp 1644511149
transform 1 0 45264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_487
timestamp 1644511149
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1644511149
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_116
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_128
timestamp 1644511149
transform 1 0 12880 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_140
timestamp 1644511149
transform 1 0 13984 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1644511149
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_176
timestamp 1644511149
transform 1 0 17296 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_184
timestamp 1644511149
transform 1 0 18032 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_253
timestamp 1644511149
transform 1 0 24380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_284
timestamp 1644511149
transform 1 0 27232 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_292
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_313
timestamp 1644511149
transform 1 0 29900 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_321
timestamp 1644511149
transform 1 0 30636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1644511149
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_341
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_348
timestamp 1644511149
transform 1 0 33120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_360
timestamp 1644511149
transform 1 0 34224 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_368
timestamp 1644511149
transform 1 0 34960 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_378
timestamp 1644511149
transform 1 0 35880 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1644511149
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_421
timestamp 1644511149
transform 1 0 39836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_425
timestamp 1644511149
transform 1 0 40204 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_437
timestamp 1644511149
transform 1 0 41308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1644511149
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1644511149
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_122
timestamp 1644511149
transform 1 0 12328 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1644511149
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_151
timestamp 1644511149
transform 1 0 14996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_168
timestamp 1644511149
transform 1 0 16560 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_200
timestamp 1644511149
transform 1 0 19504 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_213
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_217
timestamp 1644511149
transform 1 0 21068 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_226
timestamp 1644511149
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1644511149
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_256
timestamp 1644511149
transform 1 0 24656 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1644511149
transform 1 0 26036 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1644511149
transform 1 0 27048 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1644511149
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1644511149
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_313
timestamp 1644511149
transform 1 0 29900 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_329
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_337
timestamp 1644511149
transform 1 0 32108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_375
timestamp 1644511149
transform 1 0 35604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_387
timestamp 1644511149
transform 1 0 36708 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_399
timestamp 1644511149
transform 1 0 37812 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_411
timestamp 1644511149
transform 1 0 38916 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_97
timestamp 1644511149
transform 1 0 10028 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_121
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_128
timestamp 1644511149
transform 1 0 12880 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_152
timestamp 1644511149
transform 1 0 15088 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 1644511149
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_194
timestamp 1644511149
transform 1 0 18952 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1644511149
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_233
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_255
timestamp 1644511149
transform 1 0 24564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_267
timestamp 1644511149
transform 1 0 25668 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_286
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_294
timestamp 1644511149
transform 1 0 28152 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_300
timestamp 1644511149
transform 1 0 28704 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_308
timestamp 1644511149
transform 1 0 29440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_314
timestamp 1644511149
transform 1 0 29992 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_322
timestamp 1644511149
transform 1 0 30728 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_326
timestamp 1644511149
transform 1 0 31096 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_340
timestamp 1644511149
transform 1 0 32384 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_351
timestamp 1644511149
transform 1 0 33396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_101
timestamp 1644511149
transform 1 0 10396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_113
timestamp 1644511149
transform 1 0 11500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_117
timestamp 1644511149
transform 1 0 11868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_122
timestamp 1644511149
transform 1 0 12328 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1644511149
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_148
timestamp 1644511149
transform 1 0 14720 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_157
timestamp 1644511149
transform 1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_172
timestamp 1644511149
transform 1 0 16928 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_180
timestamp 1644511149
transform 1 0 17664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_215
timestamp 1644511149
transform 1 0 20884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_228
timestamp 1644511149
transform 1 0 22080 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_236
timestamp 1644511149
transform 1 0 22816 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_258
timestamp 1644511149
transform 1 0 24840 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_266
timestamp 1644511149
transform 1 0 25576 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_286
timestamp 1644511149
transform 1 0 27416 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_300
timestamp 1644511149
transform 1 0 28704 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_318
timestamp 1644511149
transform 1 0 30360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_326
timestamp 1644511149
transform 1 0 31096 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_339
timestamp 1644511149
transform 1 0 32292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_349
timestamp 1644511149
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1644511149
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_507
timestamp 1644511149
transform 1 0 47748 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_515
timestamp 1644511149
transform 1 0 48484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_118
timestamp 1644511149
transform 1 0 11960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_130
timestamp 1644511149
transform 1 0 13064 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_138
timestamp 1644511149
transform 1 0 13800 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_144
timestamp 1644511149
transform 1 0 14352 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_156
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_211
timestamp 1644511149
transform 1 0 20516 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1644511149
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_244
timestamp 1644511149
transform 1 0 23552 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_251
timestamp 1644511149
transform 1 0 24196 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_263
timestamp 1644511149
transform 1 0 25300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_272
timestamp 1644511149
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1644511149
transform 1 0 28520 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_310
timestamp 1644511149
transform 1 0 29624 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_322
timestamp 1644511149
transform 1 0 30728 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 1644511149
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_124
timestamp 1644511149
transform 1 0 12512 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_132
timestamp 1644511149
transform 1 0 13248 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_145
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_157
timestamp 1644511149
transform 1 0 15548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_169
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_181
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1644511149
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_222
timestamp 1644511149
transform 1 0 21528 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_234
timestamp 1644511149
transform 1 0 22632 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_273
timestamp 1644511149
transform 1 0 26220 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_278
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1644511149
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_316
timestamp 1644511149
transform 1 0 30176 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_328
timestamp 1644511149
transform 1 0 31280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_338
timestamp 1644511149
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_350
timestamp 1644511149
transform 1 0 33304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1644511149
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_99
timestamp 1644511149
transform 1 0 10212 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_104
timestamp 1644511149
transform 1 0 10672 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_120
timestamp 1644511149
transform 1 0 12144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1644511149
transform 1 0 12788 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_148
timestamp 1644511149
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_155
timestamp 1644511149
transform 1 0 15364 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_190
timestamp 1644511149
transform 1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_214
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1644511149
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_234
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_246
timestamp 1644511149
transform 1 0 23736 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_258
timestamp 1644511149
transform 1 0 24840 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_288
timestamp 1644511149
transform 1 0 27600 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_296
timestamp 1644511149
transform 1 0 28336 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_318
timestamp 1644511149
transform 1 0 30360 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_326
timestamp 1644511149
transform 1 0 31096 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_359
timestamp 1644511149
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_371
timestamp 1644511149
transform 1 0 35236 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_383
timestamp 1644511149
transform 1 0 36340 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_93
timestamp 1644511149
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_99
timestamp 1644511149
transform 1 0 10212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_106
timestamp 1644511149
transform 1 0 10856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_113
timestamp 1644511149
transform 1 0 11500 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_125
timestamp 1644511149
transform 1 0 12604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1644511149
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_161
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_168
timestamp 1644511149
transform 1 0 16560 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_179
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_187
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_217
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_228
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_237
timestamp 1644511149
transform 1 0 22908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_276
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_292
timestamp 1644511149
transform 1 0 27968 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_300
timestamp 1644511149
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_317
timestamp 1644511149
transform 1 0 30268 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_326
timestamp 1644511149
transform 1 0 31096 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_332
timestamp 1644511149
transform 1 0 31648 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_339
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_347
timestamp 1644511149
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1644511149
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_368
timestamp 1644511149
transform 1 0 34960 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_380
timestamp 1644511149
transform 1 0 36064 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_392
timestamp 1644511149
transform 1 0 37168 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_404
timestamp 1644511149
transform 1 0 38272 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_416
timestamp 1644511149
transform 1 0 39376 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_507
timestamp 1644511149
transform 1 0 47748 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_515
timestamp 1644511149
transform 1 0 48484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1644511149
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_134
timestamp 1644511149
transform 1 0 13432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_142
timestamp 1644511149
transform 1 0 14168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_190
timestamp 1644511149
transform 1 0 18584 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_199
timestamp 1644511149
transform 1 0 19412 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_209
timestamp 1644511149
transform 1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1644511149
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_228
timestamp 1644511149
transform 1 0 22080 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_240
timestamp 1644511149
transform 1 0 23184 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_291
timestamp 1644511149
transform 1 0 27876 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_298
timestamp 1644511149
transform 1 0 28520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_306
timestamp 1644511149
transform 1 0 29256 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_311
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_319
timestamp 1644511149
transform 1 0 30452 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_347
timestamp 1644511149
transform 1 0 33028 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_355
timestamp 1644511149
transform 1 0 33764 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_377
timestamp 1644511149
transform 1 0 35788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1644511149
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_144
timestamp 1644511149
transform 1 0 14352 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_169
timestamp 1644511149
transform 1 0 16652 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_181
timestamp 1644511149
transform 1 0 17756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1644511149
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_217
timestamp 1644511149
transform 1 0 21068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_237
timestamp 1644511149
transform 1 0 22908 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1644511149
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_262
timestamp 1644511149
transform 1 0 25208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_269
timestamp 1644511149
transform 1 0 25852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_285
timestamp 1644511149
transform 1 0 27324 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_293
timestamp 1644511149
transform 1 0 28060 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_317
timestamp 1644511149
transform 1 0 30268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_323
timestamp 1644511149
transform 1 0 30820 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_334
timestamp 1644511149
transform 1 0 31832 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_344
timestamp 1644511149
transform 1 0 32752 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1644511149
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_155
timestamp 1644511149
transform 1 0 15364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_198
timestamp 1644511149
transform 1 0 19320 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_253
timestamp 1644511149
transform 1 0 24380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_264
timestamp 1644511149
transform 1 0 25392 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1644511149
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_286
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_298
timestamp 1644511149
transform 1 0 28520 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1644511149
transform 1 0 29624 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_322
timestamp 1644511149
transform 1 0 30728 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_326
timestamp 1644511149
transform 1 0 31096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1644511149
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_347
timestamp 1644511149
transform 1 0 33028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_360
timestamp 1644511149
transform 1 0 34224 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_364
timestamp 1644511149
transform 1 0 34592 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_368
timestamp 1644511149
transform 1 0 34960 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_380
timestamp 1644511149
transform 1 0 36064 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_205
timestamp 1644511149
transform 1 0 19964 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_214
timestamp 1644511149
transform 1 0 20792 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_222
timestamp 1644511149
transform 1 0 21528 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_239
timestamp 1644511149
transform 1 0 23092 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1644511149
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_264
timestamp 1644511149
transform 1 0 25392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_271
timestamp 1644511149
transform 1 0 26036 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_279
timestamp 1644511149
transform 1 0 26772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_288
timestamp 1644511149
transform 1 0 27600 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_296
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_300
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_329
timestamp 1644511149
transform 1 0 31372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_342
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_351
timestamp 1644511149
transform 1 0 33396 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1644511149
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_385
timestamp 1644511149
transform 1 0 36524 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_397
timestamp 1644511149
transform 1 0 37628 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_409
timestamp 1644511149
transform 1 0 38732 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_417
timestamp 1644511149
transform 1 0 39468 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_495
timestamp 1644511149
transform 1 0 46644 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_509
timestamp 1644511149
transform 1 0 47932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_515
timestamp 1644511149
transform 1 0 48484 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1644511149
transform 1 0 20240 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_239
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_243
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_250
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_260
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_268
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_313
timestamp 1644511149
transform 1 0 29900 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_321
timestamp 1644511149
transform 1 0 30636 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_7
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_14
timestamp 1644511149
transform 1 0 2392 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1644511149
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_50
timestamp 1644511149
transform 1 0 5704 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_62
timestamp 1644511149
transform 1 0 6808 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_74
timestamp 1644511149
transform 1 0 7912 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1644511149
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_182
timestamp 1644511149
transform 1 0 17848 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_201
timestamp 1644511149
transform 1 0 19596 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_213
timestamp 1644511149
transform 1 0 20700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_230
timestamp 1644511149
transform 1 0 22264 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_240
timestamp 1644511149
transform 1 0 23184 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_263
timestamp 1644511149
transform 1 0 25300 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_291
timestamp 1644511149
transform 1 0 27876 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_298
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1644511149
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_316
timestamp 1644511149
transform 1 0 30176 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_328
timestamp 1644511149
transform 1 0 31280 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_352
timestamp 1644511149
transform 1 0 33488 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_28
timestamp 1644511149
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_40
timestamp 1644511149
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_213
timestamp 1644511149
transform 1 0 20700 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_235
timestamp 1644511149
transform 1 0 22724 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_245
timestamp 1644511149
transform 1 0 23644 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_262
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_274
timestamp 1644511149
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_284
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_294
timestamp 1644511149
transform 1 0 28152 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_310
timestamp 1644511149
transform 1 0 29624 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_358
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_370
timestamp 1644511149
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1644511149
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1644511149
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_13
timestamp 1644511149
transform 1 0 2300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1644511149
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1644511149
transform 1 0 4048 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1644511149
transform 1 0 5152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1644511149
transform 1 0 6256 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1644511149
transform 1 0 7360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_217
timestamp 1644511149
transform 1 0 21068 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_225
timestamp 1644511149
transform 1 0 21804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_240
timestamp 1644511149
transform 1 0 23184 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_259
timestamp 1644511149
transform 1 0 24932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_271
timestamp 1644511149
transform 1 0 26036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_279
timestamp 1644511149
transform 1 0 26772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_290
timestamp 1644511149
transform 1 0 27784 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_297
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1644511149
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_316
timestamp 1644511149
transform 1 0 30176 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_324
timestamp 1644511149
transform 1 0 30912 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_331
timestamp 1644511149
transform 1 0 31556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_343
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_355
timestamp 1644511149
transform 1 0 33764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_498
timestamp 1644511149
transform 1 0 46920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_6
timestamp 1644511149
transform 1 0 1656 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_33
timestamp 1644511149
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1644511149
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1644511149
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_201
timestamp 1644511149
transform 1 0 19596 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_206
timestamp 1644511149
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_218
timestamp 1644511149
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_231
timestamp 1644511149
transform 1 0 22356 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_243
timestamp 1644511149
transform 1 0 23460 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_267
timestamp 1644511149
transform 1 0 25668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_301
timestamp 1644511149
transform 1 0 28796 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_323
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_493
timestamp 1644511149
transform 1 0 46460 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_511
timestamp 1644511149
transform 1 0 48116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_515
timestamp 1644511149
transform 1 0 48484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_203
timestamp 1644511149
transform 1 0 19780 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_211
timestamp 1644511149
transform 1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1644511149
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_234
timestamp 1644511149
transform 1 0 22632 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_242
timestamp 1644511149
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1644511149
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_281
timestamp 1644511149
transform 1 0 26956 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_287
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_295
timestamp 1644511149
transform 1 0 28244 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_302
timestamp 1644511149
transform 1 0 28888 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_315
timestamp 1644511149
transform 1 0 30084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_323
timestamp 1644511149
transform 1 0 30820 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_331
timestamp 1644511149
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1644511149
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_355
timestamp 1644511149
transform 1 0 33764 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_189
timestamp 1644511149
transform 1 0 18492 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_210
timestamp 1644511149
transform 1 0 20424 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1644511149
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_233
timestamp 1644511149
transform 1 0 22540 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_242
timestamp 1644511149
transform 1 0 23368 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_254
timestamp 1644511149
transform 1 0 24472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_258
timestamp 1644511149
transform 1 0 24840 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_270
timestamp 1644511149
transform 1 0 25944 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1644511149
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_291
timestamp 1644511149
transform 1 0 27876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_299
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_304
timestamp 1644511149
transform 1 0 29072 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_308
timestamp 1644511149
transform 1 0 29440 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_314
timestamp 1644511149
transform 1 0 29992 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_324
timestamp 1644511149
transform 1 0 30912 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_217
timestamp 1644511149
transform 1 0 21068 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_230
timestamp 1644511149
transform 1 0 22264 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_238
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1644511149
transform 1 0 24840 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_270
timestamp 1644511149
transform 1 0 25944 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_300
timestamp 1644511149
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_316
timestamp 1644511149
transform 1 0 30176 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_329
timestamp 1644511149
transform 1 0 31372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_342
timestamp 1644511149
transform 1 0 32568 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_354
timestamp 1644511149
transform 1 0 33672 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1644511149
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_216
timestamp 1644511149
transform 1 0 20976 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_234
timestamp 1644511149
transform 1 0 22632 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_244
timestamp 1644511149
transform 1 0 23552 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_252
timestamp 1644511149
transform 1 0 24288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_258
timestamp 1644511149
transform 1 0 24840 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_268
timestamp 1644511149
transform 1 0 25760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_290
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_299
timestamp 1644511149
transform 1 0 28612 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_319
timestamp 1644511149
transform 1 0 30452 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 1644511149
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_357
timestamp 1644511149
transform 1 0 33948 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_369
timestamp 1644511149
transform 1 0 35052 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_381
timestamp 1644511149
transform 1 0 36156 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1644511149
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1644511149
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_203
timestamp 1644511149
transform 1 0 19780 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_207
timestamp 1644511149
transform 1 0 20148 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_235
timestamp 1644511149
transform 1 0 22724 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1644511149
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_260
timestamp 1644511149
transform 1 0 25024 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1644511149
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_296
timestamp 1644511149
transform 1 0 28336 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_316
timestamp 1644511149
transform 1 0 30176 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_325
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1644511149
transform 1 0 32292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1644511149
transform 1 0 33396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_231
timestamp 1644511149
transform 1 0 22356 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_243
timestamp 1644511149
transform 1 0 23460 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_255
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_260
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1644511149
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_288
timestamp 1644511149
transform 1 0 27600 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_300
timestamp 1644511149
transform 1 0 28704 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_308
timestamp 1644511149
transform 1 0 29440 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_203
timestamp 1644511149
transform 1 0 19780 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_215
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_223
timestamp 1644511149
transform 1 0 21620 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_228
timestamp 1644511149
transform 1 0 22080 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_240
timestamp 1644511149
transform 1 0 23184 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_258
timestamp 1644511149
transform 1 0 24840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_268
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_276
timestamp 1644511149
transform 1 0 26496 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_280
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_209
timestamp 1644511149
transform 1 0 20332 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_216
timestamp 1644511149
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_257
timestamp 1644511149
transform 1 0 24748 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_263
timestamp 1644511149
transform 1 0 25300 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_267
timestamp 1644511149
transform 1 0 25668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_301
timestamp 1644511149
transform 1 0 28796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_308
timestamp 1644511149
transform 1 0 29440 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_320
timestamp 1644511149
transform 1 0 30544 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1644511149
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_185
timestamp 1644511149
transform 1 0 18124 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_192
timestamp 1644511149
transform 1 0 18768 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_222
timestamp 1644511149
transform 1 0 21528 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_234
timestamp 1644511149
transform 1 0 22632 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_240
timestamp 1644511149
transform 1 0 23184 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1644511149
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_273
timestamp 1644511149
transform 1 0 26220 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_285
timestamp 1644511149
transform 1 0 27324 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_294
timestamp 1644511149
transform 1 0 28152 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1644511149
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_507
timestamp 1644511149
transform 1 0 47748 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_515
timestamp 1644511149
transform 1 0 48484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_209
timestamp 1644511149
transform 1 0 20332 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1644511149
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_248
timestamp 1644511149
transform 1 0 23920 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_229
timestamp 1644511149
transform 1 0 22172 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_235
timestamp 1644511149
transform 1 0 22724 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1644511149
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_257
timestamp 1644511149
transform 1 0 24748 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_267
timestamp 1644511149
transform 1 0 25668 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_279
timestamp 1644511149
transform 1 0 26772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_291
timestamp 1644511149
transform 1 0 27876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_303
timestamp 1644511149
transform 1 0 28980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_499
timestamp 1644511149
transform 1 0 47012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_488
timestamp 1644511149
transform 1 0 46000 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_495
timestamp 1644511149
transform 1 0 46644 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1644511149
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_282
timestamp 1644511149
transform 1 0 27048 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_294
timestamp 1644511149
transform 1 0 28152 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1644511149
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_428
timestamp 1644511149
transform 1 0 40480 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_440
timestamp 1644511149
transform 1 0 41584 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_472
timestamp 1644511149
transform 1 0 44528 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_407
timestamp 1644511149
transform 1 0 38548 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_411
timestamp 1644511149
transform 1 0 38916 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_453
timestamp 1644511149
transform 1 0 42780 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_458
timestamp 1644511149
transform 1 0 43240 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_466
timestamp 1644511149
transform 1 0 43976 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_485
timestamp 1644511149
transform 1 0 45724 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_14
timestamp 1644511149
transform 1 0 2392 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_26
timestamp 1644511149
transform 1 0 3496 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_38
timestamp 1644511149
transform 1 0 4600 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 1644511149
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_101
timestamp 1644511149
transform 1 0 10396 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_269
timestamp 1644511149
transform 1 0 25852 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_274
timestamp 1644511149
transform 1 0 26312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_452
timestamp 1644511149
transform 1 0 42688 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_460
timestamp 1644511149
transform 1 0 43424 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_464
timestamp 1644511149
transform 1 0 43792 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_489
timestamp 1644511149
transform 1 0 46092 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1644511149
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_33
timestamp 1644511149
transform 1 0 4140 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_37
timestamp 1644511149
transform 1 0 4508 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_46
timestamp 1644511149
transform 1 0 5336 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_58
timestamp 1644511149
transform 1 0 6440 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_70
timestamp 1644511149
transform 1 0 7544 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1644511149
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_122
timestamp 1644511149
transform 1 0 12328 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_134
timestamp 1644511149
transform 1 0 13432 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_188
timestamp 1644511149
transform 1 0 18400 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_203
timestamp 1644511149
transform 1 0 19780 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_228
timestamp 1644511149
transform 1 0 22080 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_240
timestamp 1644511149
transform 1 0 23184 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_261
timestamp 1644511149
transform 1 0 25116 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_290
timestamp 1644511149
transform 1 0 27784 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_302
timestamp 1644511149
transform 1 0 28888 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_458
timestamp 1644511149
transform 1 0 43240 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_464
timestamp 1644511149
transform 1 0 43792 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_13
timestamp 1644511149
transform 1 0 2300 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_20
timestamp 1644511149
transform 1 0 2944 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_28
timestamp 1644511149
transform 1 0 3680 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_132
timestamp 1644511149
transform 1 0 13248 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_157
timestamp 1644511149
transform 1 0 15548 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_165
timestamp 1644511149
transform 1 0 16284 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_189
timestamp 1644511149
transform 1 0 18492 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_195
timestamp 1644511149
transform 1 0 19044 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_266
timestamp 1644511149
transform 1 0 25576 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_275
timestamp 1644511149
transform 1 0 26404 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_302
timestamp 1644511149
transform 1 0 28888 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_314
timestamp 1644511149
transform 1 0 29992 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_326
timestamp 1644511149
transform 1 0 31096 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_358
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_370
timestamp 1644511149
transform 1 0 35144 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_382
timestamp 1644511149
transform 1 0 36248 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_390
timestamp 1644511149
transform 1 0 36984 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1644511149
transform 1 0 6900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_118
timestamp 1644511149
transform 1 0 11960 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1644511149
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_151
timestamp 1644511149
transform 1 0 14996 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_159
timestamp 1644511149
transform 1 0 15732 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_207
timestamp 1644511149
transform 1 0 20148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_214
timestamp 1644511149
transform 1 0 20792 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_222
timestamp 1644511149
transform 1 0 21528 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_228
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_240
timestamp 1644511149
transform 1 0 23184 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_444
timestamp 1644511149
transform 1 0 41952 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32660 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31188 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0601_
timestamp 1644511149
transform 1 0 32936 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0603_
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0604_
timestamp 1644511149
transform 1 0 24748 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0605_
timestamp 1644511149
transform 1 0 23092 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0606_
timestamp 1644511149
transform 1 0 30360 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0607_
timestamp 1644511149
transform 1 0 25208 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0608_
timestamp 1644511149
transform 1 0 25392 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0611_
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0612_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0614_
timestamp 1644511149
transform 1 0 26864 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0615_
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1644511149
transform 1 0 26772 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0620_
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0621_
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0622_
timestamp 1644511149
transform 1 0 22264 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0623_
timestamp 1644511149
transform 1 0 19504 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0624_
timestamp 1644511149
transform 1 0 21528 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0625_
timestamp 1644511149
transform 1 0 14076 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0626_
timestamp 1644511149
transform 1 0 15364 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0627_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0628_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0630_
timestamp 1644511149
transform 1 0 28336 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1644511149
transform 1 0 27048 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0633_
timestamp 1644511149
transform 1 0 27968 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0634_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1644511149
transform 1 0 25392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0639_
timestamp 1644511149
transform 1 0 24748 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0641_
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0642_
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0643_
timestamp 1644511149
transform 1 0 21988 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0644_
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0646_
timestamp 1644511149
transform 1 0 20240 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0648_
timestamp 1644511149
transform 1 0 20424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0651_
timestamp 1644511149
transform 1 0 17112 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0653_
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1644511149
transform 1 0 14536 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 1644511149
transform 1 0 15088 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0656_
timestamp 1644511149
transform 1 0 11960 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0657_
timestamp 1644511149
transform 1 0 16560 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1644511149
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1644511149
transform 1 0 18216 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0660_
timestamp 1644511149
transform 1 0 14352 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 1644511149
transform 1 0 13340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0665_
timestamp 1644511149
transform 1 0 14904 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1644511149
transform 1 0 14076 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0670_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1644511149
transform 1 0 12512 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0674_
timestamp 1644511149
transform 1 0 11224 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1644511149
transform 1 0 12328 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 1644511149
transform 1 0 10580 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0677_
timestamp 1644511149
transform 1 0 10396 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1644511149
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0680_
timestamp 1644511149
transform 1 0 10120 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0682_
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0683_
timestamp 1644511149
transform 1 0 12788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0684_
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1644511149
transform 1 0 10672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0687_
timestamp 1644511149
transform 1 0 12420 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0688_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1644511149
transform 1 0 11960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0690_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11224 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0692_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0694_
timestamp 1644511149
transform 1 0 10396 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0695_
timestamp 1644511149
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1644511149
transform 1 0 16744 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0698_
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0701_
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0702_
timestamp 1644511149
transform 1 0 14536 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0704_
timestamp 1644511149
transform 1 0 14536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 1644511149
transform 1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1644511149
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0707_
timestamp 1644511149
transform 1 0 14076 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1644511149
transform 1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0709_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0710_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0711_
timestamp 1644511149
transform 1 0 18400 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0712_
timestamp 1644511149
transform 1 0 17296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0713_
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0714_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1644511149
transform 1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0716_
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0717_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 20240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0719_
timestamp 1644511149
transform 1 0 18124 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0721_
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0722_
timestamp 1644511149
transform 1 0 22080 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 1644511149
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 24656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_
timestamp 1644511149
transform 1 0 22816 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23736 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0728_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1644511149
transform 1 0 23092 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0733_
timestamp 1644511149
transform 1 0 25760 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1644511149
transform 1 0 28796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0735_
timestamp 1644511149
transform 1 0 25576 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1644511149
transform 1 0 25944 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0738_
timestamp 1644511149
transform 1 0 29624 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0739_
timestamp 1644511149
transform 1 0 30728 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0740_
timestamp 1644511149
transform 1 0 28152 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0743_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0744_
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1644511149
transform 1 0 28244 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0746_
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1644511149
transform 1 0 26956 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0748_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0749_
timestamp 1644511149
transform 1 0 27784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0750_
timestamp 1644511149
transform 1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0751_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0752_
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26404 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0755_
timestamp 1644511149
transform 1 0 23276 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0756_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0757_
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0758_
timestamp 1644511149
transform 1 0 28704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0759_
timestamp 1644511149
transform 1 0 22908 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0761_
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0762_
timestamp 1644511149
transform 1 0 23000 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0763_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0764_
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0765_
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0766_
timestamp 1644511149
transform 1 0 26864 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0767_
timestamp 1644511149
transform 1 0 27968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1644511149
transform 1 0 20240 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0771_
timestamp 1644511149
transform 1 0 28336 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0773_
timestamp 1644511149
transform 1 0 20700 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0774_
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0775_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0776_
timestamp 1644511149
transform 1 0 30452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0777_
timestamp 1644511149
transform 1 0 27048 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0778_
timestamp 1644511149
transform 1 0 20148 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0779_
timestamp 1644511149
transform 1 0 20700 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0780_
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1644511149
transform 1 0 20056 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0783_
timestamp 1644511149
transform 1 0 19504 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0784_
timestamp 1644511149
transform 1 0 20792 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0786_
timestamp 1644511149
transform 1 0 24472 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0787_
timestamp 1644511149
transform 1 0 23000 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0788_
timestamp 1644511149
transform 1 0 21252 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0789_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0790_
timestamp 1644511149
transform 1 0 25208 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0792_
timestamp 1644511149
transform 1 0 24472 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1644511149
transform 1 0 22908 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0795_
timestamp 1644511149
transform 1 0 27140 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1644511149
transform 1 0 30360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0797_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0798_
timestamp 1644511149
transform 1 0 23552 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0799_
timestamp 1644511149
transform 1 0 24288 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1644511149
transform 1 0 28060 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0801_
timestamp 1644511149
transform 1 0 29900 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0803_
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0805_
timestamp 1644511149
transform 1 0 27140 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0806_
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0807_
timestamp 1644511149
transform 1 0 30084 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0808_
timestamp 1644511149
transform 1 0 27508 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0809_
timestamp 1644511149
transform 1 0 26220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0810_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0811_
timestamp 1644511149
transform 1 0 27048 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0812_
timestamp 1644511149
transform 1 0 23000 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0813_
timestamp 1644511149
transform 1 0 29532 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0814_
timestamp 1644511149
transform 1 0 30820 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0815_
timestamp 1644511149
transform 1 0 30728 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0816_
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1644511149
transform 1 0 30544 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0818_
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0819_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0820_
timestamp 1644511149
transform 1 0 31188 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1644511149
transform 1 0 31280 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0822_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0823_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0824_
timestamp 1644511149
transform 1 0 28980 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0825_
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0826_
timestamp 1644511149
transform 1 0 28888 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0827_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0829_
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0830_
timestamp 1644511149
transform 1 0 30820 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1644511149
transform 1 0 22632 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0832_
timestamp 1644511149
transform 1 0 25760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0833_
timestamp 1644511149
transform 1 0 26036 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0834_
timestamp 1644511149
transform 1 0 26956 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1644511149
transform 1 0 26956 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0837_
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0838_
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0839_
timestamp 1644511149
transform 1 0 24472 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0840_
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0841_
timestamp 1644511149
transform 1 0 23552 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0842_
timestamp 1644511149
transform 1 0 23184 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0843_
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1644511149
transform 1 0 23828 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0845_
timestamp 1644511149
transform 1 0 25024 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0847_
timestamp 1644511149
transform 1 0 20976 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0848_
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0849_
timestamp 1644511149
transform 1 0 21896 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0850_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0851_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0852_
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0853_
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0854_
timestamp 1644511149
transform 1 0 21988 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0855_
timestamp 1644511149
transform 1 0 21988 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0856_
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0857_
timestamp 1644511149
transform 1 0 23092 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0858_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0859_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1644511149
transform 1 0 33764 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0861_
timestamp 1644511149
transform 1 0 31372 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 1644511149
transform 1 0 30820 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32200 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0864_
timestamp 1644511149
transform 1 0 33396 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0866_
timestamp 1644511149
transform 1 0 29624 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0867_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0868_
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0869_
timestamp 1644511149
transform 1 0 31280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0870_
timestamp 1644511149
transform 1 0 31556 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0872_
timestamp 1644511149
transform 1 0 32016 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1644511149
transform 1 0 31004 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0874_
timestamp 1644511149
transform 1 0 32108 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0875_
timestamp 1644511149
transform 1 0 31188 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0876_
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0877_
timestamp 1644511149
transform 1 0 32384 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0878_
timestamp 1644511149
transform 1 0 33304 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0879_
timestamp 1644511149
transform 1 0 32752 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0880_
timestamp 1644511149
transform 1 0 31648 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0881_
timestamp 1644511149
transform 1 0 33764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0883_
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1644511149
transform 1 0 30728 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1644511149
transform 1 0 31004 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1644511149
transform 1 0 30360 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0887_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0889_
timestamp 1644511149
transform 1 0 33856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0890_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 39928 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 43792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 45632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 26036 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 5060 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0908_
timestamp 1644511149
transform 1 0 35052 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 27508 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 46736 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0914_
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _0915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 21620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 45540 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 15640 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0921_
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 11960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 11040 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 12052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0927_
timestamp 1644511149
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0933_
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 22816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 14996 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0939_
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 22448 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0946_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 24748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0952_
timestamp 1644511149
transform 1 0 19228 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0958_
timestamp 1644511149
transform 1 0 19228 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 43516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 43332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 38640 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0964_
timestamp 1644511149
transform 1 0 18216 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 18216 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 19504 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 10488 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 2116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0970_
timestamp 1644511149
transform 1 0 20700 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 17756 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0976_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0977_
timestamp 1644511149
transform 1 0 17664 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 17296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 15088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 17296 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0983_
timestamp 1644511149
transform 1 0 42136 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 39376 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 33672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 46736 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0989_
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 42964 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0995_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1001_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 34408 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1644511149
transform 1 0 23184 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33488 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform 1 0 34592 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35604 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46000 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1015_
timestamp 1644511149
transform 1 0 46368 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1016_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1644511149
transform 1 0 47932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1644511149
transform 1 0 45448 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1020_
timestamp 1644511149
transform 1 0 46184 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _1021_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1644511149
transform 1 0 45632 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1023_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1024_
timestamp 1644511149
transform 1 0 40020 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1026_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1644511149
transform 1 0 39008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1029_
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1644511149
transform 1 0 40664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21620 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _1032_
timestamp 1644511149
transform 1 0 43240 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1644511149
transform 1 0 44068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1644511149
transform 1 0 44068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1035_
timestamp 1644511149
transform 1 0 42872 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1036_
timestamp 1644511149
transform 1 0 44160 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1644511149
transform 1 0 45632 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1644511149
transform 1 0 27140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 1644511149
transform 1 0 27784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1040_
timestamp 1644511149
transform 1 0 28704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 1644511149
transform 1 0 27140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1042_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1043_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1044_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1045_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43516 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1644511149
transform 1 0 43148 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1047_
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43332 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1049_
timestamp 1644511149
transform 1 0 43332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1644511149
transform 1 0 44528 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1644511149
transform 1 0 42504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1052_
timestamp 1644511149
transform 1 0 42964 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 1644511149
transform 1 0 43884 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1644511149
transform 1 0 44068 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44160 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1056_
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1057_
timestamp 1644511149
transform 1 0 43608 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1058_
timestamp 1644511149
transform 1 0 29072 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 28428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1060_
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1061_
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1644511149
transform 1 0 29624 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1064_
timestamp 1644511149
transform 1 0 30452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1065_
timestamp 1644511149
transform 1 0 29992 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 1644511149
transform 1 0 30820 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1644511149
transform 1 0 43332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1071_
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1072_
timestamp 1644511149
transform 1 0 40480 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1073_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1644511149
transform 1 0 33028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1075_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1077_
timestamp 1644511149
transform 1 0 2668 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1079_
timestamp 1644511149
transform 1 0 46276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1081_
timestamp 1644511149
transform -1 0 34500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1083_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1085_
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1644511149
transform 1 0 44252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1087_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1644511149
transform 1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1089_
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 32844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1093_
timestamp 1644511149
transform 1 0 28152 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1644511149
transform 1 0 33212 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 33488 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 34684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1099_
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1644511149
transform 1 0 19504 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1644511149
transform 1 0 19320 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 19780 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1644511149
transform 1 0 24564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1644511149
transform 1 0 28428 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 25576 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1644511149
transform 1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 28244 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 29992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1111_
timestamp 1644511149
transform 1 0 24472 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 30728 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1644511149
transform 1 0 32016 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 27876 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 25392 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1117_
timestamp 1644511149
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1644511149
transform 1 0 20700 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1644511149
transform 1 0 19872 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1644511149
transform 1 0 19136 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 19688 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1123_
timestamp 1644511149
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1644511149
transform 1 0 23184 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1128_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1129_
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1130_
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1132_
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1133_
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1134_
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1135_
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1136_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1644511149
transform 1 0 15088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1138_
timestamp 1644511149
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1644511149
transform 1 0 13248 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1141_
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1142_
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1143_
timestamp 1644511149
transform 1 0 10488 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1144_
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1145_
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1146_
timestamp 1644511149
transform 1 0 10120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1147_
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1644511149
transform 1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1149_
timestamp 1644511149
transform 1 0 10304 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1150_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1152_
timestamp 1644511149
transform 1 0 12512 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1153_
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1154_
timestamp 1644511149
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1155_
timestamp 1644511149
transform 1 0 17296 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1156_
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1644511149
transform 1 0 18308 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1158_
timestamp 1644511149
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1159_
timestamp 1644511149
transform 1 0 19412 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1160_
timestamp 1644511149
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1161_
timestamp 1644511149
transform 1 0 23828 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1162_
timestamp 1644511149
transform 1 0 28152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1163_
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1644511149
transform 1 0 23460 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1644511149
transform 1 0 30728 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1644511149
transform 1 0 32384 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1644511149
transform 1 0 33948 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1644511149
transform 1 0 32292 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1644511149
transform 1 0 28520 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1644511149
transform 1 0 18584 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1644511149
transform 1 0 23276 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1644511149
transform 1 0 24656 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1644511149
transform 1 0 26036 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1644511149
transform 1 0 29532 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1644511149
transform 1 0 27232 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1644511149
transform 1 0 22080 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1644511149
transform 1 0 19136 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1644511149
transform 1 0 18952 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1644511149
transform 1 0 24656 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1198_
timestamp 1644511149
transform 1 0 26772 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1199_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1200_
timestamp 1644511149
transform 1 0 23184 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1201_
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1644511149
transform 1 0 21252 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1203_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1204_
timestamp 1644511149
transform 1 0 19228 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1644511149
transform 1 0 16836 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1206_
timestamp 1644511149
transform 1 0 14536 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1210_
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1644511149
transform 1 0 9476 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1215_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1216_
timestamp 1644511149
transform 1 0 10580 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1644511149
transform 1 0 13248 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1644511149
transform 1 0 16652 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1222_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1223_
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 1644511149
transform 1 0 22264 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1226_
timestamp 1644511149
transform 1 0 24472 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1228_
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1644511149
transform 1 0 28704 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1230_
timestamp 1644511149
transform 1 0 21988 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1231__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1232__82
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1233__83
timestamp 1644511149
transform 1 0 17572 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1234__84
timestamp 1644511149
transform 1 0 47472 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1235__85
timestamp 1644511149
transform 1 0 47472 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1236__86
timestamp 1644511149
transform 1 0 20516 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1237__87
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1238__88
timestamp 1644511149
transform 1 0 25300 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1239__89
timestamp 1644511149
transform 1 0 10488 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1240__90
timestamp 1644511149
transform 1 0 26128 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1241__91
timestamp 1644511149
transform 1 0 47472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1242__92
timestamp 1644511149
transform 1 0 2668 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1243__93
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1244__94
timestamp 1644511149
transform 1 0 4232 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1245__95
timestamp 1644511149
transform 1 0 1472 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1246__96
timestamp 1644511149
transform 1 0 43792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1247__97
timestamp 1644511149
transform 1 0 46368 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1248__98
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1249__99
timestamp 1644511149
transform 1 0 47840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1250__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1251__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1252__102
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1253__103
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1254__104
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1255__105
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1256__106
timestamp 1644511149
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1257__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1258__108
timestamp 1644511149
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1259__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1260__110
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1261__111
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1262__112
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1263__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1264__114
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1265__115
timestamp 1644511149
transform 1 0 25392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1266__116
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1267__117
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1268__118
timestamp 1644511149
transform 1 0 12972 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1269__119
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1270__120
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1271__121
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1272__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1273__123
timestamp 1644511149
transform 1 0 46644 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1274__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1275__125
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1276__126
timestamp 1644511149
transform 1 0 18768 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1277__127
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1278__128
timestamp 1644511149
transform 1 0 47472 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1279__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1280__130
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1281__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1282__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1283__133
timestamp 1644511149
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1284__134
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1285__135
timestamp 1644511149
transform 1 0 44252 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31280 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 31188 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 43608 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 44436 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 45172 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 43332 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 38548 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 18308 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 20148 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 10488 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 10396 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 42780 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1315_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1316_
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1317_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1318_
timestamp 1644511149
transform 1 0 35052 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1319_
timestamp 1644511149
transform 1 0 30820 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1320_
timestamp 1644511149
transform 1 0 11684 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1321_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1322_
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1323_
timestamp 1644511149
transform 1 0 19412 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1324_
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1325_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1326_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1327_
timestamp 1644511149
transform 1 0 16744 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1328_
timestamp 1644511149
transform 1 0 16836 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1329_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1330_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1331_
timestamp 1644511149
transform 1 0 14260 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1332_
timestamp 1644511149
transform 1 0 8188 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1333_
timestamp 1644511149
transform 1 0 11776 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1334_
timestamp 1644511149
transform 1 0 14720 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1335_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1336_
timestamp 1644511149
transform 1 0 8280 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1337_
timestamp 1644511149
transform 1 0 14260 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1338_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1339_
timestamp 1644511149
transform 1 0 16836 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1340_
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1341_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1342_
timestamp 1644511149
transform 1 0 16376 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1343_
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1344_
timestamp 1644511149
transform 1 0 19412 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1345_
timestamp 1644511149
transform 1 0 23276 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1346_
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 32752 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 30176 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 9108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 21896 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 13616 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 6532 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 46276 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1372_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1373_
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1374_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1375_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1376_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1377_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1378_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1379_
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1380_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1381_
timestamp 1644511149
transform 1 0 44160 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27324 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 24840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 29532 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 23092 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 47288 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 45540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1644511149
transform 1 0 46736 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1644511149
transform 1 0 47288 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1644511149
transform 1 0 46184 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1644511149
transform 1 0 12328 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 46460 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 15364 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 45356 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 11592 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46184 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 45632 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 40848 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 39192 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39652 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 15088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 20424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 26036 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2208 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42228 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37536 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 30452 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 26036 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45448 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 34868 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46736 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 38272 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 32292 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 32200 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 34868 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45632 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45540 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 40020 0 -1 22848
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
