magic
tech sky130A
magscale 1 2
timestamp 1654258427
<< viali >>
rect 3065 47209 3099 47243
rect 29929 47209 29963 47243
rect 31033 47209 31067 47243
rect 5089 47141 5123 47175
rect 22477 47141 22511 47175
rect 44097 47141 44131 47175
rect 47961 47141 47995 47175
rect 2053 47073 2087 47107
rect 11713 47073 11747 47107
rect 11989 47073 12023 47107
rect 14105 47073 14139 47107
rect 14381 47073 14415 47107
rect 47041 47073 47075 47107
rect 1777 47005 1811 47039
rect 3801 47005 3835 47039
rect 4813 47005 4847 47039
rect 6377 47005 6411 47039
rect 7389 47005 7423 47039
rect 9413 47005 9447 47039
rect 13001 47005 13035 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 21097 47005 21131 47039
rect 22017 47005 22051 47039
rect 22661 47005 22695 47039
rect 24777 47005 24811 47039
rect 25513 47005 25547 47039
rect 28549 47005 28583 47039
rect 29745 47005 29779 47039
rect 31217 47005 31251 47039
rect 38393 47005 38427 47039
rect 42717 47005 42751 47039
rect 43269 47005 43303 47039
rect 43913 47005 43947 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 2789 46937 2823 46971
rect 4077 46937 4111 46971
rect 6653 46937 6687 46971
rect 7573 46937 7607 46971
rect 9597 46937 9631 46971
rect 19717 46937 19751 46971
rect 20085 46937 20119 46971
rect 28733 46937 28767 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 43453 46937 43487 46971
rect 45385 46937 45419 46971
rect 13185 46869 13219 46903
rect 5825 46597 5859 46631
rect 1409 46529 1443 46563
rect 19441 46529 19475 46563
rect 24593 46529 24627 46563
rect 38117 46529 38151 46563
rect 47961 46529 47995 46563
rect 3985 46461 4019 46495
rect 4169 46461 4203 46495
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 12173 46461 12207 46495
rect 13829 46461 13863 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 31585 46461 31619 46495
rect 32137 46461 32171 46495
rect 32321 46461 32355 46495
rect 32597 46461 32631 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46765 46461 46799 46495
rect 1593 46325 1627 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 4353 46121 4387 46155
rect 5089 46121 5123 46155
rect 13553 46121 13587 46155
rect 14197 46121 14231 46155
rect 20085 46121 20119 46155
rect 24685 46121 24719 46155
rect 31861 46121 31895 46155
rect 38301 46121 38335 46155
rect 43729 46121 43763 46155
rect 44373 46121 44407 46155
rect 20821 45985 20855 46019
rect 21281 45985 21315 46019
rect 25237 45985 25271 46019
rect 25789 45985 25823 46019
rect 41337 45985 41371 46019
rect 41889 45985 41923 46019
rect 47041 45985 47075 46019
rect 2053 45917 2087 45951
rect 4997 45917 5031 45951
rect 12541 45917 12575 45951
rect 14105 45917 14139 45951
rect 19993 45917 20027 45951
rect 24593 45917 24627 45951
rect 31769 45917 31803 45951
rect 38209 45917 38243 45951
rect 43637 45917 43671 45951
rect 44281 45917 44315 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 21005 45849 21039 45883
rect 25421 45849 25455 45883
rect 41521 45849 41555 45883
rect 45845 45849 45879 45883
rect 46489 45849 46523 45883
rect 12357 45781 12391 45815
rect 12081 45577 12115 45611
rect 21097 45577 21131 45611
rect 25421 45577 25455 45611
rect 41521 45577 41555 45611
rect 1777 45441 1811 45475
rect 11989 45441 12023 45475
rect 21005 45441 21039 45475
rect 25329 45441 25363 45475
rect 27169 45441 27203 45475
rect 41429 45441 41463 45475
rect 44925 45441 44959 45475
rect 47593 45441 47627 45475
rect 1961 45373 1995 45407
rect 2789 45373 2823 45407
rect 42625 45373 42659 45407
rect 42809 45373 42843 45407
rect 44097 45373 44131 45407
rect 45109 45373 45143 45407
rect 45661 45373 45695 45407
rect 27261 45237 27295 45271
rect 47777 45237 47811 45271
rect 2237 45033 2271 45067
rect 42809 45033 42843 45067
rect 43545 45033 43579 45067
rect 44373 45033 44407 45067
rect 45753 45033 45787 45067
rect 45201 44965 45235 44999
rect 27261 44897 27295 44931
rect 48145 44897 48179 44931
rect 2145 44829 2179 44863
rect 27077 44829 27111 44863
rect 42717 44829 42751 44863
rect 44281 44829 44315 44863
rect 45661 44829 45695 44863
rect 46305 44829 46339 44863
rect 28917 44761 28951 44795
rect 46489 44761 46523 44795
rect 27077 44489 27111 44523
rect 46305 44489 46339 44523
rect 47685 44421 47719 44455
rect 26985 44353 27019 44387
rect 45109 44353 45143 44387
rect 45753 44353 45787 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 46949 44149 46983 44183
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 1409 43265 1443 43299
rect 47041 43265 47075 43299
rect 1685 43197 1719 43231
rect 47777 43061 47811 43095
rect 46305 42721 46339 42755
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 46949 42313 46983 42347
rect 46857 42177 46891 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 47685 41973 47719 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46489 41633 46523 41667
rect 46305 41565 46339 41599
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 2145 41225 2179 41259
rect 2053 41089 2087 41123
rect 47961 41089 47995 41123
rect 48053 40885 48087 40919
rect 47685 40681 47719 40715
rect 22293 40477 22327 40511
rect 1869 40409 1903 40443
rect 1961 40341 1995 40375
rect 22109 40341 22143 40375
rect 22937 40137 22971 40171
rect 20361 40069 20395 40103
rect 20545 40069 20579 40103
rect 22293 40001 22327 40035
rect 22661 40001 22695 40035
rect 23305 40001 23339 40035
rect 24041 40001 24075 40035
rect 23397 39933 23431 39967
rect 23489 39933 23523 39967
rect 20729 39797 20763 39831
rect 47777 39797 47811 39831
rect 21649 39457 21683 39491
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 19901 39389 19935 39423
rect 21373 39389 21407 39423
rect 45017 39389 45051 39423
rect 46489 39321 46523 39355
rect 20085 39253 20119 39287
rect 23121 39253 23155 39287
rect 45109 39253 45143 39287
rect 20269 39049 20303 39083
rect 22017 39049 22051 39083
rect 23121 39049 23155 39083
rect 45201 38981 45235 39015
rect 46857 38981 46891 39015
rect 20085 38913 20119 38947
rect 21925 38913 21959 38947
rect 22753 38913 22787 38947
rect 23581 38913 23615 38947
rect 27813 38913 27847 38947
rect 43637 38913 43671 38947
rect 47777 38913 47811 38947
rect 22661 38845 22695 38879
rect 44373 38845 44407 38879
rect 45017 38845 45051 38879
rect 23673 38709 23707 38743
rect 27905 38709 27939 38743
rect 47869 38709 47903 38743
rect 46949 38505 46983 38539
rect 19533 38369 19567 38403
rect 21925 38369 21959 38403
rect 24409 38369 24443 38403
rect 26617 38369 26651 38403
rect 44281 38369 44315 38403
rect 16313 38301 16347 38335
rect 16497 38301 16531 38335
rect 43545 38301 43579 38335
rect 45017 38301 45051 38335
rect 46857 38301 46891 38335
rect 19809 38233 19843 38267
rect 22201 38233 22235 38267
rect 24685 38233 24719 38267
rect 26893 38233 26927 38267
rect 45937 38233 45971 38267
rect 16405 38165 16439 38199
rect 21281 38165 21315 38199
rect 23673 38165 23707 38199
rect 26157 38165 26191 38199
rect 28365 38165 28399 38199
rect 17601 37961 17635 37995
rect 18705 37961 18739 37995
rect 20637 37961 20671 37995
rect 24777 37961 24811 37995
rect 25605 37961 25639 37995
rect 26985 37961 27019 37995
rect 19717 37893 19751 37927
rect 17417 37825 17451 37859
rect 17703 37815 17737 37849
rect 18153 37825 18187 37859
rect 18337 37825 18371 37859
rect 18429 37825 18463 37859
rect 18567 37825 18601 37859
rect 19613 37815 19647 37849
rect 20005 37825 20039 37859
rect 20545 37825 20579 37859
rect 22845 37825 22879 37859
rect 23121 37825 23155 37859
rect 23765 37825 23799 37859
rect 24961 37825 24995 37859
rect 25513 37825 25547 37859
rect 27169 37825 27203 37859
rect 27261 37825 27295 37859
rect 27537 37825 27571 37859
rect 44097 37825 44131 37859
rect 19831 37757 19865 37791
rect 22937 37757 22971 37791
rect 44465 37757 44499 37791
rect 19993 37689 20027 37723
rect 17233 37621 17267 37655
rect 22845 37621 22879 37655
rect 23305 37621 23339 37655
rect 23857 37621 23891 37655
rect 27445 37621 27479 37655
rect 47777 37621 47811 37655
rect 15945 37417 15979 37451
rect 20913 37417 20947 37451
rect 23305 37417 23339 37451
rect 24961 37417 24995 37451
rect 26893 37417 26927 37451
rect 44281 37417 44315 37451
rect 20821 37349 20855 37383
rect 24869 37349 24903 37383
rect 16865 37281 16899 37315
rect 21005 37281 21039 37315
rect 26525 37281 26559 37315
rect 45385 37281 45419 37315
rect 48145 37281 48179 37315
rect 2053 37213 2087 37247
rect 15669 37213 15703 37247
rect 15761 37213 15795 37247
rect 16037 37213 16071 37247
rect 16589 37213 16623 37247
rect 19257 37213 19291 37247
rect 20729 37213 20763 37247
rect 22845 37213 22879 37247
rect 23213 37213 23247 37247
rect 23397 37213 23431 37247
rect 26709 37213 26743 37247
rect 27353 37213 27387 37247
rect 27537 37213 27571 37247
rect 28825 37213 28859 37247
rect 44097 37213 44131 37247
rect 45109 37213 45143 37247
rect 46305 37213 46339 37247
rect 19349 37145 19383 37179
rect 24501 37145 24535 37179
rect 46489 37145 46523 37179
rect 15485 37077 15519 37111
rect 18337 37077 18371 37111
rect 23029 37077 23063 37111
rect 27721 37077 27755 37111
rect 28917 37077 28951 37111
rect 18153 36873 18187 36907
rect 22661 36873 22695 36907
rect 24133 36873 24167 36907
rect 27077 36873 27111 36907
rect 27261 36873 27295 36907
rect 47685 36873 47719 36907
rect 16773 36805 16807 36839
rect 23765 36805 23799 36839
rect 23981 36805 24015 36839
rect 1777 36737 1811 36771
rect 16681 36737 16715 36771
rect 17785 36737 17819 36771
rect 22845 36737 22879 36771
rect 23029 36737 23063 36771
rect 23121 36737 23155 36771
rect 24961 36737 24995 36771
rect 27202 36737 27236 36771
rect 28457 36737 28491 36771
rect 47593 36737 47627 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 13921 36669 13955 36703
rect 14197 36669 14231 36703
rect 17877 36669 17911 36703
rect 27721 36669 27755 36703
rect 28733 36669 28767 36703
rect 15669 36533 15703 36567
rect 23949 36533 23983 36567
rect 25145 36533 25179 36567
rect 27629 36533 27663 36567
rect 30205 36533 30239 36567
rect 2237 36329 2271 36363
rect 15669 36329 15703 36363
rect 22845 36329 22879 36363
rect 25053 36329 25087 36363
rect 25513 36329 25547 36363
rect 27077 36329 27111 36363
rect 15209 36261 15243 36295
rect 16037 36261 16071 36295
rect 14933 36193 14967 36227
rect 24777 36193 24811 36227
rect 24869 36193 24903 36227
rect 25973 36193 26007 36227
rect 2145 36125 2179 36159
rect 14841 36125 14875 36159
rect 15853 36125 15887 36159
rect 16129 36125 16163 36159
rect 20545 36125 20579 36159
rect 22017 36125 22051 36159
rect 23029 36125 23063 36159
rect 23213 36125 23247 36159
rect 23489 36125 23523 36159
rect 24409 36125 24443 36159
rect 25697 36125 25731 36159
rect 25789 36125 25823 36159
rect 26065 36125 26099 36159
rect 26985 36125 27019 36159
rect 27077 36125 27111 36159
rect 27905 36125 27939 36159
rect 27997 36125 28031 36159
rect 28181 36125 28215 36159
rect 28273 36125 28307 36159
rect 22201 36057 22235 36091
rect 23121 36057 23155 36091
rect 23331 36057 23365 36091
rect 26801 36057 26835 36091
rect 20637 35989 20671 36023
rect 22385 35989 22419 36023
rect 27261 35989 27295 36023
rect 27721 35989 27755 36023
rect 23397 35785 23431 35819
rect 24133 35785 24167 35819
rect 26341 35785 26375 35819
rect 27353 35785 27387 35819
rect 29285 35785 29319 35819
rect 22937 35717 22971 35751
rect 30021 35717 30055 35751
rect 1593 35649 1627 35683
rect 17141 35649 17175 35683
rect 17969 35649 18003 35683
rect 19533 35649 19567 35683
rect 22293 35649 22327 35683
rect 23213 35649 23247 35683
rect 23857 35649 23891 35683
rect 23949 35649 23983 35683
rect 24777 35649 24811 35683
rect 25513 35649 25547 35683
rect 26249 35649 26283 35683
rect 26433 35649 26467 35683
rect 26985 35649 27019 35683
rect 28549 35649 28583 35683
rect 28733 35649 28767 35683
rect 29101 35649 29135 35683
rect 29837 35649 29871 35683
rect 30113 35649 30147 35683
rect 30205 35649 30239 35683
rect 18153 35581 18187 35615
rect 18245 35581 18279 35615
rect 19809 35581 19843 35615
rect 23029 35581 23063 35615
rect 24133 35581 24167 35615
rect 27077 35581 27111 35615
rect 28825 35581 28859 35615
rect 28917 35581 28951 35615
rect 25697 35513 25731 35547
rect 1409 35445 1443 35479
rect 17233 35445 17267 35479
rect 17785 35445 17819 35479
rect 21281 35445 21315 35479
rect 22385 35445 22419 35479
rect 23029 35445 23063 35479
rect 24869 35445 24903 35479
rect 26985 35445 27019 35479
rect 30389 35445 30423 35479
rect 20637 35241 20671 35275
rect 21097 35241 21131 35275
rect 22385 35241 22419 35275
rect 26157 35173 26191 35207
rect 27537 35173 27571 35207
rect 16773 35105 16807 35139
rect 21189 35105 21223 35139
rect 22017 35105 22051 35139
rect 22477 35105 22511 35139
rect 26801 35105 26835 35139
rect 26985 35105 27019 35139
rect 30389 35105 30423 35139
rect 19889 35037 19923 35071
rect 20085 35035 20119 35069
rect 20177 35037 20211 35071
rect 20269 35037 20303 35071
rect 20464 35037 20498 35071
rect 21373 35037 21407 35071
rect 22201 35037 22235 35071
rect 24409 35037 24443 35071
rect 25789 35037 25823 35071
rect 25973 35037 26007 35071
rect 26249 35037 26283 35071
rect 26709 35037 26743 35071
rect 27445 35037 27479 35071
rect 27629 35037 27663 35071
rect 48145 35037 48179 35071
rect 17049 34969 17083 35003
rect 21097 34969 21131 35003
rect 26985 34969 27019 35003
rect 30665 34969 30699 35003
rect 18521 34901 18555 34935
rect 21557 34901 21591 34935
rect 24593 34901 24627 34935
rect 32137 34901 32171 34935
rect 47961 34901 47995 34935
rect 17969 34697 18003 34731
rect 22845 34697 22879 34731
rect 23397 34697 23431 34731
rect 24041 34697 24075 34731
rect 25881 34697 25915 34731
rect 30757 34697 30791 34731
rect 32229 34697 32263 34731
rect 14289 34629 14323 34663
rect 18429 34629 18463 34663
rect 22753 34629 22787 34663
rect 31125 34629 31159 34663
rect 14197 34561 14231 34595
rect 15025 34561 15059 34595
rect 15117 34561 15151 34595
rect 15393 34561 15427 34595
rect 17233 34561 17267 34595
rect 17417 34561 17451 34595
rect 17601 34561 17635 34595
rect 17785 34561 17819 34595
rect 18613 34561 18647 34595
rect 19625 34561 19659 34595
rect 20361 34561 20395 34595
rect 21833 34561 21867 34595
rect 22017 34561 22051 34595
rect 22201 34561 22235 34595
rect 26065 34561 26099 34595
rect 26157 34561 26191 34595
rect 26433 34561 26467 34595
rect 29929 34561 29963 34595
rect 30941 34561 30975 34595
rect 31217 34561 31251 34595
rect 32137 34561 32171 34595
rect 48145 34561 48179 34595
rect 15301 34493 15335 34527
rect 17509 34493 17543 34527
rect 20637 34493 20671 34527
rect 24133 34493 24167 34527
rect 24317 34493 24351 34527
rect 29837 34493 29871 34527
rect 30297 34425 30331 34459
rect 14841 34357 14875 34391
rect 18797 34357 18831 34391
rect 19809 34357 19843 34391
rect 20637 34357 20671 34391
rect 20913 34357 20947 34391
rect 23673 34357 23707 34391
rect 26341 34357 26375 34391
rect 47961 34357 47995 34391
rect 17601 34153 17635 34187
rect 20637 34153 20671 34187
rect 27261 34153 27295 34187
rect 48053 34153 48087 34187
rect 17877 34085 17911 34119
rect 14105 34017 14139 34051
rect 21189 34017 21223 34051
rect 1593 33949 1627 33983
rect 16313 33949 16347 33983
rect 16497 33949 16531 33983
rect 17325 33949 17359 33983
rect 17693 33949 17727 33983
rect 20453 33949 20487 33983
rect 21465 33949 21499 33983
rect 23213 33949 23247 33983
rect 23673 33949 23707 33983
rect 24409 33949 24443 33983
rect 25513 33949 25547 33983
rect 27813 33949 27847 33983
rect 30389 33949 30423 33983
rect 31033 33949 31067 33983
rect 14381 33881 14415 33915
rect 25789 33881 25823 33915
rect 30205 33881 30239 33915
rect 47961 33881 47995 33915
rect 1409 33813 1443 33847
rect 15853 33813 15887 33847
rect 16405 33813 16439 33847
rect 23029 33813 23063 33847
rect 23765 33813 23799 33847
rect 24593 33813 24627 33847
rect 27997 33813 28031 33847
rect 30573 33813 30607 33847
rect 31125 33813 31159 33847
rect 13921 33609 13955 33643
rect 14381 33609 14415 33643
rect 18337 33609 18371 33643
rect 26341 33609 26375 33643
rect 27629 33609 27663 33643
rect 28825 33609 28859 33643
rect 21097 33541 21131 33575
rect 22477 33541 22511 33575
rect 24961 33541 24995 33575
rect 30113 33541 30147 33575
rect 13645 33473 13679 33507
rect 14565 33473 14599 33507
rect 14749 33473 14783 33507
rect 14841 33473 14875 33507
rect 15853 33473 15887 33507
rect 16865 33473 16899 33507
rect 17877 33473 17911 33507
rect 18153 33473 18187 33507
rect 22201 33473 22235 33507
rect 25605 33473 25639 33507
rect 26249 33473 26283 33507
rect 27537 33473 27571 33507
rect 28181 33473 28215 33507
rect 28328 33473 28362 33507
rect 29377 33473 29411 33507
rect 29653 33473 29687 33507
rect 30573 33473 30607 33507
rect 32137 33473 32171 33507
rect 47041 33473 47075 33507
rect 47593 33473 47627 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 13921 33405 13955 33439
rect 16037 33405 16071 33439
rect 16129 33405 16163 33439
rect 17141 33405 17175 33439
rect 18061 33405 18095 33439
rect 28549 33405 28583 33439
rect 30849 33405 30883 33439
rect 30941 33405 30975 33439
rect 32413 33405 32447 33439
rect 48053 33405 48087 33439
rect 15669 33337 15703 33371
rect 25697 33337 25731 33371
rect 28457 33337 28491 33371
rect 29469 33337 29503 33371
rect 13737 33269 13771 33303
rect 17049 33269 17083 33303
rect 17417 33269 17451 33303
rect 17877 33269 17911 33303
rect 21189 33269 21223 33303
rect 23949 33269 23983 33303
rect 25053 33269 25087 33303
rect 30665 33269 30699 33303
rect 31033 33269 31067 33303
rect 33885 33269 33919 33303
rect 46857 33269 46891 33303
rect 47869 33269 47903 33303
rect 1961 33065 1995 33099
rect 14473 33065 14507 33099
rect 15301 33065 15335 33099
rect 16497 33065 16531 33099
rect 16681 33065 16715 33099
rect 26065 33065 26099 33099
rect 32229 33065 32263 33099
rect 32965 33065 32999 33099
rect 14841 32997 14875 33031
rect 23673 32997 23707 33031
rect 2329 32929 2363 32963
rect 14565 32929 14599 32963
rect 23397 32929 23431 32963
rect 29929 32929 29963 32963
rect 31769 32929 31803 32963
rect 47133 32929 47167 32963
rect 47685 32929 47719 32963
rect 1869 32861 1903 32895
rect 2973 32861 3007 32895
rect 14473 32861 14507 32895
rect 15301 32861 15335 32895
rect 15485 32861 15519 32895
rect 15577 32861 15611 32895
rect 16405 32861 16439 32895
rect 16497 32861 16531 32895
rect 17141 32861 17175 32895
rect 17325 32861 17359 32895
rect 17417 32861 17451 32895
rect 17509 32861 17543 32895
rect 17693 32861 17727 32895
rect 18521 32861 18555 32895
rect 19993 32861 20027 32895
rect 22201 32861 22235 32895
rect 23305 32861 23339 32895
rect 27077 32861 27111 32895
rect 29653 32861 29687 32895
rect 31493 32861 31527 32895
rect 31677 32861 31711 32895
rect 31861 32861 31895 32895
rect 32045 32861 32079 32895
rect 32873 32861 32907 32895
rect 46581 32861 46615 32895
rect 16221 32793 16255 32827
rect 20269 32793 20303 32827
rect 22293 32793 22327 32827
rect 24777 32793 24811 32827
rect 27261 32793 27295 32827
rect 47225 32793 47259 32827
rect 2789 32725 2823 32759
rect 15761 32725 15795 32759
rect 17877 32725 17911 32759
rect 18613 32725 18647 32759
rect 21741 32725 21775 32759
rect 17049 32521 17083 32555
rect 19257 32521 19291 32555
rect 21281 32521 21315 32555
rect 24241 32521 24275 32555
rect 24409 32521 24443 32555
rect 29561 32521 29595 32555
rect 48053 32521 48087 32555
rect 2237 32453 2271 32487
rect 16865 32453 16899 32487
rect 17785 32453 17819 32487
rect 24041 32453 24075 32487
rect 29193 32453 29227 32487
rect 2053 32385 2087 32419
rect 16681 32385 16715 32419
rect 20545 32385 20579 32419
rect 20729 32385 20763 32419
rect 21097 32385 21131 32419
rect 24961 32385 24995 32419
rect 25789 32385 25823 32419
rect 26985 32385 27019 32419
rect 29377 32385 29411 32419
rect 30021 32385 30055 32419
rect 30113 32385 30147 32419
rect 32137 32385 32171 32419
rect 46857 32385 46891 32419
rect 47961 32385 47995 32419
rect 3893 32317 3927 32351
rect 17509 32317 17543 32351
rect 20821 32317 20855 32351
rect 20913 32317 20947 32351
rect 25697 32317 25731 32351
rect 27261 32317 27295 32351
rect 28733 32317 28767 32351
rect 32413 32317 32447 32351
rect 25145 32249 25179 32283
rect 1593 32181 1627 32215
rect 24225 32181 24259 32215
rect 26157 32181 26191 32215
rect 30113 32181 30147 32215
rect 30389 32181 30423 32215
rect 33885 32181 33919 32215
rect 46949 32181 46983 32215
rect 19901 31977 19935 32011
rect 23305 31977 23339 32011
rect 23489 31977 23523 32011
rect 25789 31977 25823 32011
rect 26801 31977 26835 32011
rect 28825 31977 28859 32011
rect 30297 31977 30331 32011
rect 32229 31977 32263 32011
rect 32873 31977 32907 32011
rect 17049 31909 17083 31943
rect 21005 31909 21039 31943
rect 27813 31909 27847 31943
rect 30573 31909 30607 31943
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 14381 31841 14415 31875
rect 14657 31841 14691 31875
rect 15853 31841 15887 31875
rect 20545 31841 20579 31875
rect 24777 31841 24811 31875
rect 27261 31841 27295 31875
rect 28273 31841 28307 31875
rect 31769 31841 31803 31875
rect 31861 31841 31895 31875
rect 46305 31841 46339 31875
rect 46489 31841 46523 31875
rect 48145 31841 48179 31875
rect 14289 31773 14323 31807
rect 15669 31773 15703 31807
rect 17049 31773 17083 31807
rect 17233 31773 17267 31807
rect 17693 31773 17727 31807
rect 17785 31773 17819 31807
rect 19809 31773 19843 31807
rect 20637 31773 20671 31807
rect 24961 31773 24995 31807
rect 25697 31773 25731 31807
rect 26985 31773 27019 31807
rect 27137 31773 27171 31807
rect 27353 31773 27387 31807
rect 27997 31773 28031 31807
rect 28089 31773 28123 31807
rect 28365 31773 28399 31807
rect 28825 31773 28859 31807
rect 29009 31773 29043 31807
rect 30021 31773 30055 31807
rect 30297 31773 30331 31807
rect 31493 31773 31527 31807
rect 31677 31773 31711 31807
rect 32045 31773 32079 31807
rect 32781 31773 32815 31807
rect 23351 31739 23385 31773
rect 1593 31705 1627 31739
rect 23121 31705 23155 31739
rect 25237 31705 25271 31739
rect 25145 31637 25179 31671
rect 2237 31433 2271 31467
rect 15577 31433 15611 31467
rect 24777 31433 24811 31467
rect 28917 31433 28951 31467
rect 30573 31433 30607 31467
rect 3065 31365 3099 31399
rect 4721 31365 4755 31399
rect 20729 31365 20763 31399
rect 29929 31365 29963 31399
rect 2145 31297 2179 31331
rect 17049 31297 17083 31331
rect 17877 31297 17911 31331
rect 20085 31297 20119 31331
rect 20913 31297 20947 31331
rect 23581 31297 23615 31331
rect 24593 31297 24627 31331
rect 25789 31297 25823 31331
rect 25973 31297 26007 31331
rect 27537 31297 27571 31331
rect 28641 31297 28675 31331
rect 28733 31297 28767 31331
rect 29653 31297 29687 31331
rect 29745 31297 29779 31331
rect 30389 31297 30423 31331
rect 30665 31297 30699 31331
rect 32137 31297 32171 31331
rect 2881 31229 2915 31263
rect 13829 31229 13863 31263
rect 14105 31229 14139 31263
rect 16865 31229 16899 31263
rect 23305 31229 23339 31263
rect 29929 31229 29963 31263
rect 17233 31093 17267 31127
rect 18061 31093 18095 31127
rect 20177 31093 20211 31127
rect 21097 31093 21131 31127
rect 25789 31093 25823 31127
rect 27721 31093 27755 31127
rect 30389 31093 30423 31127
rect 32229 31093 32263 31127
rect 15117 30889 15151 30923
rect 15669 30889 15703 30923
rect 17325 30889 17359 30923
rect 18521 30889 18555 30923
rect 21833 30889 21867 30923
rect 24777 30889 24811 30923
rect 28917 30889 28951 30923
rect 32597 30889 32631 30923
rect 24961 30821 24995 30855
rect 19257 30753 19291 30787
rect 19533 30753 19567 30787
rect 21925 30753 21959 30787
rect 25421 30753 25455 30787
rect 27997 30753 28031 30787
rect 30849 30753 30883 30787
rect 47133 30753 47167 30787
rect 14473 30685 14507 30719
rect 14566 30685 14600 30719
rect 14979 30685 15013 30719
rect 15577 30685 15611 30719
rect 17141 30685 17175 30719
rect 17417 30685 17451 30719
rect 18337 30685 18371 30719
rect 21649 30685 21683 30719
rect 22569 30685 22603 30719
rect 23581 30685 23615 30719
rect 24409 30685 24443 30719
rect 24777 30685 24811 30719
rect 27813 30685 27847 30719
rect 28733 30685 28767 30719
rect 29745 30685 29779 30719
rect 29837 30685 29871 30719
rect 30021 30685 30055 30719
rect 30113 30685 30147 30719
rect 14749 30617 14783 30651
rect 14841 30617 14875 30651
rect 25697 30617 25731 30651
rect 31125 30617 31159 30651
rect 46857 30617 46891 30651
rect 46949 30617 46983 30651
rect 16957 30549 16991 30583
rect 21005 30549 21039 30583
rect 21465 30549 21499 30583
rect 22661 30549 22695 30583
rect 23765 30549 23799 30583
rect 27169 30549 27203 30583
rect 29561 30549 29595 30583
rect 14657 30345 14691 30379
rect 18429 30345 18463 30379
rect 20637 30345 20671 30379
rect 26341 30345 26375 30379
rect 20361 30277 20395 30311
rect 24317 30277 24351 30311
rect 27077 30277 27111 30311
rect 28181 30277 28215 30311
rect 29469 30277 29503 30311
rect 14565 30209 14599 30243
rect 14749 30209 14783 30243
rect 19349 30209 19383 30243
rect 19533 30209 19567 30243
rect 19993 30209 20027 30243
rect 20086 30209 20120 30243
rect 20269 30209 20303 30243
rect 20499 30209 20533 30243
rect 21097 30209 21131 30243
rect 21281 30209 21315 30243
rect 24501 30209 24535 30243
rect 25697 30209 25731 30243
rect 25845 30209 25879 30243
rect 25973 30209 26007 30243
rect 26065 30209 26099 30243
rect 26203 30209 26237 30243
rect 26985 30209 27019 30243
rect 28089 30209 28123 30243
rect 29653 30209 29687 30243
rect 29929 30209 29963 30243
rect 32965 30209 32999 30243
rect 16681 30141 16715 30175
rect 16957 30141 16991 30175
rect 19441 30141 19475 30175
rect 22017 30141 22051 30175
rect 22293 30141 22327 30175
rect 33149 30141 33183 30175
rect 33425 30141 33459 30175
rect 21189 30005 21223 30039
rect 23765 30005 23799 30039
rect 29837 30005 29871 30039
rect 16681 29801 16715 29835
rect 20453 29801 20487 29835
rect 21465 29801 21499 29835
rect 22845 29801 22879 29835
rect 24593 29801 24627 29835
rect 29653 29801 29687 29835
rect 30021 29801 30055 29835
rect 33149 29801 33183 29835
rect 28825 29733 28859 29767
rect 21373 29665 21407 29699
rect 22385 29665 22419 29699
rect 29653 29665 29687 29699
rect 16037 29597 16071 29631
rect 16185 29597 16219 29631
rect 16313 29597 16347 29631
rect 16502 29597 16536 29631
rect 17233 29597 17267 29631
rect 17325 29597 17359 29631
rect 20269 29597 20303 29631
rect 20453 29597 20487 29631
rect 21097 29597 21131 29631
rect 22109 29597 22143 29631
rect 22293 29597 22327 29631
rect 22477 29597 22511 29631
rect 22661 29597 22695 29631
rect 24409 29597 24443 29631
rect 25145 29597 25179 29631
rect 29837 29597 29871 29631
rect 30665 29597 30699 29631
rect 30849 29597 30883 29631
rect 30941 29597 30975 29631
rect 33057 29597 33091 29631
rect 48145 29597 48179 29631
rect 16405 29529 16439 29563
rect 28641 29529 28675 29563
rect 29561 29529 29595 29563
rect 17509 29461 17543 29495
rect 20637 29461 20671 29495
rect 21649 29461 21683 29495
rect 25329 29461 25363 29495
rect 30481 29461 30515 29495
rect 47961 29461 47995 29495
rect 25973 29257 26007 29291
rect 27353 29257 27387 29291
rect 29837 29257 29871 29291
rect 30297 29257 30331 29291
rect 17601 29189 17635 29223
rect 17325 29121 17359 29155
rect 17418 29121 17452 29155
rect 17690 29121 17724 29155
rect 17829 29121 17863 29155
rect 19993 29121 20027 29155
rect 20177 29121 20211 29155
rect 20361 29121 20395 29155
rect 25789 29121 25823 29155
rect 26065 29121 26099 29155
rect 28365 29121 28399 29155
rect 28549 29121 28583 29155
rect 29285 29121 29319 29155
rect 29469 29121 29503 29155
rect 29561 29121 29595 29155
rect 29653 29121 29687 29155
rect 30481 29121 30515 29155
rect 27445 29053 27479 29087
rect 27629 29053 27663 29087
rect 30757 29053 30791 29087
rect 32321 29053 32355 29087
rect 32505 29053 32539 29087
rect 32781 29053 32815 29087
rect 26985 28985 27019 29019
rect 30665 28985 30699 29019
rect 17969 28917 18003 28951
rect 25605 28917 25639 28951
rect 28457 28917 28491 28951
rect 17509 28713 17543 28747
rect 25973 28713 26007 28747
rect 27353 28713 27387 28747
rect 29009 28713 29043 28747
rect 31309 28713 31343 28747
rect 32505 28713 32539 28747
rect 27905 28645 27939 28679
rect 17325 28577 17359 28611
rect 19625 28577 19659 28611
rect 19717 28577 19751 28611
rect 29561 28577 29595 28611
rect 29837 28577 29871 28611
rect 15025 28509 15059 28543
rect 15669 28509 15703 28543
rect 17233 28509 17267 28543
rect 19349 28509 19383 28543
rect 19521 28511 19555 28545
rect 19901 28509 19935 28543
rect 24869 28509 24903 28543
rect 25881 28509 25915 28543
rect 27169 28509 27203 28543
rect 27905 28509 27939 28543
rect 28181 28509 28215 28543
rect 28641 28509 28675 28543
rect 32413 28509 32447 28543
rect 47685 28509 47719 28543
rect 28825 28441 28859 28475
rect 15117 28373 15151 28407
rect 15761 28373 15795 28407
rect 20085 28373 20119 28407
rect 24961 28373 24995 28407
rect 28089 28373 28123 28407
rect 18797 28169 18831 28203
rect 25881 28169 25915 28203
rect 30573 28169 30607 28203
rect 35633 28169 35667 28203
rect 14473 28101 14507 28135
rect 20545 28101 20579 28135
rect 21833 28101 21867 28135
rect 22017 28101 22051 28135
rect 28641 28101 28675 28135
rect 19441 28033 19475 28067
rect 20177 28033 20211 28067
rect 20361 28033 20395 28067
rect 21005 28033 21039 28067
rect 21189 28033 21223 28067
rect 23351 28033 23385 28067
rect 23486 28033 23520 28067
rect 23581 28036 23615 28070
rect 23765 28033 23799 28067
rect 24225 28033 24259 28067
rect 25421 28033 25455 28067
rect 25605 28033 25639 28067
rect 27445 28033 27479 28067
rect 28457 28033 28491 28067
rect 30205 28033 30239 28067
rect 47593 28033 47627 28067
rect 14289 27965 14323 27999
rect 15853 27965 15887 27999
rect 17049 27965 17083 27999
rect 17325 27965 17359 27999
rect 19717 27965 19751 27999
rect 24317 27965 24351 27999
rect 25973 27965 26007 27999
rect 27629 27965 27663 27999
rect 30297 27965 30331 27999
rect 33885 27965 33919 27999
rect 34161 27965 34195 27999
rect 19625 27897 19659 27931
rect 22201 27897 22235 27931
rect 19257 27829 19291 27863
rect 21005 27829 21039 27863
rect 23121 27829 23155 27863
rect 24225 27829 24259 27863
rect 24593 27829 24627 27863
rect 28825 27829 28859 27863
rect 47685 27829 47719 27863
rect 19441 27625 19475 27659
rect 19809 27625 19843 27659
rect 21281 27625 21315 27659
rect 21373 27625 21407 27659
rect 22017 27625 22051 27659
rect 26138 27625 26172 27659
rect 27629 27625 27663 27659
rect 28733 27625 28767 27659
rect 34161 27625 34195 27659
rect 18613 27557 18647 27591
rect 29837 27557 29871 27591
rect 33057 27557 33091 27591
rect 35081 27557 35115 27591
rect 15117 27489 15151 27523
rect 15853 27489 15887 27523
rect 22109 27489 22143 27523
rect 23489 27489 23523 27523
rect 25881 27489 25915 27523
rect 33885 27489 33919 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 14933 27421 14967 27455
rect 18521 27421 18555 27455
rect 19441 27421 19475 27455
rect 19625 27421 19659 27455
rect 21097 27421 21131 27455
rect 21189 27421 21223 27455
rect 21557 27421 21591 27455
rect 22293 27421 22327 27455
rect 23121 27421 23155 27455
rect 24777 27421 24811 27455
rect 28181 27421 28215 27455
rect 28549 27421 28583 27455
rect 29745 27421 29779 27455
rect 32965 27421 32999 27455
rect 33793 27421 33827 27455
rect 34989 27421 35023 27455
rect 22017 27353 22051 27387
rect 23397 27353 23431 27387
rect 23606 27353 23640 27387
rect 24409 27353 24443 27387
rect 24593 27353 24627 27387
rect 28365 27353 28399 27387
rect 28457 27353 28491 27387
rect 20821 27285 20855 27319
rect 22477 27285 22511 27319
rect 23765 27285 23799 27319
rect 20729 27081 20763 27115
rect 22201 27081 22235 27115
rect 25789 27081 25823 27115
rect 27353 27081 27387 27115
rect 29745 27081 29779 27115
rect 33885 27081 33919 27115
rect 19257 27013 19291 27047
rect 21833 27013 21867 27047
rect 22017 27013 22051 27047
rect 23213 27013 23247 27047
rect 34529 27013 34563 27047
rect 12265 26945 12299 26979
rect 23029 26945 23063 26979
rect 23305 26945 23339 26979
rect 23397 26945 23431 26979
rect 24041 26945 24075 26979
rect 27261 26945 27295 26979
rect 27997 26945 28031 26979
rect 31309 26945 31343 26979
rect 34345 26945 34379 26979
rect 34621 26945 34655 26979
rect 12357 26877 12391 26911
rect 16681 26877 16715 26911
rect 16865 26877 16899 26911
rect 17141 26877 17175 26911
rect 18981 26877 19015 26911
rect 24317 26877 24351 26911
rect 28273 26877 28307 26911
rect 31585 26877 31619 26911
rect 32137 26877 32171 26911
rect 32413 26877 32447 26911
rect 12633 26809 12667 26843
rect 23581 26809 23615 26843
rect 34345 26741 34379 26775
rect 12633 26537 12667 26571
rect 15301 26537 15335 26571
rect 20085 26537 20119 26571
rect 23397 26537 23431 26571
rect 24777 26537 24811 26571
rect 25329 26537 25363 26571
rect 28365 26537 28399 26571
rect 29653 26537 29687 26571
rect 32689 26537 32723 26571
rect 34161 26537 34195 26571
rect 18705 26469 18739 26503
rect 27537 26469 27571 26503
rect 16313 26401 16347 26435
rect 21649 26401 21683 26435
rect 21925 26401 21959 26435
rect 24409 26401 24443 26435
rect 31033 26401 31067 26435
rect 32413 26401 32447 26435
rect 39313 26401 39347 26435
rect 11897 26333 11931 26367
rect 12541 26333 12575 26367
rect 12725 26333 12759 26367
rect 13185 26333 13219 26367
rect 14105 26333 14139 26367
rect 15209 26333 15243 26367
rect 15853 26333 15887 26367
rect 18521 26333 18555 26367
rect 19257 26333 19291 26367
rect 19993 26333 20027 26367
rect 24593 26333 24627 26367
rect 25237 26333 25271 26367
rect 27353 26333 27387 26367
rect 28549 26333 28583 26367
rect 29561 26333 29595 26367
rect 30481 26333 30515 26367
rect 32321 26333 32355 26367
rect 33609 26333 33643 26367
rect 33977 26333 34011 26367
rect 34713 26333 34747 26367
rect 37473 26333 37507 26367
rect 11989 26265 12023 26299
rect 14197 26265 14231 26299
rect 16037 26265 16071 26299
rect 33793 26265 33827 26299
rect 34989 26265 35023 26299
rect 37657 26265 37691 26299
rect 13277 26197 13311 26231
rect 19441 26197 19475 26231
rect 33885 26197 33919 26231
rect 36461 26197 36495 26231
rect 22569 25993 22603 26027
rect 23121 25993 23155 26027
rect 32597 25993 32631 26027
rect 33517 25993 33551 26027
rect 34989 25993 35023 26027
rect 35633 25993 35667 26027
rect 37657 25993 37691 26027
rect 12725 25925 12759 25959
rect 34069 25925 34103 25959
rect 34269 25925 34303 25959
rect 11897 25857 11931 25891
rect 14933 25857 14967 25891
rect 15761 25857 15795 25891
rect 17233 25857 17267 25891
rect 18061 25857 18095 25891
rect 22477 25857 22511 25891
rect 23305 25857 23339 25891
rect 23397 25857 23431 25891
rect 23581 25857 23615 25891
rect 23673 25857 23707 25891
rect 25421 25857 25455 25891
rect 32505 25857 32539 25891
rect 33333 25857 33367 25891
rect 34897 25857 34931 25891
rect 35081 25857 35115 25891
rect 35541 25857 35575 25891
rect 37565 25857 37599 25891
rect 41521 25857 41555 25891
rect 48145 25857 48179 25891
rect 12449 25789 12483 25823
rect 14197 25789 14231 25823
rect 15209 25789 15243 25823
rect 25973 25789 26007 25823
rect 29745 25789 29779 25823
rect 29929 25789 29963 25823
rect 31585 25789 31619 25823
rect 15117 25721 15151 25755
rect 18245 25721 18279 25755
rect 11713 25653 11747 25687
rect 14749 25653 14783 25687
rect 15853 25653 15887 25687
rect 17417 25653 17451 25687
rect 34253 25653 34287 25687
rect 34437 25653 34471 25687
rect 41613 25653 41647 25687
rect 47961 25653 47995 25687
rect 16405 25449 16439 25483
rect 17233 25449 17267 25483
rect 32781 25449 32815 25483
rect 39221 25449 39255 25483
rect 17969 25381 18003 25415
rect 47961 25381 47995 25415
rect 11713 25313 11747 25347
rect 11989 25313 12023 25347
rect 14933 25313 14967 25347
rect 25973 25313 26007 25347
rect 26893 25313 26927 25347
rect 32137 25313 32171 25347
rect 41705 25313 41739 25347
rect 42165 25313 42199 25347
rect 42349 25313 42383 25347
rect 46857 25313 46891 25347
rect 14657 25245 14691 25279
rect 17049 25245 17083 25279
rect 17785 25245 17819 25279
rect 19349 25245 19383 25279
rect 19533 25245 19567 25279
rect 21189 25245 21223 25279
rect 21373 25245 21407 25279
rect 24501 25245 24535 25279
rect 25145 25245 25179 25279
rect 26617 25245 26651 25279
rect 27813 25245 27847 25279
rect 29653 25245 29687 25279
rect 30389 25245 30423 25279
rect 32597 25245 32631 25279
rect 39129 25245 39163 25279
rect 39865 25245 39899 25279
rect 45477 25245 45511 25279
rect 1869 25177 1903 25211
rect 27629 25177 27663 25211
rect 40049 25177 40083 25211
rect 44005 25177 44039 25211
rect 45661 25177 45695 25211
rect 1961 25109 1995 25143
rect 13461 25109 13495 25143
rect 19717 25109 19751 25143
rect 21281 25109 21315 25143
rect 24593 25109 24627 25143
rect 29837 25109 29871 25143
rect 13093 24905 13127 24939
rect 14749 24905 14783 24939
rect 19441 24905 19475 24939
rect 20821 24905 20855 24939
rect 29837 24905 29871 24939
rect 12173 24837 12207 24871
rect 14657 24837 14691 24871
rect 14841 24837 14875 24871
rect 19625 24837 19659 24871
rect 40233 24837 40267 24871
rect 12081 24769 12115 24803
rect 12449 24769 12483 24803
rect 13185 24769 13219 24803
rect 13277 24769 13311 24803
rect 13461 24769 13495 24803
rect 15485 24769 15519 24803
rect 15669 24769 15703 24803
rect 16865 24769 16899 24803
rect 16957 24769 16991 24803
rect 17601 24769 17635 24803
rect 19533 24769 19567 24803
rect 20637 24769 20671 24803
rect 20913 24769 20947 24803
rect 21833 24769 21867 24803
rect 23213 24769 23247 24803
rect 26157 24769 26191 24803
rect 26985 24769 27019 24803
rect 27813 24769 27847 24803
rect 28457 24769 28491 24803
rect 29745 24769 29779 24803
rect 30389 24769 30423 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 34069 24769 34103 24803
rect 34897 24769 34931 24803
rect 38761 24769 38795 24803
rect 39405 24769 39439 24803
rect 39497 24769 39531 24803
rect 44925 24769 44959 24803
rect 45017 24769 45051 24803
rect 47593 24769 47627 24803
rect 12265 24701 12299 24735
rect 15577 24701 15611 24735
rect 23857 24701 23891 24735
rect 24041 24701 24075 24735
rect 25697 24701 25731 24735
rect 31125 24701 31159 24735
rect 34161 24701 34195 24735
rect 34437 24701 34471 24735
rect 35173 24701 35207 24735
rect 36645 24701 36679 24735
rect 40049 24701 40083 24735
rect 41245 24701 41279 24735
rect 12909 24633 12943 24667
rect 14473 24633 14507 24667
rect 19257 24633 19291 24667
rect 20637 24633 20671 24667
rect 23305 24633 23339 24667
rect 12449 24565 12483 24599
rect 15025 24565 15059 24599
rect 17693 24565 17727 24599
rect 19809 24565 19843 24599
rect 21833 24565 21867 24599
rect 26341 24565 26375 24599
rect 26985 24565 27019 24599
rect 27905 24565 27939 24599
rect 28549 24565 28583 24599
rect 32137 24565 32171 24599
rect 38853 24565 38887 24599
rect 47041 24565 47075 24599
rect 47685 24565 47719 24599
rect 12449 24361 12483 24395
rect 15209 24361 15243 24395
rect 20729 24361 20763 24395
rect 32413 24361 32447 24395
rect 34069 24361 34103 24395
rect 35909 24361 35943 24395
rect 13553 24293 13587 24327
rect 33425 24293 33459 24327
rect 35265 24293 35299 24327
rect 21281 24225 21315 24259
rect 21557 24225 21591 24259
rect 25697 24225 25731 24259
rect 28641 24225 28675 24259
rect 38577 24225 38611 24259
rect 39957 24225 39991 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 12449 24157 12483 24191
rect 12633 24157 12667 24191
rect 15117 24157 15151 24191
rect 15945 24157 15979 24191
rect 16957 24157 16991 24191
rect 19717 24157 19751 24191
rect 20453 24157 20487 24191
rect 20545 24157 20579 24191
rect 24593 24157 24627 24191
rect 25789 24157 25823 24191
rect 26617 24157 26651 24191
rect 29653 24157 29687 24191
rect 30481 24157 30515 24191
rect 33149 24157 33183 24191
rect 33241 24157 33275 24191
rect 33977 24157 34011 24191
rect 35173 24157 35207 24191
rect 35817 24157 35851 24191
rect 37013 24157 37047 24191
rect 40049 24157 40083 24191
rect 42993 24157 43027 24191
rect 43177 24157 43211 24191
rect 13369 24089 13403 24123
rect 17233 24089 17267 24123
rect 19349 24089 19383 24123
rect 19625 24089 19659 24123
rect 26893 24089 26927 24123
rect 31217 24089 31251 24123
rect 32229 24089 32263 24123
rect 32445 24089 32479 24123
rect 37197 24089 37231 24123
rect 15945 24021 15979 24055
rect 18705 24021 18739 24055
rect 19533 24021 19567 24055
rect 19901 24021 19935 24055
rect 23029 24021 23063 24055
rect 24685 24021 24719 24055
rect 26157 24021 26191 24055
rect 29745 24021 29779 24055
rect 32597 24021 32631 24055
rect 40417 24021 40451 24055
rect 43085 24021 43119 24055
rect 18429 23817 18463 23851
rect 20361 23817 20395 23851
rect 20545 23817 20579 23851
rect 20729 23817 20763 23851
rect 22845 23817 22879 23851
rect 26341 23817 26375 23851
rect 31407 23817 31441 23851
rect 32781 23817 32815 23851
rect 33149 23817 33183 23851
rect 36093 23817 36127 23851
rect 37381 23817 37415 23851
rect 16037 23749 16071 23783
rect 20177 23749 20211 23783
rect 23949 23749 23983 23783
rect 31309 23749 31343 23783
rect 33793 23749 33827 23783
rect 39037 23749 39071 23783
rect 40693 23749 40727 23783
rect 1869 23681 1903 23715
rect 11897 23681 11931 23715
rect 15117 23681 15151 23715
rect 15945 23681 15979 23715
rect 16681 23681 16715 23715
rect 19073 23681 19107 23715
rect 20453 23681 20487 23715
rect 21833 23681 21867 23715
rect 22753 23681 22787 23715
rect 26341 23681 26375 23715
rect 26985 23681 27019 23715
rect 29653 23681 29687 23715
rect 30665 23681 30699 23715
rect 31493 23681 31527 23715
rect 31585 23681 31619 23715
rect 32873 23681 32907 23715
rect 32965 23681 32999 23715
rect 33609 23681 33643 23715
rect 33885 23681 33919 23715
rect 37289 23681 37323 23715
rect 41337 23681 41371 23715
rect 43177 23681 43211 23715
rect 43545 23681 43579 23715
rect 45937 23681 45971 23715
rect 46121 23681 46155 23715
rect 46581 23681 46615 23715
rect 47593 23681 47627 23715
rect 15209 23613 15243 23647
rect 16957 23613 16991 23647
rect 19165 23613 19199 23647
rect 23673 23613 23707 23647
rect 25697 23613 25731 23647
rect 27261 23613 27295 23647
rect 28733 23613 28767 23647
rect 34345 23613 34379 23647
rect 34621 23613 34655 23647
rect 38853 23613 38887 23647
rect 41245 23613 41279 23647
rect 44649 23613 44683 23647
rect 2053 23545 2087 23579
rect 15485 23545 15519 23579
rect 19441 23545 19475 23579
rect 32597 23545 32631 23579
rect 46029 23545 46063 23579
rect 11805 23477 11839 23511
rect 21833 23477 21867 23511
rect 29837 23477 29871 23511
rect 30757 23477 30791 23511
rect 33609 23477 33643 23511
rect 41613 23477 41647 23511
rect 46857 23477 46891 23511
rect 47041 23477 47075 23511
rect 47685 23477 47719 23511
rect 17141 23273 17175 23307
rect 23213 23273 23247 23307
rect 27169 23273 27203 23307
rect 32781 23273 32815 23307
rect 34713 23273 34747 23307
rect 43177 23273 43211 23307
rect 15669 23205 15703 23239
rect 24961 23205 24995 23239
rect 30297 23205 30331 23239
rect 11529 23137 11563 23171
rect 13553 23137 13587 23171
rect 19349 23137 19383 23171
rect 20269 23137 20303 23171
rect 21465 23137 21499 23171
rect 26341 23137 26375 23171
rect 28457 23137 28491 23171
rect 28917 23137 28951 23171
rect 31033 23137 31067 23171
rect 31309 23137 31343 23171
rect 33977 23137 34011 23171
rect 40509 23137 40543 23171
rect 46305 23137 46339 23171
rect 46489 23137 46523 23171
rect 48145 23137 48179 23171
rect 15485 23069 15519 23103
rect 17325 23069 17359 23103
rect 19533 23069 19567 23103
rect 19809 23069 19843 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 20729 23069 20763 23103
rect 24869 23069 24903 23103
rect 25053 23069 25087 23103
rect 25697 23069 25731 23103
rect 26525 23069 26559 23103
rect 26709 23069 26743 23103
rect 27353 23069 27387 23103
rect 28549 23069 28583 23103
rect 30113 23069 30147 23103
rect 33885 23069 33919 23103
rect 34069 23069 34103 23103
rect 34713 23069 34747 23103
rect 40049 23069 40083 23103
rect 42901 23069 42935 23103
rect 42993 23069 43027 23103
rect 43637 23069 43671 23103
rect 43821 23069 43855 23103
rect 45845 23069 45879 23103
rect 11805 23001 11839 23035
rect 21741 23001 21775 23035
rect 25513 23001 25547 23035
rect 25881 23001 25915 23035
rect 40693 23001 40727 23035
rect 42349 23001 42383 23035
rect 19717 22933 19751 22967
rect 39865 22933 39899 22967
rect 43729 22933 43763 22967
rect 45661 22933 45695 22967
rect 13093 22729 13127 22763
rect 22845 22729 22879 22763
rect 30481 22729 30515 22763
rect 32229 22729 32263 22763
rect 40693 22729 40727 22763
rect 29009 22661 29043 22695
rect 42533 22661 42567 22695
rect 42717 22661 42751 22695
rect 43361 22661 43395 22695
rect 45385 22661 45419 22695
rect 11713 22593 11747 22627
rect 13001 22593 13035 22627
rect 15117 22593 15151 22627
rect 22753 22593 22787 22627
rect 25605 22593 25639 22627
rect 27905 22593 27939 22627
rect 31125 22593 31159 22627
rect 32137 22593 32171 22627
rect 40233 22593 40267 22627
rect 42809 22593 42843 22627
rect 43269 22593 43303 22627
rect 43453 22593 43487 22627
rect 44741 22593 44775 22627
rect 45201 22593 45235 22627
rect 47593 22593 47627 22627
rect 11805 22525 11839 22559
rect 12081 22525 12115 22559
rect 28733 22525 28767 22559
rect 45753 22525 45787 22559
rect 47869 22525 47903 22559
rect 42533 22457 42567 22491
rect 48145 22457 48179 22491
rect 15209 22389 15243 22423
rect 25421 22389 25455 22423
rect 28089 22389 28123 22423
rect 31309 22389 31343 22423
rect 40325 22389 40359 22423
rect 44557 22389 44591 22423
rect 47685 22389 47719 22423
rect 26157 22185 26191 22219
rect 29561 22185 29595 22219
rect 35081 22185 35115 22219
rect 35541 22185 35575 22219
rect 13185 22117 13219 22151
rect 25973 22117 26007 22151
rect 26709 22117 26743 22151
rect 30849 22117 30883 22151
rect 14841 22049 14875 22083
rect 15025 22049 15059 22083
rect 15301 22049 15335 22083
rect 24409 22049 24443 22083
rect 30573 22049 30607 22083
rect 31309 22049 31343 22083
rect 31585 22049 31619 22083
rect 45201 22049 45235 22083
rect 45385 22049 45419 22083
rect 45753 22049 45787 22083
rect 47501 22049 47535 22083
rect 11805 21981 11839 22015
rect 12357 21981 12391 22015
rect 12541 21981 12575 22015
rect 13001 21981 13035 22015
rect 17141 21981 17175 22015
rect 18521 21981 18555 22015
rect 19257 21981 19291 22015
rect 20361 21981 20395 22015
rect 22477 21981 22511 22015
rect 24685 21981 24719 22015
rect 26617 21981 26651 22015
rect 28365 21981 28399 22015
rect 29745 21981 29779 22015
rect 30481 21981 30515 22015
rect 34805 21981 34839 22015
rect 40325 21981 40359 22015
rect 40417 21981 40451 22015
rect 43361 21981 43395 22015
rect 43545 21981 43579 22015
rect 44189 21981 44223 22015
rect 44373 21981 44407 22015
rect 47685 21981 47719 22015
rect 20913 21913 20947 21947
rect 22845 21913 22879 21947
rect 25697 21913 25731 21947
rect 28641 21913 28675 21947
rect 40601 21913 40635 21947
rect 48053 21913 48087 21947
rect 11805 21845 11839 21879
rect 12449 21845 12483 21879
rect 17233 21845 17267 21879
rect 18613 21845 18647 21879
rect 19349 21845 19383 21879
rect 33057 21845 33091 21879
rect 35265 21845 35299 21879
rect 43453 21845 43487 21879
rect 44373 21845 44407 21879
rect 47777 21845 47811 21879
rect 47869 21845 47903 21879
rect 22385 21641 22419 21675
rect 25053 21641 25087 21675
rect 25697 21641 25731 21675
rect 27537 21641 27571 21675
rect 32229 21641 32263 21675
rect 10885 21573 10919 21607
rect 11713 21573 11747 21607
rect 16865 21573 16899 21607
rect 19625 21573 19659 21607
rect 21281 21573 21315 21607
rect 35265 21573 35299 21607
rect 42809 21573 42843 21607
rect 45201 21573 45235 21607
rect 47593 21573 47627 21607
rect 47777 21573 47811 21607
rect 10793 21505 10827 21539
rect 16681 21505 16715 21539
rect 22293 21505 22327 21539
rect 23213 21505 23247 21539
rect 23397 21505 23431 21539
rect 24869 21505 24903 21539
rect 24961 21505 24995 21539
rect 25237 21505 25271 21539
rect 25881 21505 25915 21539
rect 26157 21505 26191 21539
rect 27353 21505 27387 21539
rect 28273 21505 28307 21539
rect 30665 21505 30699 21539
rect 32137 21505 32171 21539
rect 34621 21505 34655 21539
rect 42993 21505 43027 21539
rect 43913 21505 43947 21539
rect 46213 21505 46247 21539
rect 11529 21437 11563 21471
rect 11989 21437 12023 21471
rect 14289 21437 14323 21471
rect 14473 21437 14507 21471
rect 14749 21437 14783 21471
rect 17141 21437 17175 21471
rect 19441 21437 19475 21471
rect 25973 21437 26007 21471
rect 26065 21437 26099 21471
rect 28457 21437 28491 21471
rect 29009 21437 29043 21471
rect 31493 21437 31527 21471
rect 35173 21437 35207 21471
rect 36185 21437 36219 21471
rect 44649 21437 44683 21471
rect 46489 21437 46523 21471
rect 24685 21369 24719 21403
rect 34437 21369 34471 21403
rect 47961 21369 47995 21403
rect 43177 21301 43211 21335
rect 43729 21301 43763 21335
rect 14105 21097 14139 21131
rect 15669 21097 15703 21131
rect 27169 21097 27203 21131
rect 28641 21097 28675 21131
rect 45385 21097 45419 21131
rect 23765 21029 23799 21063
rect 24961 21029 24995 21063
rect 24409 20961 24443 20995
rect 25697 20961 25731 20995
rect 30021 20961 30055 20995
rect 36553 20961 36587 20995
rect 48145 20961 48179 20995
rect 11529 20893 11563 20927
rect 14381 20893 14415 20927
rect 14841 20893 14875 20927
rect 15577 20893 15611 20927
rect 16589 20893 16623 20927
rect 17325 20893 17359 20927
rect 18061 20893 18095 20927
rect 19257 20893 19291 20927
rect 21097 20893 21131 20927
rect 21649 20893 21683 20927
rect 21741 20893 21775 20927
rect 24685 20893 24719 20927
rect 25421 20893 25455 20927
rect 27997 20893 28031 20927
rect 28549 20893 28583 20927
rect 29561 20893 29595 20927
rect 42349 20893 42383 20927
rect 42533 20893 42567 20927
rect 43085 20893 43119 20927
rect 43453 20893 43487 20927
rect 45201 20893 45235 20927
rect 46305 20893 46339 20927
rect 11805 20825 11839 20859
rect 14105 20825 14139 20859
rect 19441 20825 19475 20859
rect 23213 20825 23247 20859
rect 23581 20825 23615 20859
rect 24593 20825 24627 20859
rect 29745 20825 29779 20859
rect 35541 20825 35575 20859
rect 35633 20825 35667 20859
rect 45017 20825 45051 20859
rect 46489 20825 46523 20859
rect 13277 20757 13311 20791
rect 14289 20757 14323 20791
rect 15025 20757 15059 20791
rect 16773 20757 16807 20791
rect 17509 20757 17543 20791
rect 18153 20757 18187 20791
rect 21925 20757 21959 20791
rect 23397 20757 23431 20791
rect 23489 20757 23523 20791
rect 24777 20757 24811 20791
rect 27997 20757 28031 20791
rect 42533 20757 42567 20791
rect 44097 20757 44131 20791
rect 24317 20553 24351 20587
rect 25513 20553 25547 20587
rect 27169 20553 27203 20587
rect 29193 20553 29227 20587
rect 42625 20553 42659 20587
rect 43361 20553 43395 20587
rect 43453 20553 43487 20587
rect 48053 20553 48087 20587
rect 14933 20485 14967 20519
rect 15133 20485 15167 20519
rect 18981 20485 19015 20519
rect 19197 20485 19231 20519
rect 19993 20485 20027 20519
rect 20193 20485 20227 20519
rect 23949 20485 23983 20519
rect 24165 20485 24199 20519
rect 45385 20485 45419 20519
rect 47961 20485 47995 20519
rect 11989 20417 12023 20451
rect 16773 20417 16807 20451
rect 17601 20417 17635 20451
rect 17877 20417 17911 20451
rect 18061 20417 18095 20451
rect 21833 20417 21867 20451
rect 25513 20417 25547 20451
rect 26065 20417 26099 20451
rect 26985 20417 27019 20451
rect 29101 20417 29135 20451
rect 30481 20417 30515 20451
rect 33425 20417 33459 20451
rect 42441 20417 42475 20451
rect 42625 20417 42659 20451
rect 43085 20417 43119 20451
rect 43269 20417 43303 20451
rect 43637 20417 43671 20451
rect 44373 20417 44407 20451
rect 44557 20417 44591 20451
rect 12173 20349 12207 20383
rect 12633 20349 12667 20383
rect 12909 20349 12943 20383
rect 14381 20349 14415 20383
rect 44097 20349 44131 20383
rect 45201 20349 45235 20383
rect 45753 20349 45787 20383
rect 15301 20281 15335 20315
rect 19349 20281 19383 20315
rect 15117 20213 15151 20247
rect 16865 20213 16899 20247
rect 17417 20213 17451 20247
rect 19165 20213 19199 20247
rect 20177 20213 20211 20247
rect 20361 20213 20395 20247
rect 22017 20213 22051 20247
rect 24133 20213 24167 20247
rect 26157 20213 26191 20247
rect 30573 20213 30607 20247
rect 33241 20213 33275 20247
rect 44373 20213 44407 20247
rect 12909 20009 12943 20043
rect 14105 20009 14139 20043
rect 14657 20009 14691 20043
rect 16313 20009 16347 20043
rect 19809 20009 19843 20043
rect 43085 20009 43119 20043
rect 45845 20009 45879 20043
rect 15485 19941 15519 19975
rect 16497 19941 16531 19975
rect 20821 19941 20855 19975
rect 23581 19941 23615 19975
rect 43913 19941 43947 19975
rect 16957 19873 16991 19907
rect 17233 19873 17267 19907
rect 24961 19873 24995 19907
rect 25421 19873 25455 19907
rect 30481 19873 30515 19907
rect 30665 19873 30699 19907
rect 33149 19873 33183 19907
rect 45201 19873 45235 19907
rect 46305 19873 46339 19907
rect 2053 19805 2087 19839
rect 12817 19805 12851 19839
rect 14286 19805 14320 19839
rect 14749 19805 14783 19839
rect 15209 19805 15243 19839
rect 19441 19805 19475 19839
rect 20269 19805 20303 19839
rect 20637 19805 20671 19839
rect 21741 19805 21775 19839
rect 23857 19805 23891 19839
rect 25053 19805 25087 19839
rect 25973 19805 26007 19839
rect 29745 19805 29779 19839
rect 43085 19805 43119 19839
rect 43269 19805 43303 19839
rect 43821 19805 43855 19839
rect 44005 19805 44039 19839
rect 16129 19737 16163 19771
rect 16329 19737 16363 19771
rect 19257 19737 19291 19771
rect 19533 19737 19567 19771
rect 20453 19737 20487 19771
rect 23581 19737 23615 19771
rect 23765 19737 23799 19771
rect 32321 19737 32355 19771
rect 33241 19737 33275 19771
rect 34161 19737 34195 19771
rect 46489 19737 46523 19771
rect 48145 19737 48179 19771
rect 14289 19669 14323 19703
rect 15669 19669 15703 19703
rect 18705 19669 18739 19703
rect 19625 19669 19659 19703
rect 20545 19669 20579 19703
rect 21833 19669 21867 19703
rect 26065 19669 26099 19703
rect 29561 19669 29595 19703
rect 13737 19465 13771 19499
rect 15485 19465 15519 19499
rect 19625 19465 19659 19499
rect 26065 19465 26099 19499
rect 28089 19465 28123 19499
rect 29653 19465 29687 19499
rect 45477 19465 45511 19499
rect 47685 19465 47719 19499
rect 17417 19397 17451 19431
rect 28641 19397 28675 19431
rect 29101 19397 29135 19431
rect 32321 19397 32355 19431
rect 46305 19397 46339 19431
rect 46489 19397 46523 19431
rect 1777 19329 1811 19363
rect 12817 19329 12851 19363
rect 13645 19329 13679 19363
rect 15301 19329 15335 19363
rect 15577 19329 15611 19363
rect 17233 19329 17267 19363
rect 19073 19329 19107 19363
rect 19533 19329 19567 19363
rect 20729 19329 20763 19363
rect 23857 19329 23891 19363
rect 26985 19329 27019 19363
rect 28457 19329 28491 19363
rect 29469 19329 29503 19363
rect 43085 19329 43119 19363
rect 45661 19329 45695 19363
rect 46397 19329 46431 19363
rect 47593 19329 47627 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 12909 19261 12943 19295
rect 15117 19261 15151 19295
rect 20821 19261 20855 19295
rect 21833 19261 21867 19295
rect 22109 19261 22143 19295
rect 24317 19261 24351 19295
rect 24593 19261 24627 19295
rect 28825 19261 28859 19295
rect 29285 19261 29319 19295
rect 32229 19261 32263 19295
rect 32505 19261 32539 19295
rect 46673 19261 46707 19295
rect 21097 19193 21131 19227
rect 33609 19193 33643 19227
rect 46121 19193 46155 19227
rect 13185 19125 13219 19159
rect 27077 19125 27111 19159
rect 43177 19125 43211 19159
rect 2237 18921 2271 18955
rect 16957 18921 16991 18955
rect 21465 18921 21499 18955
rect 23489 18921 23523 18955
rect 24869 18921 24903 18955
rect 27169 18921 27203 18955
rect 33149 18921 33183 18955
rect 33425 18921 33459 18955
rect 48053 18921 48087 18955
rect 11713 18785 11747 18819
rect 12449 18785 12483 18819
rect 23029 18785 23063 18819
rect 25697 18785 25731 18819
rect 29653 18785 29687 18819
rect 30113 18785 30147 18819
rect 42809 18785 42843 18819
rect 45845 18785 45879 18819
rect 2145 18717 2179 18751
rect 14749 18717 14783 18751
rect 15209 18717 15243 18751
rect 21465 18717 21499 18751
rect 22937 18717 22971 18751
rect 23489 18717 23523 18751
rect 23673 18717 23707 18751
rect 24777 18717 24811 18751
rect 25421 18717 25455 18751
rect 28457 18717 28491 18751
rect 28641 18717 28675 18751
rect 29745 18717 29779 18751
rect 30665 18717 30699 18751
rect 32965 18717 32999 18751
rect 42625 18717 42659 18751
rect 45201 18717 45235 18751
rect 45385 18717 45419 18751
rect 46213 18717 46247 18751
rect 46489 18717 46523 18751
rect 46857 18717 46891 18751
rect 47317 18717 47351 18751
rect 47961 18717 47995 18751
rect 11897 18649 11931 18683
rect 15485 18649 15519 18683
rect 28549 18649 28583 18683
rect 30849 18649 30883 18683
rect 32505 18649 32539 18683
rect 44465 18649 44499 18683
rect 46121 18649 46155 18683
rect 14565 18581 14599 18615
rect 45293 18581 45327 18615
rect 47409 18581 47443 18615
rect 47961 18377 47995 18411
rect 11897 18309 11931 18343
rect 13645 18309 13679 18343
rect 15945 18309 15979 18343
rect 16773 18309 16807 18343
rect 22845 18309 22879 18343
rect 23581 18309 23615 18343
rect 28089 18309 28123 18343
rect 45385 18309 45419 18343
rect 47777 18309 47811 18343
rect 1869 18241 1903 18275
rect 11805 18241 11839 18275
rect 15669 18241 15703 18275
rect 16681 18241 16715 18275
rect 22753 18241 22787 18275
rect 27629 18241 27663 18275
rect 27905 18241 27939 18275
rect 28733 18241 28767 18275
rect 32137 18241 32171 18275
rect 33241 18241 33275 18275
rect 41245 18241 41279 18275
rect 41429 18241 41463 18275
rect 41705 18241 41739 18275
rect 43729 18241 43763 18275
rect 47593 18241 47627 18275
rect 13369 18173 13403 18207
rect 17693 18173 17727 18207
rect 17969 18173 18003 18207
rect 23397 18173 23431 18207
rect 25237 18173 25271 18207
rect 27997 18173 28031 18207
rect 28549 18173 28583 18207
rect 29745 18173 29779 18207
rect 29929 18173 29963 18207
rect 31125 18173 31159 18207
rect 32597 18173 32631 18207
rect 44649 18173 44683 18207
rect 45201 18173 45235 18207
rect 45661 18173 45695 18207
rect 19441 18105 19475 18139
rect 41613 18105 41647 18139
rect 1961 18037 1995 18071
rect 15117 18037 15151 18071
rect 27721 18037 27755 18071
rect 28917 18037 28951 18071
rect 32229 18037 32263 18071
rect 33057 18037 33091 18071
rect 14381 17833 14415 17867
rect 17509 17833 17543 17867
rect 18613 17833 18647 17867
rect 19809 17833 19843 17867
rect 23305 17833 23339 17867
rect 30205 17833 30239 17867
rect 45661 17833 45695 17867
rect 11713 17697 11747 17731
rect 12449 17697 12483 17731
rect 19349 17697 19383 17731
rect 41429 17697 41463 17731
rect 41613 17697 41647 17731
rect 41889 17697 41923 17731
rect 45017 17697 45051 17731
rect 46305 17697 46339 17731
rect 14289 17629 14323 17663
rect 17325 17629 17359 17663
rect 18521 17629 18555 17663
rect 19441 17629 19475 17663
rect 20545 17629 20579 17663
rect 27077 17629 27111 17663
rect 27905 17629 27939 17663
rect 30113 17629 30147 17663
rect 31033 17629 31067 17663
rect 44097 17629 44131 17663
rect 45385 17629 45419 17663
rect 45477 17629 45511 17663
rect 11897 17561 11931 17595
rect 23121 17561 23155 17595
rect 23337 17561 23371 17595
rect 27261 17561 27295 17595
rect 28089 17561 28123 17595
rect 28457 17561 28491 17595
rect 31217 17561 31251 17595
rect 32873 17561 32907 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 20637 17493 20671 17527
rect 23489 17493 23523 17527
rect 27445 17493 27479 17527
rect 28181 17493 28215 17527
rect 28273 17493 28307 17527
rect 44189 17493 44223 17527
rect 11897 17289 11931 17323
rect 27261 17289 27295 17323
rect 46857 17289 46891 17323
rect 47685 17289 47719 17323
rect 14013 17221 14047 17255
rect 20361 17221 20395 17255
rect 20577 17221 20611 17255
rect 44281 17221 44315 17255
rect 11805 17153 11839 17187
rect 13921 17153 13955 17187
rect 15853 17153 15887 17187
rect 17509 17153 17543 17187
rect 24225 17153 24259 17187
rect 25237 17153 25271 17187
rect 25973 17153 26007 17187
rect 27077 17153 27111 17187
rect 27261 17153 27295 17187
rect 27997 17153 28031 17187
rect 28089 17153 28123 17187
rect 28273 17153 28307 17187
rect 28825 17153 28859 17187
rect 29193 17153 29227 17187
rect 46765 17153 46799 17187
rect 46949 17153 46983 17187
rect 47593 17153 47627 17187
rect 17601 17085 17635 17119
rect 18153 17085 18187 17119
rect 18429 17085 18463 17119
rect 21833 17085 21867 17119
rect 22109 17085 22143 17119
rect 44097 17085 44131 17119
rect 44557 17085 44591 17119
rect 19901 17017 19935 17051
rect 20729 17017 20763 17051
rect 2053 16949 2087 16983
rect 15945 16949 15979 16983
rect 20545 16949 20579 16983
rect 23581 16949 23615 16983
rect 24225 16949 24259 16983
rect 25237 16949 25271 16983
rect 26065 16949 26099 16983
rect 30665 16949 30699 16983
rect 18521 16745 18555 16779
rect 22937 16745 22971 16779
rect 19533 16677 19567 16711
rect 28549 16677 28583 16711
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 15669 16609 15703 16643
rect 15853 16609 15887 16643
rect 24409 16609 24443 16643
rect 24685 16609 24719 16643
rect 26157 16609 26191 16643
rect 42625 16609 42659 16643
rect 46305 16609 46339 16643
rect 18521 16541 18555 16575
rect 18705 16541 18739 16575
rect 19717 16541 19751 16575
rect 19809 16541 19843 16575
rect 20637 16541 20671 16575
rect 23121 16541 23155 16575
rect 23397 16541 23431 16575
rect 23581 16541 23615 16575
rect 26617 16541 26651 16575
rect 27813 16541 27847 16575
rect 27997 16541 28031 16575
rect 28457 16541 28491 16575
rect 31217 16541 31251 16575
rect 45017 16541 45051 16575
rect 1593 16473 1627 16507
rect 17509 16473 17543 16507
rect 19533 16473 19567 16507
rect 20821 16473 20855 16507
rect 22477 16473 22511 16507
rect 42809 16473 42843 16507
rect 44465 16473 44499 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 26709 16405 26743 16439
rect 27997 16405 28031 16439
rect 31309 16405 31343 16439
rect 45109 16405 45143 16439
rect 2145 16201 2179 16235
rect 19349 16201 19383 16235
rect 22017 16201 22051 16235
rect 25605 16201 25639 16235
rect 27169 16201 27203 16235
rect 28549 16201 28583 16235
rect 42901 16201 42935 16235
rect 16037 16133 16071 16167
rect 16865 16133 16899 16167
rect 44097 16133 44131 16167
rect 2053 16065 2087 16099
rect 15945 16065 15979 16099
rect 19257 16065 19291 16099
rect 22017 16065 22051 16099
rect 25237 16065 25271 16099
rect 27077 16065 27111 16099
rect 27261 16065 27295 16099
rect 28365 16065 28399 16099
rect 28549 16065 28583 16099
rect 42809 16065 42843 16099
rect 47777 16065 47811 16099
rect 16681 15997 16715 16031
rect 17141 15997 17175 16031
rect 22753 15997 22787 16031
rect 22937 15997 22971 16031
rect 24317 15997 24351 16031
rect 25145 15997 25179 16031
rect 43913 15997 43947 16031
rect 45109 15997 45143 16031
rect 21833 15657 21867 15691
rect 23213 15657 23247 15691
rect 23397 15657 23431 15691
rect 24501 15657 24535 15691
rect 47685 15657 47719 15691
rect 25329 15521 25363 15555
rect 27077 15521 27111 15555
rect 30389 15521 30423 15555
rect 30573 15521 30607 15555
rect 2053 15453 2087 15487
rect 21741 15453 21775 15487
rect 24409 15453 24443 15487
rect 24593 15453 24627 15487
rect 23029 15385 23063 15419
rect 25605 15385 25639 15419
rect 32229 15385 32263 15419
rect 23239 15317 23273 15351
rect 23397 15113 23431 15147
rect 1777 14977 1811 15011
rect 23305 14977 23339 15011
rect 24409 14977 24443 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 24317 14909 24351 14943
rect 24777 14909 24811 14943
rect 2329 14569 2363 14603
rect 2237 14365 2271 14399
rect 22017 13345 22051 13379
rect 23673 13345 23707 13379
rect 47685 13277 47719 13311
rect 22201 13209 22235 13243
rect 22477 12937 22511 12971
rect 1409 12801 1443 12835
rect 22385 12801 22419 12835
rect 1593 12597 1627 12631
rect 47777 12597 47811 12631
rect 46305 12257 46339 12291
rect 48145 12257 48179 12291
rect 46489 12121 46523 12155
rect 47685 11849 47719 11883
rect 46673 11713 46707 11747
rect 47593 11713 47627 11747
rect 46765 11509 46799 11543
rect 46305 11169 46339 11203
rect 46489 11169 46523 11203
rect 48145 11033 48179 11067
rect 47593 10625 47627 10659
rect 47041 10421 47075 10455
rect 47685 10421 47719 10455
rect 46305 10081 46339 10115
rect 46489 10081 46523 10115
rect 48145 10081 48179 10115
rect 47869 9537 47903 9571
rect 48053 9401 48087 9435
rect 47777 8857 47811 8891
rect 47869 8789 47903 8823
rect 48145 8449 48179 8483
rect 47961 8245 47995 8279
rect 45569 7905 45603 7939
rect 46581 7905 46615 7939
rect 47133 7905 47167 7939
rect 47409 7905 47443 7939
rect 45661 7769 45695 7803
rect 47225 7769 47259 7803
rect 47593 7497 47627 7531
rect 46305 7361 46339 7395
rect 47777 7361 47811 7395
rect 46765 7293 46799 7327
rect 45937 7225 45971 7259
rect 46397 7157 46431 7191
rect 41797 6817 41831 6851
rect 47317 6817 47351 6851
rect 47593 6817 47627 6851
rect 40325 6681 40359 6715
rect 40785 6681 40819 6715
rect 40877 6681 40911 6715
rect 40693 6409 40727 6443
rect 48053 6409 48087 6443
rect 40877 6273 40911 6307
rect 47961 6273 47995 6307
rect 41889 5729 41923 5763
rect 42717 5729 42751 5763
rect 41981 5593 42015 5627
rect 40693 5321 40727 5355
rect 21833 5185 21867 5219
rect 22477 5185 22511 5219
rect 40233 5185 40267 5219
rect 47777 5185 47811 5219
rect 21925 5049 21959 5083
rect 47961 5049 47995 5083
rect 22569 4981 22603 5015
rect 40325 4981 40359 5015
rect 22109 4641 22143 4675
rect 22753 4641 22787 4675
rect 37933 4641 37967 4675
rect 47593 4641 47627 4675
rect 7389 4573 7423 4607
rect 20729 4573 20763 4607
rect 21373 4573 21407 4607
rect 22017 4573 22051 4607
rect 22661 4573 22695 4607
rect 23489 4573 23523 4607
rect 39957 4573 39991 4607
rect 40601 4573 40635 4607
rect 46673 4573 46707 4607
rect 47317 4573 47351 4607
rect 36553 4505 36587 4539
rect 36921 4505 36955 4539
rect 37013 4505 37047 4539
rect 7481 4437 7515 4471
rect 20821 4437 20855 4471
rect 21465 4437 21499 4471
rect 23305 4437 23339 4471
rect 40049 4437 40083 4471
rect 40693 4437 40727 4471
rect 46765 4437 46799 4471
rect 21925 4233 21959 4267
rect 23213 4233 23247 4267
rect 36553 4233 36587 4267
rect 25513 4165 25547 4199
rect 37657 4165 37691 4199
rect 38577 4165 38611 4199
rect 46581 4165 46615 4199
rect 47777 4165 47811 4199
rect 2053 4097 2087 4131
rect 12081 4097 12115 4131
rect 13737 4097 13771 4131
rect 16681 4097 16715 4131
rect 17693 4097 17727 4131
rect 18337 4097 18371 4131
rect 19441 4097 19475 4131
rect 20085 4097 20119 4131
rect 20729 4097 20763 4131
rect 21833 4097 21867 4131
rect 22477 4097 22511 4131
rect 23121 4097 23155 4131
rect 23765 4097 23799 4131
rect 23857 4097 23891 4131
rect 24593 4097 24627 4131
rect 36737 4097 36771 4131
rect 39405 4097 39439 4131
rect 42993 4097 43027 4131
rect 6929 4029 6963 4063
rect 7389 4029 7423 4063
rect 7573 4029 7607 4063
rect 8401 4029 8435 4063
rect 19533 4029 19567 4063
rect 22569 4029 22603 4063
rect 25421 4029 25455 4063
rect 26433 4029 26467 4063
rect 37565 4029 37599 4063
rect 40049 4029 40083 4063
rect 40233 4029 40267 4063
rect 40509 4029 40543 4063
rect 48053 4029 48087 4063
rect 17785 3961 17819 3995
rect 46765 3961 46799 3995
rect 2145 3893 2179 3927
rect 2881 3893 2915 3927
rect 9873 3893 9907 3927
rect 12173 3893 12207 3927
rect 13829 3893 13863 3927
rect 16773 3893 16807 3927
rect 18429 3893 18463 3927
rect 20177 3893 20211 3927
rect 20821 3893 20855 3927
rect 24685 3893 24719 3927
rect 39497 3893 39531 3927
rect 43085 3893 43119 3927
rect 43821 3893 43855 3927
rect 46029 3893 46063 3927
rect 8309 3689 8343 3723
rect 17233 3689 17267 3723
rect 24961 3689 24995 3723
rect 38577 3689 38611 3723
rect 23029 3621 23063 3655
rect 39129 3621 39163 3655
rect 40509 3621 40543 3655
rect 3985 3553 4019 3587
rect 9229 3553 9263 3587
rect 9689 3553 9723 3587
rect 14933 3553 14967 3587
rect 15393 3553 15427 3587
rect 21925 3553 21959 3587
rect 40969 3553 41003 3587
rect 42625 3553 42659 3587
rect 42809 3553 42843 3587
rect 43177 3553 43211 3587
rect 46305 3553 46339 3587
rect 2697 3485 2731 3519
rect 6469 3485 6503 3519
rect 7113 3485 7147 3519
rect 7573 3485 7607 3519
rect 8217 3485 8251 3519
rect 11713 3485 11747 3519
rect 14289 3485 14323 3519
rect 15025 3485 15059 3519
rect 15853 3485 15887 3519
rect 15945 3485 15979 3519
rect 16497 3485 16531 3519
rect 17141 3485 17175 3519
rect 17785 3485 17819 3519
rect 18521 3485 18555 3519
rect 19257 3485 19291 3519
rect 20085 3485 20119 3519
rect 20545 3485 20579 3519
rect 21189 3485 21223 3519
rect 21281 3485 21315 3519
rect 21833 3485 21867 3519
rect 23857 3485 23891 3519
rect 27261 3485 27295 3519
rect 31493 3485 31527 3519
rect 32413 3485 32447 3519
rect 38485 3485 38519 3519
rect 39313 3485 39347 3519
rect 39865 3485 39899 3519
rect 40049 3485 40083 3519
rect 41153 3485 41187 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 1869 3417 1903 3451
rect 2237 3417 2271 3451
rect 9413 3417 9447 3451
rect 24869 3417 24903 3451
rect 25605 3417 25639 3451
rect 25697 3417 25731 3451
rect 26617 3417 26651 3451
rect 45753 3417 45787 3451
rect 46489 3417 46523 3451
rect 48145 3417 48179 3451
rect 2789 3349 2823 3383
rect 7665 3349 7699 3383
rect 16589 3349 16623 3383
rect 17877 3349 17911 3383
rect 18613 3349 18647 3383
rect 19349 3349 19383 3383
rect 20637 3349 20671 3383
rect 27077 3349 27111 3383
rect 31585 3349 31619 3383
rect 41613 3349 41647 3383
rect 16773 3145 16807 3179
rect 17969 3145 18003 3179
rect 18613 3145 18647 3179
rect 26157 3145 26191 3179
rect 27537 3145 27571 3179
rect 36737 3145 36771 3179
rect 39957 3145 39991 3179
rect 40969 3145 41003 3179
rect 47869 3145 47903 3179
rect 2053 3077 2087 3111
rect 7481 3077 7515 3111
rect 10149 3077 10183 3111
rect 11713 3077 11747 3111
rect 14013 3077 14047 3111
rect 19625 3077 19659 3111
rect 32413 3077 32447 3111
rect 39589 3077 39623 3111
rect 45385 3077 45419 3111
rect 1869 3009 1903 3043
rect 7297 3009 7331 3043
rect 10057 3009 10091 3043
rect 11529 3009 11563 3043
rect 13829 3009 13863 3043
rect 16681 3009 16715 3043
rect 17877 3009 17911 3043
rect 18521 3009 18555 3043
rect 19441 3009 19475 3043
rect 22201 3009 22235 3043
rect 22845 3009 22879 3043
rect 25697 3009 25731 3043
rect 27445 3009 27479 3043
rect 32229 3009 32263 3043
rect 36277 3009 36311 3043
rect 39773 3009 39807 3043
rect 40417 3009 40451 3043
rect 41613 3033 41647 3067
rect 42441 3009 42475 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2329 2941 2363 2975
rect 7757 2941 7791 2975
rect 11989 2941 12023 2975
rect 14289 2941 14323 2975
rect 19901 2941 19935 2975
rect 23029 2941 23063 2975
rect 23581 2941 23615 2975
rect 33425 2941 33459 2975
rect 40693 2941 40727 2975
rect 42625 2941 42659 2975
rect 42901 2941 42935 2975
rect 47041 2941 47075 2975
rect 22385 2873 22419 2907
rect 41429 2873 41463 2907
rect 25789 2805 25823 2839
rect 36369 2805 36403 2839
rect 40509 2805 40543 2839
rect 5273 2601 5307 2635
rect 17877 2601 17911 2635
rect 18521 2601 18555 2635
rect 19349 2601 19383 2635
rect 19993 2601 20027 2635
rect 20913 2601 20947 2635
rect 28641 2601 28675 2635
rect 29745 2601 29779 2635
rect 35541 2601 35575 2635
rect 36369 2601 36403 2635
rect 39129 2601 39163 2635
rect 41705 2601 41739 2635
rect 17325 2533 17359 2567
rect 22017 2533 22051 2567
rect 45569 2533 45603 2567
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2881 2465 2915 2499
rect 6561 2465 6595 2499
rect 6745 2465 6779 2499
rect 7021 2465 7055 2499
rect 24501 2465 24535 2499
rect 24685 2465 24719 2499
rect 25145 2465 25179 2499
rect 27261 2465 27295 2499
rect 40509 2465 40543 2499
rect 46489 2465 46523 2499
rect 47869 2465 47903 2499
rect 3801 2397 3835 2431
rect 5457 2397 5491 2431
rect 15301 2397 15335 2431
rect 15577 2397 15611 2431
rect 17785 2397 17819 2431
rect 18429 2397 18463 2431
rect 19257 2397 19291 2431
rect 19901 2397 19935 2431
rect 22385 2397 22419 2431
rect 22845 2397 22879 2431
rect 26985 2397 27019 2431
rect 28457 2397 28491 2431
rect 29929 2397 29963 2431
rect 35725 2397 35759 2431
rect 38117 2397 38151 2431
rect 39313 2397 39347 2431
rect 41889 2397 41923 2431
rect 43637 2397 43671 2431
rect 43913 2397 43947 2431
rect 46213 2397 46247 2431
rect 47685 2397 47719 2431
rect 9413 2329 9447 2363
rect 17141 2329 17175 2363
rect 20821 2329 20855 2363
rect 36277 2329 36311 2363
rect 40325 2329 40359 2363
rect 41061 2329 41095 2363
rect 45385 2329 45419 2363
rect 3985 2261 4019 2295
rect 9689 2261 9723 2295
rect 38301 2261 38335 2295
rect 41153 2261 41187 2295
<< metal1 >>
rect 15930 47540 15936 47592
rect 15988 47580 15994 47592
rect 20070 47580 20076 47592
rect 15988 47552 20076 47580
rect 15988 47540 15994 47552
rect 20070 47540 20076 47552
rect 20128 47540 20134 47592
rect 20254 47540 20260 47592
rect 20312 47580 20318 47592
rect 28258 47580 28264 47592
rect 20312 47552 28264 47580
rect 20312 47540 20318 47552
rect 28258 47540 28264 47552
rect 28316 47540 28322 47592
rect 3050 47472 3056 47524
rect 3108 47512 3114 47524
rect 35434 47512 35440 47524
rect 3108 47484 35440 47512
rect 3108 47472 3114 47484
rect 35434 47472 35440 47484
rect 35492 47472 35498 47524
rect 2038 47404 2044 47456
rect 2096 47444 2102 47456
rect 40126 47444 40132 47456
rect 2096 47416 40132 47444
rect 2096 47404 2102 47416
rect 40126 47404 40132 47416
rect 40184 47404 40190 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 3050 47240 3056 47252
rect 3011 47212 3056 47240
rect 3050 47200 3056 47212
rect 3108 47200 3114 47252
rect 3326 47200 3332 47252
rect 3384 47240 3390 47252
rect 21818 47240 21824 47252
rect 3384 47212 21824 47240
rect 3384 47200 3390 47212
rect 21818 47200 21824 47212
rect 21876 47200 21882 47252
rect 28994 47200 29000 47252
rect 29052 47240 29058 47252
rect 29917 47243 29975 47249
rect 29917 47240 29929 47243
rect 29052 47212 29929 47240
rect 29052 47200 29058 47212
rect 29917 47209 29929 47212
rect 29963 47209 29975 47243
rect 29917 47203 29975 47209
rect 30190 47200 30196 47252
rect 30248 47240 30254 47252
rect 31021 47243 31079 47249
rect 31021 47240 31033 47243
rect 30248 47212 31033 47240
rect 30248 47200 30254 47212
rect 31021 47209 31033 47212
rect 31067 47209 31079 47243
rect 31021 47203 31079 47209
rect 41690 47200 41696 47252
rect 41748 47240 41754 47252
rect 46842 47240 46848 47252
rect 41748 47212 46848 47240
rect 41748 47200 41754 47212
rect 46842 47200 46848 47212
rect 46900 47200 46906 47252
rect 5077 47175 5135 47181
rect 5077 47141 5089 47175
rect 5123 47172 5135 47175
rect 20254 47172 20260 47184
rect 5123 47144 20260 47172
rect 5123 47141 5135 47144
rect 5077 47135 5135 47141
rect 20254 47132 20260 47144
rect 20312 47132 20318 47184
rect 20346 47132 20352 47184
rect 20404 47172 20410 47184
rect 22465 47175 22523 47181
rect 22465 47172 22477 47175
rect 20404 47144 22477 47172
rect 20404 47132 20410 47144
rect 22465 47141 22477 47144
rect 22511 47141 22523 47175
rect 44085 47175 44143 47181
rect 44085 47172 44097 47175
rect 22465 47135 22523 47141
rect 26206 47144 44097 47172
rect 2038 47104 2044 47116
rect 1999 47076 2044 47104
rect 2038 47064 2044 47076
rect 2096 47064 2102 47116
rect 11606 47064 11612 47116
rect 11664 47104 11670 47116
rect 11701 47107 11759 47113
rect 11701 47104 11713 47107
rect 11664 47076 11713 47104
rect 11664 47064 11670 47076
rect 11701 47073 11713 47076
rect 11747 47073 11759 47107
rect 11701 47067 11759 47073
rect 11977 47107 12035 47113
rect 11977 47073 11989 47107
rect 12023 47104 12035 47107
rect 12023 47076 13768 47104
rect 12023 47073 12035 47076
rect 11977 47067 12035 47073
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47036 1823 47039
rect 1946 47036 1952 47048
rect 1811 47008 1952 47036
rect 1811 47005 1823 47008
rect 1765 46999 1823 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4798 47036 4804 47048
rect 4759 47008 4804 47036
rect 3789 46999 3847 47005
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 5868 47008 6377 47036
rect 5868 46996 5874 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 7374 47036 7380 47048
rect 7335 47008 7380 47036
rect 6365 46999 6423 47005
rect 7374 46996 7380 47008
rect 7432 46996 7438 47048
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 9401 46999 9459 47005
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 12989 47039 13047 47045
rect 12989 47036 13001 47039
rect 12952 47008 13001 47036
rect 12952 46996 12958 47008
rect 12989 47005 13001 47008
rect 13035 47005 13047 47039
rect 13740 47036 13768 47076
rect 13814 47064 13820 47116
rect 13872 47104 13878 47116
rect 14093 47107 14151 47113
rect 14093 47104 14105 47107
rect 13872 47076 14105 47104
rect 13872 47064 13878 47076
rect 14093 47073 14105 47076
rect 14139 47073 14151 47107
rect 14093 47067 14151 47073
rect 14369 47107 14427 47113
rect 14369 47073 14381 47107
rect 14415 47104 14427 47107
rect 17402 47104 17408 47116
rect 14415 47076 17408 47104
rect 14415 47073 14427 47076
rect 14369 47067 14427 47073
rect 17402 47064 17408 47076
rect 17460 47064 17466 47116
rect 20070 47064 20076 47116
rect 20128 47104 20134 47116
rect 26206 47104 26234 47144
rect 44085 47141 44097 47144
rect 44131 47141 44143 47175
rect 44085 47135 44143 47141
rect 47854 47132 47860 47184
rect 47912 47172 47918 47184
rect 47949 47175 48007 47181
rect 47949 47172 47961 47175
rect 47912 47144 47961 47172
rect 47912 47132 47918 47144
rect 47949 47141 47961 47144
rect 47995 47141 48007 47175
rect 47949 47135 48007 47141
rect 44450 47104 44456 47116
rect 20128 47076 26234 47104
rect 43272 47076 44456 47104
rect 20128 47064 20134 47076
rect 14458 47036 14464 47048
rect 13740 47008 14464 47036
rect 12989 46999 13047 47005
rect 14458 46996 14464 47008
rect 14516 46996 14522 47048
rect 16574 46996 16580 47048
rect 16632 47036 16638 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16632 47008 16681 47036
rect 16632 46996 16638 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 16945 47039 17003 47045
rect 16945 47005 16957 47039
rect 16991 47036 17003 47039
rect 18598 47036 18604 47048
rect 16991 47008 18604 47036
rect 16991 47005 17003 47008
rect 16945 46999 17003 47005
rect 18598 46996 18604 47008
rect 18656 46996 18662 47048
rect 21082 47036 21088 47048
rect 21043 47008 21088 47036
rect 21082 46996 21088 47008
rect 21140 46996 21146 47048
rect 22002 47036 22008 47048
rect 21963 47008 22008 47036
rect 22002 46996 22008 47008
rect 22060 46996 22066 47048
rect 22649 47039 22707 47045
rect 22649 47005 22661 47039
rect 22695 47005 22707 47039
rect 22649 46999 22707 47005
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 2777 46931 2835 46937
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 2792 46900 2820 46931
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 6638 46968 6644 46980
rect 6599 46940 6644 46968
rect 6638 46928 6644 46940
rect 6696 46928 6702 46980
rect 7466 46928 7472 46980
rect 7524 46968 7530 46980
rect 7561 46971 7619 46977
rect 7561 46968 7573 46971
rect 7524 46940 7573 46968
rect 7524 46928 7530 46940
rect 7561 46937 7573 46940
rect 7607 46937 7619 46971
rect 7561 46931 7619 46937
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 19426 46968 19432 46980
rect 9585 46931 9643 46937
rect 13188 46940 19432 46968
rect 13188 46909 13216 46940
rect 19426 46928 19432 46940
rect 19484 46928 19490 46980
rect 19705 46971 19763 46977
rect 19705 46937 19717 46971
rect 19751 46937 19763 46971
rect 19705 46931 19763 46937
rect 2648 46872 2820 46900
rect 13173 46903 13231 46909
rect 2648 46860 2654 46872
rect 13173 46869 13185 46903
rect 13219 46869 13231 46903
rect 13173 46863 13231 46869
rect 16114 46860 16120 46912
rect 16172 46900 16178 46912
rect 16574 46900 16580 46912
rect 16172 46872 16580 46900
rect 16172 46860 16178 46872
rect 16574 46860 16580 46872
rect 16632 46860 16638 46912
rect 18690 46860 18696 46912
rect 18748 46900 18754 46912
rect 19720 46900 19748 46931
rect 19978 46928 19984 46980
rect 20036 46968 20042 46980
rect 20073 46971 20131 46977
rect 20073 46968 20085 46971
rect 20036 46940 20085 46968
rect 20036 46928 20042 46940
rect 20073 46937 20085 46940
rect 20119 46937 20131 46971
rect 22664 46968 22692 46999
rect 24578 46996 24584 47048
rect 24636 47036 24642 47048
rect 24765 47039 24823 47045
rect 24765 47036 24777 47039
rect 24636 47008 24777 47036
rect 24636 46996 24642 47008
rect 24765 47005 24777 47008
rect 24811 47005 24823 47039
rect 25498 47036 25504 47048
rect 25459 47008 25504 47036
rect 24765 46999 24823 47005
rect 25498 46996 25504 47008
rect 25556 46996 25562 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28537 47039 28595 47045
rect 28537 47036 28549 47039
rect 28408 47008 28549 47036
rect 28408 46996 28414 47008
rect 28537 47005 28549 47008
rect 28583 47005 28595 47039
rect 28537 46999 28595 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 30926 46996 30932 47048
rect 30984 47036 30990 47048
rect 31205 47039 31263 47045
rect 31205 47036 31217 47039
rect 30984 47008 31217 47036
rect 30984 46996 30990 47008
rect 31205 47005 31217 47008
rect 31251 47005 31263 47039
rect 31205 46999 31263 47005
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 42702 47036 42708 47048
rect 42663 47008 42708 47036
rect 38381 46999 38439 47005
rect 42702 46996 42708 47008
rect 42760 46996 42766 47048
rect 43272 47045 43300 47076
rect 44450 47064 44456 47076
rect 44508 47064 44514 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 43257 47039 43315 47045
rect 43257 47005 43269 47039
rect 43303 47005 43315 47039
rect 43257 46999 43315 47005
rect 43806 46996 43812 47048
rect 43864 47036 43870 47048
rect 43901 47039 43959 47045
rect 43901 47036 43913 47039
rect 43864 47008 43913 47036
rect 43864 46996 43870 47008
rect 43901 47005 43913 47008
rect 43947 47005 43959 47039
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 43901 46999 43959 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 20073 46931 20131 46937
rect 22020 46940 22692 46968
rect 18748 46872 19748 46900
rect 18748 46860 18754 46872
rect 20162 46860 20168 46912
rect 20220 46900 20226 46912
rect 22020 46900 22048 46940
rect 27798 46928 27804 46980
rect 27856 46968 27862 46980
rect 28721 46971 28779 46977
rect 28721 46968 28733 46971
rect 27856 46940 28733 46968
rect 27856 46928 27862 46940
rect 28721 46937 28733 46940
rect 28767 46937 28779 46971
rect 28721 46931 28779 46937
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 20220 46872 22048 46900
rect 20220 46860 20226 46872
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 40497 46931 40555 46937
rect 43346 46928 43352 46980
rect 43404 46968 43410 46980
rect 43441 46971 43499 46977
rect 43441 46968 43453 46971
rect 43404 46940 43453 46968
rect 43404 46928 43410 46940
rect 43441 46937 43453 46940
rect 43487 46937 43499 46971
rect 43441 46931 43499 46937
rect 45373 46971 45431 46977
rect 45373 46937 45385 46971
rect 45419 46968 45431 46971
rect 45462 46968 45468 46980
rect 45419 46940 45468 46968
rect 45419 46937 45431 46940
rect 45373 46931 45431 46937
rect 45462 46928 45468 46940
rect 45520 46928 45526 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 3878 46588 3884 46640
rect 3936 46628 3942 46640
rect 5813 46631 5871 46637
rect 5813 46628 5825 46631
rect 3936 46600 5825 46628
rect 3936 46588 3942 46600
rect 5813 46597 5825 46600
rect 5859 46597 5871 46631
rect 22002 46628 22008 46640
rect 5813 46591 5871 46597
rect 19444 46600 22008 46628
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 19444 46569 19472 46600
rect 22002 46588 22008 46600
rect 22060 46588 22066 46640
rect 19429 46563 19487 46569
rect 19429 46529 19441 46563
rect 19475 46529 19487 46563
rect 24578 46560 24584 46572
rect 24539 46532 24584 46560
rect 19429 46523 19487 46529
rect 24578 46520 24584 46532
rect 24636 46520 24642 46572
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 47946 46560 47952 46572
rect 47907 46532 47952 46560
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 3970 46492 3976 46504
rect 3931 46464 3976 46492
rect 3970 46452 3976 46464
rect 4028 46452 4034 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46492 4215 46495
rect 5074 46492 5080 46504
rect 4203 46464 5080 46492
rect 4203 46461 4215 46464
rect 4157 46455 4215 46461
rect 5074 46452 5080 46464
rect 5132 46452 5138 46504
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11517 46455 11575 46461
rect 11701 46495 11759 46501
rect 11701 46461 11713 46495
rect 11747 46492 11759 46495
rect 12066 46492 12072 46504
rect 11747 46464 12072 46492
rect 11747 46461 11759 46464
rect 11701 46455 11759 46461
rect 12066 46452 12072 46464
rect 12124 46452 12130 46504
rect 12161 46495 12219 46501
rect 12161 46461 12173 46495
rect 12207 46461 12219 46495
rect 12161 46455 12219 46461
rect 12176 46424 12204 46455
rect 13538 46452 13544 46504
rect 13596 46492 13602 46504
rect 13817 46495 13875 46501
rect 13817 46492 13829 46495
rect 13596 46464 13829 46492
rect 13596 46452 13602 46464
rect 13817 46461 13829 46464
rect 13863 46461 13875 46495
rect 13817 46455 13875 46461
rect 14001 46495 14059 46501
rect 14001 46461 14013 46495
rect 14047 46492 14059 46495
rect 14182 46492 14188 46504
rect 14047 46464 14188 46492
rect 14047 46461 14059 46464
rect 14001 46455 14059 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 19613 46495 19671 46501
rect 14332 46464 14377 46492
rect 14332 46452 14338 46464
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 20070 46492 20076 46504
rect 19659 46464 20076 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 20070 46452 20076 46464
rect 20128 46452 20134 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 31573 46495 31631 46501
rect 31573 46461 31585 46495
rect 31619 46492 31631 46495
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 31619 46464 32137 46492
rect 31619 46461 31631 46464
rect 31573 46455 31631 46461
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32306 46492 32312 46504
rect 32267 46464 32312 46492
rect 32125 46455 32183 46461
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46461 32643 46495
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 32585 46455 32643 46461
rect 10980 46396 12204 46424
rect 10980 46368 11008 46396
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 32600 46424 32628 46455
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 42889 46455 42947 46461
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45370 46492 45376 46504
rect 45331 46464 45376 46492
rect 45189 46455 45247 46461
rect 32272 46396 32628 46424
rect 32272 46384 32278 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 42576 46396 42932 46424
rect 45204 46424 45232 46455
rect 45370 46452 45376 46464
rect 45428 46452 45434 46504
rect 46750 46492 46756 46504
rect 46711 46464 46756 46492
rect 46750 46452 46756 46464
rect 46808 46452 46814 46504
rect 45646 46424 45652 46436
rect 45204 46396 45652 46424
rect 42576 46384 42582 46396
rect 45646 46384 45652 46396
rect 45704 46384 45710 46436
rect 1581 46359 1639 46365
rect 1581 46325 1593 46359
rect 1627 46356 1639 46359
rect 1670 46356 1676 46368
rect 1627 46328 1676 46356
rect 1627 46325 1639 46328
rect 1581 46319 1639 46325
rect 1670 46316 1676 46328
rect 1728 46316 1734 46368
rect 10962 46316 10968 46368
rect 11020 46316 11026 46368
rect 41233 46359 41291 46365
rect 41233 46325 41245 46359
rect 41279 46356 41291 46359
rect 41322 46356 41328 46368
rect 41279 46328 41328 46356
rect 41279 46325 41291 46328
rect 41233 46319 41291 46325
rect 41322 46316 41328 46328
rect 41380 46316 41386 46368
rect 48038 46356 48044 46368
rect 47999 46328 48044 46356
rect 48038 46316 48044 46328
rect 48096 46316 48102 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3970 46112 3976 46164
rect 4028 46152 4034 46164
rect 4341 46155 4399 46161
rect 4341 46152 4353 46155
rect 4028 46124 4353 46152
rect 4028 46112 4034 46124
rect 4341 46121 4353 46124
rect 4387 46121 4399 46155
rect 5074 46152 5080 46164
rect 5035 46124 5080 46152
rect 4341 46115 4399 46121
rect 5074 46112 5080 46124
rect 5132 46112 5138 46164
rect 13538 46152 13544 46164
rect 13499 46124 13544 46152
rect 13538 46112 13544 46124
rect 13596 46112 13602 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 20070 46152 20076 46164
rect 20031 46124 20076 46152
rect 20070 46112 20076 46124
rect 20128 46112 20134 46164
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 31849 46155 31907 46161
rect 31849 46121 31861 46155
rect 31895 46152 31907 46155
rect 32306 46152 32312 46164
rect 31895 46124 32312 46152
rect 31895 46121 31907 46124
rect 31849 46115 31907 46121
rect 32306 46112 32312 46124
rect 32364 46112 32370 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 42610 46112 42616 46164
rect 42668 46152 42674 46164
rect 43717 46155 43775 46161
rect 43717 46152 43729 46155
rect 42668 46124 43729 46152
rect 42668 46112 42674 46124
rect 43717 46121 43729 46124
rect 43763 46121 43775 46155
rect 43717 46115 43775 46121
rect 44361 46155 44419 46161
rect 44361 46121 44373 46155
rect 44407 46152 44419 46155
rect 45370 46152 45376 46164
rect 44407 46124 45376 46152
rect 44407 46121 44419 46124
rect 44361 46115 44419 46121
rect 45370 46112 45376 46124
rect 45428 46112 45434 46164
rect 6886 46056 24624 46084
rect 1762 45908 1768 45960
rect 1820 45948 1826 45960
rect 2041 45951 2099 45957
rect 2041 45948 2053 45951
rect 1820 45920 2053 45948
rect 1820 45908 1826 45920
rect 2041 45917 2053 45920
rect 2087 45917 2099 45951
rect 2041 45911 2099 45917
rect 4985 45951 5043 45957
rect 4985 45917 4997 45951
rect 5031 45948 5043 45951
rect 6886 45948 6914 46056
rect 20809 46019 20867 46025
rect 20809 45985 20821 46019
rect 20855 46016 20867 46019
rect 21082 46016 21088 46028
rect 20855 45988 21088 46016
rect 20855 45985 20867 45988
rect 20809 45979 20867 45985
rect 21082 45976 21088 45988
rect 21140 45976 21146 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 5031 45920 6914 45948
rect 5031 45917 5043 45920
rect 4985 45911 5043 45917
rect 12250 45908 12256 45960
rect 12308 45948 12314 45960
rect 12529 45951 12587 45957
rect 12529 45948 12541 45951
rect 12308 45920 12541 45948
rect 12308 45908 12314 45920
rect 12529 45917 12541 45920
rect 12575 45917 12587 45951
rect 14090 45948 14096 45960
rect 14003 45920 14096 45948
rect 12529 45911 12587 45917
rect 14090 45908 14096 45920
rect 14148 45948 14154 45960
rect 19981 45951 20039 45957
rect 19981 45948 19993 45951
rect 14148 45920 19993 45948
rect 14148 45908 14154 45920
rect 19981 45917 19993 45920
rect 20027 45948 20039 45951
rect 20622 45948 20628 45960
rect 20027 45920 20628 45948
rect 20027 45917 20039 45920
rect 19981 45911 20039 45917
rect 20622 45908 20628 45920
rect 20680 45908 20686 45960
rect 24596 45957 24624 46056
rect 39942 46044 39948 46096
rect 40000 46084 40006 46096
rect 40000 46056 44312 46084
rect 40000 46044 40006 46056
rect 25225 46019 25283 46025
rect 25225 45985 25237 46019
rect 25271 46016 25283 46019
rect 25498 46016 25504 46028
rect 25271 45988 25504 46016
rect 25271 45985 25283 45988
rect 25225 45979 25283 45985
rect 25498 45976 25504 45988
rect 25556 45976 25562 46028
rect 25774 46016 25780 46028
rect 25735 45988 25780 46016
rect 25774 45976 25780 45988
rect 25832 45976 25838 46028
rect 41322 46016 41328 46028
rect 41283 45988 41328 46016
rect 41322 45976 41328 45988
rect 41380 45976 41386 46028
rect 41874 46016 41880 46028
rect 41835 45988 41880 46016
rect 41874 45976 41880 45988
rect 41932 45976 41938 46028
rect 24581 45951 24639 45957
rect 24581 45917 24593 45951
rect 24627 45917 24639 45951
rect 31754 45948 31760 45960
rect 24581 45911 24639 45917
rect 29932 45920 31760 45948
rect 20993 45883 21051 45889
rect 20993 45849 21005 45883
rect 21039 45880 21051 45883
rect 21082 45880 21088 45892
rect 21039 45852 21088 45880
rect 21039 45849 21051 45852
rect 20993 45843 21051 45849
rect 21082 45840 21088 45852
rect 21140 45840 21146 45892
rect 12342 45812 12348 45824
rect 12303 45784 12348 45812
rect 12342 45772 12348 45784
rect 12400 45772 12406 45824
rect 24596 45812 24624 45911
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 29932 45880 29960 45920
rect 31754 45908 31760 45920
rect 31812 45908 31818 45960
rect 38197 45951 38255 45957
rect 38197 45917 38209 45951
rect 38243 45948 38255 45951
rect 39942 45948 39948 45960
rect 38243 45920 39948 45948
rect 38243 45917 38255 45920
rect 38197 45911 38255 45917
rect 39942 45908 39948 45920
rect 40000 45908 40006 45960
rect 44284 45957 44312 46056
rect 45738 46016 45744 46028
rect 45664 45988 45744 46016
rect 45664 45957 45692 45988
rect 45738 45976 45744 45988
rect 45796 45976 45802 46028
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 43625 45951 43683 45957
rect 43625 45917 43637 45951
rect 43671 45917 43683 45951
rect 43625 45911 43683 45917
rect 44269 45951 44327 45957
rect 44269 45917 44281 45951
rect 44315 45917 44327 45951
rect 44269 45911 44327 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45917 45707 45951
rect 46290 45948 46296 45960
rect 46251 45920 46296 45948
rect 45649 45911 45707 45917
rect 41506 45880 41512 45892
rect 26206 45852 29960 45880
rect 41467 45852 41512 45880
rect 26206 45812 26234 45852
rect 41506 45840 41512 45852
rect 41564 45840 41570 45892
rect 43640 45880 43668 45911
rect 46290 45908 46296 45920
rect 46348 45908 46354 45960
rect 45370 45880 45376 45892
rect 43640 45852 45376 45880
rect 45370 45840 45376 45852
rect 45428 45840 45434 45892
rect 45830 45880 45836 45892
rect 45791 45852 45836 45880
rect 45830 45840 45836 45852
rect 45888 45840 45894 45892
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 24596 45784 26234 45812
rect 45094 45772 45100 45824
rect 45152 45812 45158 45824
rect 45554 45812 45560 45824
rect 45152 45784 45560 45812
rect 45152 45772 45158 45784
rect 45554 45772 45560 45784
rect 45612 45772 45618 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 12066 45608 12072 45620
rect 12027 45580 12072 45608
rect 12066 45568 12072 45580
rect 12124 45568 12130 45620
rect 21082 45608 21088 45620
rect 21043 45580 21088 45608
rect 21082 45568 21088 45580
rect 21140 45568 21146 45620
rect 25406 45608 25412 45620
rect 25367 45580 25412 45608
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 41506 45608 41512 45620
rect 41467 45580 41512 45608
rect 41506 45568 41512 45580
rect 41564 45568 41570 45620
rect 46382 45568 46388 45620
rect 46440 45608 46446 45620
rect 46440 45580 47624 45608
rect 46440 45568 46446 45580
rect 42794 45500 42800 45552
rect 42852 45540 42858 45552
rect 42852 45512 44956 45540
rect 42852 45500 42858 45512
rect 1762 45472 1768 45484
rect 1723 45444 1768 45472
rect 1762 45432 1768 45444
rect 1820 45432 1826 45484
rect 11974 45472 11980 45484
rect 11935 45444 11980 45472
rect 11974 45432 11980 45444
rect 12032 45432 12038 45484
rect 20993 45475 21051 45481
rect 20993 45441 21005 45475
rect 21039 45472 21051 45475
rect 25317 45475 25375 45481
rect 25317 45472 25329 45475
rect 21039 45444 25329 45472
rect 21039 45441 21051 45444
rect 20993 45435 21051 45441
rect 25317 45441 25329 45444
rect 25363 45472 25375 45475
rect 27157 45475 27215 45481
rect 27157 45472 27169 45475
rect 25363 45444 27169 45472
rect 25363 45441 25375 45444
rect 25317 45435 25375 45441
rect 27157 45441 27169 45444
rect 27203 45472 27215 45475
rect 31018 45472 31024 45484
rect 27203 45444 31024 45472
rect 27203 45441 27215 45444
rect 27157 45435 27215 45441
rect 31018 45432 31024 45444
rect 31076 45432 31082 45484
rect 41414 45472 41420 45484
rect 41375 45444 41420 45472
rect 41414 45432 41420 45444
rect 41472 45432 41478 45484
rect 44928 45481 44956 45512
rect 47596 45481 47624 45580
rect 44913 45475 44971 45481
rect 44913 45441 44925 45475
rect 44959 45441 44971 45475
rect 44913 45435 44971 45441
rect 47581 45475 47639 45481
rect 47581 45441 47593 45475
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 1949 45407 2007 45413
rect 1949 45373 1961 45407
rect 1995 45404 2007 45407
rect 2222 45404 2228 45416
rect 1995 45376 2228 45404
rect 1995 45373 2007 45376
rect 1949 45367 2007 45373
rect 2222 45364 2228 45376
rect 2280 45364 2286 45416
rect 2774 45404 2780 45416
rect 2735 45376 2780 45404
rect 2774 45364 2780 45376
rect 2832 45364 2838 45416
rect 42613 45407 42671 45413
rect 42613 45373 42625 45407
rect 42659 45373 42671 45407
rect 42794 45404 42800 45416
rect 42755 45376 42800 45404
rect 42613 45367 42671 45373
rect 42628 45336 42656 45367
rect 42794 45364 42800 45376
rect 42852 45364 42858 45416
rect 44082 45404 44088 45416
rect 44043 45376 44088 45404
rect 44082 45364 44088 45376
rect 44140 45364 44146 45416
rect 45094 45404 45100 45416
rect 45055 45376 45100 45404
rect 45094 45364 45100 45376
rect 45152 45364 45158 45416
rect 45646 45404 45652 45416
rect 45607 45376 45652 45404
rect 45646 45364 45652 45376
rect 45704 45364 45710 45416
rect 43530 45336 43536 45348
rect 42628 45308 43536 45336
rect 43530 45296 43536 45308
rect 43588 45296 43594 45348
rect 27246 45268 27252 45280
rect 27207 45240 27252 45268
rect 27246 45228 27252 45240
rect 27304 45228 27310 45280
rect 47486 45228 47492 45280
rect 47544 45268 47550 45280
rect 47765 45271 47823 45277
rect 47765 45268 47777 45271
rect 47544 45240 47777 45268
rect 47544 45228 47550 45240
rect 47765 45237 47777 45240
rect 47811 45237 47823 45271
rect 47765 45231 47823 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 2222 45064 2228 45076
rect 2183 45036 2228 45064
rect 2222 45024 2228 45036
rect 2280 45024 2286 45076
rect 42794 45064 42800 45076
rect 42755 45036 42800 45064
rect 42794 45024 42800 45036
rect 42852 45024 42858 45076
rect 43530 45064 43536 45076
rect 43491 45036 43536 45064
rect 43530 45024 43536 45036
rect 43588 45024 43594 45076
rect 44361 45067 44419 45073
rect 44361 45033 44373 45067
rect 44407 45064 44419 45067
rect 45094 45064 45100 45076
rect 44407 45036 45100 45064
rect 44407 45033 44419 45036
rect 44361 45027 44419 45033
rect 45094 45024 45100 45036
rect 45152 45024 45158 45076
rect 45741 45067 45799 45073
rect 45741 45033 45753 45067
rect 45787 45064 45799 45067
rect 46474 45064 46480 45076
rect 45787 45036 46480 45064
rect 45787 45033 45799 45036
rect 45741 45027 45799 45033
rect 46474 45024 46480 45036
rect 46532 45024 46538 45076
rect 45189 44999 45247 45005
rect 45189 44965 45201 44999
rect 45235 44996 45247 44999
rect 46290 44996 46296 45008
rect 45235 44968 46296 44996
rect 45235 44965 45247 44968
rect 45189 44959 45247 44965
rect 46290 44956 46296 44968
rect 46348 44956 46354 45008
rect 27246 44928 27252 44940
rect 27207 44900 27252 44928
rect 27246 44888 27252 44900
rect 27304 44888 27310 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 2133 44863 2191 44869
rect 2133 44829 2145 44863
rect 2179 44860 2191 44863
rect 2314 44860 2320 44872
rect 2179 44832 2320 44860
rect 2179 44829 2191 44832
rect 2133 44823 2191 44829
rect 2314 44820 2320 44832
rect 2372 44820 2378 44872
rect 27062 44860 27068 44872
rect 27023 44832 27068 44860
rect 27062 44820 27068 44832
rect 27120 44820 27126 44872
rect 42705 44863 42763 44869
rect 42705 44829 42717 44863
rect 42751 44829 42763 44863
rect 42705 44823 42763 44829
rect 44269 44863 44327 44869
rect 44269 44829 44281 44863
rect 44315 44860 44327 44863
rect 45002 44860 45008 44872
rect 44315 44832 45008 44860
rect 44315 44829 44327 44832
rect 44269 44823 44327 44829
rect 28905 44795 28963 44801
rect 28905 44761 28917 44795
rect 28951 44792 28963 44795
rect 38654 44792 38660 44804
rect 28951 44764 38660 44792
rect 28951 44761 28963 44764
rect 28905 44755 28963 44761
rect 38654 44752 38660 44764
rect 38712 44752 38718 44804
rect 42720 44792 42748 44823
rect 45002 44820 45008 44832
rect 45060 44820 45066 44872
rect 45370 44820 45376 44872
rect 45428 44860 45434 44872
rect 45649 44863 45707 44869
rect 45649 44860 45661 44863
rect 45428 44832 45661 44860
rect 45428 44820 45434 44832
rect 45649 44829 45661 44832
rect 45695 44829 45707 44863
rect 45649 44823 45707 44829
rect 46293 44863 46351 44869
rect 46293 44829 46305 44863
rect 46339 44829 46351 44863
rect 46293 44823 46351 44829
rect 46198 44792 46204 44804
rect 42720 44764 46204 44792
rect 46198 44752 46204 44764
rect 46256 44752 46262 44804
rect 46308 44724 46336 44823
rect 46474 44792 46480 44804
rect 46435 44764 46480 44792
rect 46474 44752 46480 44764
rect 46532 44752 46538 44804
rect 47026 44724 47032 44736
rect 46308 44696 47032 44724
rect 47026 44684 47032 44696
rect 47084 44684 47090 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 27062 44520 27068 44532
rect 27023 44492 27068 44520
rect 27062 44480 27068 44492
rect 27120 44480 27126 44532
rect 46293 44523 46351 44529
rect 46293 44489 46305 44523
rect 46339 44520 46351 44523
rect 46474 44520 46480 44532
rect 46339 44492 46480 44520
rect 46339 44489 46351 44492
rect 46293 44483 46351 44489
rect 46474 44480 46480 44492
rect 46532 44480 46538 44532
rect 45462 44412 45468 44464
rect 45520 44452 45526 44464
rect 47673 44455 47731 44461
rect 47673 44452 47685 44455
rect 45520 44424 47685 44452
rect 45520 44412 45526 44424
rect 47673 44421 47685 44424
rect 47719 44421 47731 44455
rect 47673 44415 47731 44421
rect 25130 44344 25136 44396
rect 25188 44384 25194 44396
rect 26973 44387 27031 44393
rect 26973 44384 26985 44387
rect 25188 44356 26985 44384
rect 25188 44344 25194 44356
rect 26973 44353 26985 44356
rect 27019 44353 27031 44387
rect 26973 44347 27031 44353
rect 45097 44387 45155 44393
rect 45097 44353 45109 44387
rect 45143 44384 45155 44387
rect 45186 44384 45192 44396
rect 45143 44356 45192 44384
rect 45143 44353 45155 44356
rect 45097 44347 45155 44353
rect 45186 44344 45192 44356
rect 45244 44344 45250 44396
rect 45738 44384 45744 44396
rect 45699 44356 45744 44384
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46201 44387 46259 44393
rect 46201 44353 46213 44387
rect 46247 44384 46259 44387
rect 46845 44387 46903 44393
rect 46845 44384 46857 44387
rect 46247 44356 46857 44384
rect 46247 44353 46259 44356
rect 46201 44347 46259 44353
rect 46845 44353 46857 44356
rect 46891 44353 46903 44387
rect 47578 44384 47584 44396
rect 47539 44356 47584 44384
rect 46845 44347 46903 44353
rect 41414 44276 41420 44328
rect 41472 44316 41478 44328
rect 46216 44316 46244 44347
rect 47578 44344 47584 44356
rect 47636 44344 47642 44396
rect 41472 44288 46244 44316
rect 41472 44276 41478 44288
rect 46934 44180 46940 44192
rect 46895 44152 46940 44180
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 46934 43840 46940 43852
rect 46523 43812 46940 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 46934 43800 46940 43812
rect 46992 43800 46998 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 1673 43231 1731 43237
rect 1673 43197 1685 43231
rect 1719 43228 1731 43231
rect 41230 43228 41236 43240
rect 1719 43200 41236 43228
rect 1719 43197 1731 43200
rect 1673 43191 1731 43197
rect 41230 43188 41236 43200
rect 41288 43188 41294 43240
rect 47762 43092 47768 43104
rect 47723 43064 47768 43092
rect 47762 43052 47768 43064
rect 47820 43052 47826 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46293 42755 46351 42761
rect 46293 42721 46305 42755
rect 46339 42752 46351 42755
rect 47762 42752 47768 42764
rect 46339 42724 47768 42752
rect 46339 42721 46351 42724
rect 46293 42715 46351 42721
rect 47762 42712 47768 42724
rect 47820 42712 47826 42764
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 46934 42616 46940 42628
rect 46523 42588 46940 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 46934 42576 46940 42588
rect 46992 42576 46998 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 46934 42344 46940 42356
rect 46895 42316 46940 42344
rect 46934 42304 46940 42316
rect 46992 42304 46998 42356
rect 44358 42236 44364 42288
rect 44416 42276 44422 42288
rect 45370 42276 45376 42288
rect 44416 42248 45376 42276
rect 44416 42236 44422 42248
rect 45370 42236 45376 42248
rect 45428 42276 45434 42288
rect 45428 42248 47624 42276
rect 45428 42236 45434 42248
rect 46198 42168 46204 42220
rect 46256 42208 46262 42220
rect 46658 42208 46664 42220
rect 46256 42180 46664 42208
rect 46256 42168 46262 42180
rect 46658 42168 46664 42180
rect 46716 42208 46722 42220
rect 47596 42217 47624 42248
rect 46845 42211 46903 42217
rect 46845 42208 46857 42211
rect 46716 42180 46857 42208
rect 46716 42168 46722 42180
rect 46845 42177 46857 42180
rect 46891 42177 46903 42211
rect 46845 42171 46903 42177
rect 47581 42211 47639 42217
rect 47581 42177 47593 42211
rect 47627 42177 47639 42211
rect 47581 42171 47639 42177
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 46474 41964 46480 42016
rect 46532 42004 46538 42016
rect 47673 42007 47731 42013
rect 47673 42004 47685 42007
rect 46532 41976 47685 42004
rect 46532 41964 46538 41976
rect 47673 41973 47685 41976
rect 47719 41973 47731 42007
rect 47673 41967 47731 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46474 41664 46480 41676
rect 46435 41636 46480 41664
rect 46474 41624 46480 41636
rect 46532 41624 46538 41676
rect 46293 41599 46351 41605
rect 46293 41565 46305 41599
rect 46339 41565 46351 41599
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 46293 41559 46351 41565
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46308 41528 46336 41559
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 47670 41528 47676 41540
rect 46308 41500 47676 41528
rect 47670 41488 47676 41500
rect 47728 41488 47734 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 2133 41219 2191 41225
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 47302 40876 47308 40928
rect 47360 40916 47366 40928
rect 48041 40919 48099 40925
rect 48041 40916 48053 40919
rect 47360 40888 48053 40916
rect 47360 40876 47366 40888
rect 48041 40885 48053 40888
rect 48087 40885 48099 40919
rect 48041 40879 48099 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 22281 40511 22339 40517
rect 22281 40477 22293 40511
rect 22327 40508 22339 40511
rect 22922 40508 22928 40520
rect 22327 40480 22928 40508
rect 22327 40477 22339 40480
rect 22281 40471 22339 40477
rect 22922 40468 22928 40480
rect 22980 40468 22986 40520
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 1949 40375 2007 40381
rect 1949 40341 1961 40375
rect 1995 40372 2007 40375
rect 10318 40372 10324 40384
rect 1995 40344 10324 40372
rect 1995 40341 2007 40344
rect 1949 40335 2007 40341
rect 10318 40332 10324 40344
rect 10376 40332 10382 40384
rect 22094 40332 22100 40384
rect 22152 40372 22158 40384
rect 22152 40344 22197 40372
rect 22152 40332 22158 40344
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 22922 40168 22928 40180
rect 22883 40140 22928 40168
rect 22922 40128 22928 40140
rect 22980 40128 22986 40180
rect 20346 40100 20352 40112
rect 20307 40072 20352 40100
rect 20346 40060 20352 40072
rect 20404 40060 20410 40112
rect 20530 40100 20536 40112
rect 20491 40072 20536 40100
rect 20530 40060 20536 40072
rect 20588 40060 20594 40112
rect 45830 40100 45836 40112
rect 24044 40072 45836 40100
rect 24044 40041 24072 40072
rect 45830 40060 45836 40072
rect 45888 40060 45894 40112
rect 22281 40035 22339 40041
rect 22281 40001 22293 40035
rect 22327 40032 22339 40035
rect 22649 40035 22707 40041
rect 22649 40032 22661 40035
rect 22327 40004 22661 40032
rect 22327 40001 22339 40004
rect 22281 39995 22339 40001
rect 22649 40001 22661 40004
rect 22695 40032 22707 40035
rect 23293 40035 23351 40041
rect 23293 40032 23305 40035
rect 22695 40004 23305 40032
rect 22695 40001 22707 40004
rect 22649 39995 22707 40001
rect 23293 40001 23305 40004
rect 23339 40032 23351 40035
rect 24029 40035 24087 40041
rect 24029 40032 24041 40035
rect 23339 40004 24041 40032
rect 23339 40001 23351 40004
rect 23293 39995 23351 40001
rect 24029 40001 24041 40004
rect 24075 40001 24087 40035
rect 24029 39995 24087 40001
rect 23106 39924 23112 39976
rect 23164 39964 23170 39976
rect 23385 39967 23443 39973
rect 23385 39964 23397 39967
rect 23164 39936 23397 39964
rect 23164 39924 23170 39936
rect 23385 39933 23397 39936
rect 23431 39933 23443 39967
rect 23385 39927 23443 39933
rect 23477 39967 23535 39973
rect 23477 39933 23489 39967
rect 23523 39933 23535 39967
rect 23477 39927 23535 39933
rect 20530 39856 20536 39908
rect 20588 39896 20594 39908
rect 23492 39896 23520 39927
rect 20588 39868 23520 39896
rect 20588 39856 20594 39868
rect 20346 39788 20352 39840
rect 20404 39828 20410 39840
rect 20717 39831 20775 39837
rect 20717 39828 20729 39831
rect 20404 39800 20729 39828
rect 20404 39788 20410 39800
rect 20717 39797 20729 39800
rect 20763 39797 20775 39831
rect 20717 39791 20775 39797
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 21637 39491 21695 39497
rect 21637 39457 21649 39491
rect 21683 39488 21695 39491
rect 22094 39488 22100 39500
rect 21683 39460 22100 39488
rect 21683 39457 21695 39460
rect 21637 39451 21695 39457
rect 22094 39448 22100 39460
rect 22152 39448 22158 39500
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 19889 39423 19947 39429
rect 19889 39389 19901 39423
rect 19935 39420 19947 39423
rect 19978 39420 19984 39432
rect 19935 39392 19984 39420
rect 19935 39389 19947 39392
rect 19889 39383 19947 39389
rect 19978 39380 19984 39392
rect 20036 39380 20042 39432
rect 21358 39420 21364 39432
rect 21319 39392 21364 39420
rect 21358 39380 21364 39392
rect 21416 39380 21422 39432
rect 45002 39420 45008 39432
rect 44963 39392 45008 39420
rect 45002 39380 45008 39392
rect 45060 39380 45066 39432
rect 22094 39312 22100 39364
rect 22152 39312 22158 39364
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 46934 39352 46940 39364
rect 46523 39324 46940 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 46934 39312 46940 39324
rect 46992 39312 46998 39364
rect 20073 39287 20131 39293
rect 20073 39253 20085 39287
rect 20119 39284 20131 39287
rect 20254 39284 20260 39296
rect 20119 39256 20260 39284
rect 20119 39253 20131 39256
rect 20073 39247 20131 39253
rect 20254 39244 20260 39256
rect 20312 39244 20318 39296
rect 22922 39244 22928 39296
rect 22980 39284 22986 39296
rect 23109 39287 23167 39293
rect 23109 39284 23121 39287
rect 22980 39256 23121 39284
rect 22980 39244 22986 39256
rect 23109 39253 23121 39256
rect 23155 39253 23167 39287
rect 23109 39247 23167 39253
rect 45097 39287 45155 39293
rect 45097 39253 45109 39287
rect 45143 39284 45155 39287
rect 45186 39284 45192 39296
rect 45143 39256 45192 39284
rect 45143 39253 45155 39256
rect 45097 39247 45155 39253
rect 45186 39244 45192 39256
rect 45244 39244 45250 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 20257 39083 20315 39089
rect 20257 39049 20269 39083
rect 20303 39049 20315 39083
rect 20257 39043 20315 39049
rect 22005 39083 22063 39089
rect 22005 39049 22017 39083
rect 22051 39080 22063 39083
rect 22094 39080 22100 39092
rect 22051 39052 22100 39080
rect 22051 39049 22063 39052
rect 22005 39043 22063 39049
rect 20272 39012 20300 39043
rect 22094 39040 22100 39052
rect 22152 39040 22158 39092
rect 23106 39080 23112 39092
rect 23067 39052 23112 39080
rect 23106 39040 23112 39052
rect 23164 39040 23170 39092
rect 45186 39012 45192 39024
rect 20272 38984 22094 39012
rect 45147 38984 45192 39012
rect 19334 38904 19340 38956
rect 19392 38944 19398 38956
rect 19978 38944 19984 38956
rect 19392 38916 19984 38944
rect 19392 38904 19398 38916
rect 19978 38904 19984 38916
rect 20036 38944 20042 38956
rect 20073 38947 20131 38953
rect 20073 38944 20085 38947
rect 20036 38916 20085 38944
rect 20036 38904 20042 38916
rect 20073 38913 20085 38916
rect 20119 38913 20131 38947
rect 20073 38907 20131 38913
rect 20254 38904 20260 38956
rect 20312 38944 20318 38956
rect 21913 38947 21971 38953
rect 21913 38944 21925 38947
rect 20312 38916 21925 38944
rect 20312 38904 20318 38916
rect 21913 38913 21925 38916
rect 21959 38913 21971 38947
rect 21913 38907 21971 38913
rect 20438 38768 20444 38820
rect 20496 38808 20502 38820
rect 22066 38808 22094 38984
rect 45186 38972 45192 38984
rect 45244 38972 45250 39024
rect 46842 39012 46848 39024
rect 46803 38984 46848 39012
rect 46842 38972 46848 38984
rect 46900 38972 46906 39024
rect 22741 38947 22799 38953
rect 22741 38913 22753 38947
rect 22787 38944 22799 38947
rect 22922 38944 22928 38956
rect 22787 38916 22928 38944
rect 22787 38913 22799 38916
rect 22741 38907 22799 38913
rect 22922 38904 22928 38916
rect 22980 38904 22986 38956
rect 23569 38947 23627 38953
rect 23569 38913 23581 38947
rect 23615 38944 23627 38947
rect 27801 38947 27859 38953
rect 27801 38944 27813 38947
rect 23615 38916 27813 38944
rect 23615 38913 23627 38916
rect 23569 38907 23627 38913
rect 27801 38913 27813 38916
rect 27847 38944 27859 38947
rect 28810 38944 28816 38956
rect 27847 38916 28816 38944
rect 27847 38913 27859 38916
rect 27801 38907 27859 38913
rect 22554 38836 22560 38888
rect 22612 38876 22618 38888
rect 22649 38879 22707 38885
rect 22649 38876 22661 38879
rect 22612 38848 22661 38876
rect 22612 38836 22618 38848
rect 22649 38845 22661 38848
rect 22695 38845 22707 38879
rect 22649 38839 22707 38845
rect 23584 38808 23612 38907
rect 28810 38904 28816 38916
rect 28868 38904 28874 38956
rect 43622 38944 43628 38956
rect 43583 38916 43628 38944
rect 43622 38904 43628 38916
rect 43680 38904 43686 38956
rect 47762 38944 47768 38956
rect 47723 38916 47768 38944
rect 47762 38904 47768 38916
rect 47820 38904 47826 38956
rect 44358 38876 44364 38888
rect 44319 38848 44364 38876
rect 44358 38836 44364 38848
rect 44416 38836 44422 38888
rect 44634 38836 44640 38888
rect 44692 38876 44698 38888
rect 45005 38879 45063 38885
rect 45005 38876 45017 38879
rect 44692 38848 45017 38876
rect 44692 38836 44698 38848
rect 45005 38845 45017 38848
rect 45051 38845 45063 38879
rect 45005 38839 45063 38845
rect 20496 38780 23612 38808
rect 20496 38768 20502 38780
rect 23474 38700 23480 38752
rect 23532 38740 23538 38752
rect 23661 38743 23719 38749
rect 23661 38740 23673 38743
rect 23532 38712 23673 38740
rect 23532 38700 23538 38712
rect 23661 38709 23673 38712
rect 23707 38709 23719 38743
rect 27890 38740 27896 38752
rect 27851 38712 27896 38740
rect 23661 38703 23719 38709
rect 27890 38700 27896 38712
rect 27948 38700 27954 38752
rect 47026 38700 47032 38752
rect 47084 38740 47090 38752
rect 47857 38743 47915 38749
rect 47857 38740 47869 38743
rect 47084 38712 47869 38740
rect 47084 38700 47090 38712
rect 47857 38709 47869 38712
rect 47903 38709 47915 38743
rect 47857 38703 47915 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 27338 38536 27344 38548
rect 17236 38508 27344 38536
rect 12342 38292 12348 38344
rect 12400 38332 12406 38344
rect 16301 38335 16359 38341
rect 16301 38332 16313 38335
rect 12400 38304 16313 38332
rect 12400 38292 12406 38304
rect 16301 38301 16313 38304
rect 16347 38301 16359 38335
rect 16482 38332 16488 38344
rect 16443 38304 16488 38332
rect 16301 38295 16359 38301
rect 16482 38292 16488 38304
rect 16540 38292 16546 38344
rect 11974 38224 11980 38276
rect 12032 38264 12038 38276
rect 17236 38264 17264 38508
rect 27338 38496 27344 38508
rect 27396 38496 27402 38548
rect 46934 38536 46940 38548
rect 46895 38508 46940 38536
rect 46934 38496 46940 38508
rect 46992 38496 46998 38548
rect 19521 38403 19579 38409
rect 19521 38369 19533 38403
rect 19567 38400 19579 38403
rect 20806 38400 20812 38412
rect 19567 38372 20812 38400
rect 19567 38369 19579 38372
rect 19521 38363 19579 38369
rect 20806 38360 20812 38372
rect 20864 38400 20870 38412
rect 21358 38400 21364 38412
rect 20864 38372 21364 38400
rect 20864 38360 20870 38372
rect 21358 38360 21364 38372
rect 21416 38400 21422 38412
rect 21913 38403 21971 38409
rect 21913 38400 21925 38403
rect 21416 38372 21925 38400
rect 21416 38360 21422 38372
rect 21913 38369 21925 38372
rect 21959 38369 21971 38403
rect 21913 38363 21971 38369
rect 24397 38403 24455 38409
rect 24397 38369 24409 38403
rect 24443 38400 24455 38403
rect 26605 38403 26663 38409
rect 26605 38400 26617 38403
rect 24443 38372 26617 38400
rect 24443 38369 24455 38372
rect 24397 38363 24455 38369
rect 26605 38369 26617 38372
rect 26651 38400 26663 38403
rect 27614 38400 27620 38412
rect 26651 38372 27620 38400
rect 26651 38369 26663 38372
rect 26605 38363 26663 38369
rect 27614 38360 27620 38372
rect 27672 38360 27678 38412
rect 39114 38360 39120 38412
rect 39172 38400 39178 38412
rect 39942 38400 39948 38412
rect 39172 38372 39948 38400
rect 39172 38360 39178 38372
rect 39942 38360 39948 38372
rect 40000 38400 40006 38412
rect 44269 38403 44327 38409
rect 44269 38400 44281 38403
rect 40000 38372 44281 38400
rect 40000 38360 40006 38372
rect 44269 38369 44281 38372
rect 44315 38369 44327 38403
rect 44269 38363 44327 38369
rect 43533 38335 43591 38341
rect 43533 38301 43545 38335
rect 43579 38332 43591 38335
rect 43622 38332 43628 38344
rect 43579 38304 43628 38332
rect 43579 38301 43591 38304
rect 43533 38295 43591 38301
rect 43622 38292 43628 38304
rect 43680 38332 43686 38344
rect 45005 38335 45063 38341
rect 45005 38332 45017 38335
rect 43680 38304 45017 38332
rect 43680 38292 43686 38304
rect 45005 38301 45017 38304
rect 45051 38301 45063 38335
rect 45005 38295 45063 38301
rect 46566 38292 46572 38344
rect 46624 38332 46630 38344
rect 46845 38335 46903 38341
rect 46845 38332 46857 38335
rect 46624 38304 46857 38332
rect 46624 38292 46630 38304
rect 46845 38301 46857 38304
rect 46891 38301 46903 38335
rect 46845 38295 46903 38301
rect 12032 38236 17264 38264
rect 19797 38267 19855 38273
rect 12032 38224 12038 38236
rect 19797 38233 19809 38267
rect 19843 38233 19855 38267
rect 19797 38227 19855 38233
rect 16393 38199 16451 38205
rect 16393 38165 16405 38199
rect 16439 38196 16451 38199
rect 18966 38196 18972 38208
rect 16439 38168 18972 38196
rect 16439 38165 16451 38168
rect 16393 38159 16451 38165
rect 18966 38156 18972 38168
rect 19024 38156 19030 38208
rect 19812 38196 19840 38227
rect 20530 38224 20536 38276
rect 20588 38224 20594 38276
rect 22186 38264 22192 38276
rect 22147 38236 22192 38264
rect 22186 38224 22192 38236
rect 22244 38224 22250 38276
rect 23474 38264 23480 38276
rect 23414 38236 23480 38264
rect 23474 38224 23480 38236
rect 23532 38224 23538 38276
rect 24673 38267 24731 38273
rect 24673 38233 24685 38267
rect 24719 38264 24731 38267
rect 24762 38264 24768 38276
rect 24719 38236 24768 38264
rect 24719 38233 24731 38236
rect 24673 38227 24731 38233
rect 24762 38224 24768 38236
rect 24820 38224 24826 38276
rect 25682 38224 25688 38276
rect 25740 38224 25746 38276
rect 26881 38267 26939 38273
rect 26881 38233 26893 38267
rect 26927 38264 26939 38267
rect 26970 38264 26976 38276
rect 26927 38236 26976 38264
rect 26927 38233 26939 38236
rect 26881 38227 26939 38233
rect 26970 38224 26976 38236
rect 27028 38224 27034 38276
rect 27890 38224 27896 38276
rect 27948 38224 27954 38276
rect 45922 38264 45928 38276
rect 45883 38236 45928 38264
rect 45922 38224 45928 38236
rect 45980 38224 45986 38276
rect 19978 38196 19984 38208
rect 19812 38168 19984 38196
rect 19978 38156 19984 38168
rect 20036 38156 20042 38208
rect 21266 38196 21272 38208
rect 21227 38168 21272 38196
rect 21266 38156 21272 38168
rect 21324 38156 21330 38208
rect 22830 38156 22836 38208
rect 22888 38196 22894 38208
rect 23198 38196 23204 38208
rect 22888 38168 23204 38196
rect 22888 38156 22894 38168
rect 23198 38156 23204 38168
rect 23256 38196 23262 38208
rect 23661 38199 23719 38205
rect 23661 38196 23673 38199
rect 23256 38168 23673 38196
rect 23256 38156 23262 38168
rect 23661 38165 23673 38168
rect 23707 38165 23719 38199
rect 23661 38159 23719 38165
rect 25958 38156 25964 38208
rect 26016 38196 26022 38208
rect 26145 38199 26203 38205
rect 26145 38196 26157 38199
rect 26016 38168 26157 38196
rect 26016 38156 26022 38168
rect 26145 38165 26157 38168
rect 26191 38165 26203 38199
rect 28350 38196 28356 38208
rect 28311 38168 28356 38196
rect 26145 38159 26203 38165
rect 28350 38156 28356 38168
rect 28408 38156 28414 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 17494 37992 17500 38004
rect 6886 37964 17500 37992
rect 2314 37884 2320 37936
rect 2372 37924 2378 37936
rect 6886 37924 6914 37964
rect 17494 37952 17500 37964
rect 17552 37952 17558 38004
rect 17589 37995 17647 38001
rect 17589 37961 17601 37995
rect 17635 37992 17647 37995
rect 18506 37992 18512 38004
rect 17635 37964 18512 37992
rect 17635 37961 17647 37964
rect 17589 37955 17647 37961
rect 18506 37952 18512 37964
rect 18564 37952 18570 38004
rect 18690 37992 18696 38004
rect 18651 37964 18696 37992
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 20530 37952 20536 38004
rect 20588 37992 20594 38004
rect 20625 37995 20683 38001
rect 20625 37992 20637 37995
rect 20588 37964 20637 37992
rect 20588 37952 20594 37964
rect 20625 37961 20637 37964
rect 20671 37961 20683 37995
rect 24762 37992 24768 38004
rect 24723 37964 24768 37992
rect 20625 37955 20683 37961
rect 24762 37952 24768 37964
rect 24820 37952 24826 38004
rect 25593 37995 25651 38001
rect 25593 37961 25605 37995
rect 25639 37992 25651 37995
rect 25682 37992 25688 38004
rect 25639 37964 25688 37992
rect 25639 37961 25651 37964
rect 25593 37955 25651 37961
rect 25682 37952 25688 37964
rect 25740 37952 25746 38004
rect 26970 37992 26976 38004
rect 26931 37964 26976 37992
rect 26970 37952 26976 37964
rect 27028 37952 27034 38004
rect 2372 37896 6914 37924
rect 2372 37884 2378 37896
rect 17678 37884 17684 37936
rect 17736 37924 17742 37936
rect 19242 37924 19248 37936
rect 17736 37896 19248 37924
rect 17736 37884 17742 37896
rect 19242 37884 19248 37896
rect 19300 37884 19306 37936
rect 19705 37927 19763 37933
rect 19705 37893 19717 37927
rect 19751 37924 19763 37927
rect 19794 37924 19800 37936
rect 19751 37896 19800 37924
rect 19751 37893 19763 37896
rect 19705 37887 19763 37893
rect 19794 37884 19800 37896
rect 19852 37884 19858 37936
rect 20162 37884 20168 37936
rect 20220 37924 20226 37936
rect 45922 37924 45928 37936
rect 20220 37896 45928 37924
rect 20220 37884 20226 37896
rect 45922 37884 45928 37896
rect 45980 37884 45986 37936
rect 17310 37816 17316 37868
rect 17368 37856 17374 37868
rect 17405 37859 17463 37865
rect 17405 37856 17417 37859
rect 17368 37828 17417 37856
rect 17368 37816 17374 37828
rect 17405 37825 17417 37828
rect 17451 37825 17463 37859
rect 18138 37856 18144 37868
rect 17691 37849 17749 37855
rect 17691 37846 17703 37849
rect 17405 37819 17463 37825
rect 17512 37818 17703 37846
rect 14458 37748 14464 37800
rect 14516 37788 14522 37800
rect 17512 37788 17540 37818
rect 17691 37815 17703 37818
rect 17737 37815 17749 37849
rect 18099 37828 18144 37856
rect 18138 37816 18144 37828
rect 18196 37816 18202 37868
rect 18325 37859 18383 37865
rect 18325 37825 18337 37859
rect 18371 37825 18383 37859
rect 18325 37819 18383 37825
rect 17691 37809 17749 37815
rect 14516 37760 17540 37788
rect 18340 37788 18368 37819
rect 18414 37816 18420 37868
rect 18472 37856 18478 37868
rect 18555 37859 18613 37865
rect 19426 37860 19432 37868
rect 18472 37828 18517 37856
rect 18472 37816 18478 37828
rect 18555 37825 18567 37859
rect 18601 37856 18613 37859
rect 19352 37856 19432 37860
rect 18601 37832 19432 37856
rect 18601 37828 19380 37832
rect 18601 37825 18613 37828
rect 18555 37819 18613 37825
rect 19426 37816 19432 37832
rect 19484 37816 19490 37868
rect 19993 37859 20051 37865
rect 19601 37849 19659 37855
rect 19601 37846 19613 37849
rect 19536 37840 19613 37846
rect 19524 37818 19613 37840
rect 19524 37812 19564 37818
rect 19601 37815 19613 37818
rect 19647 37815 19659 37849
rect 19993 37825 20005 37859
rect 20039 37856 20051 37859
rect 20039 37828 20208 37856
rect 20039 37825 20051 37828
rect 19993 37819 20051 37825
rect 19288 37788 19294 37800
rect 18340 37760 19294 37788
rect 14516 37748 14522 37760
rect 19288 37748 19294 37760
rect 19346 37748 19352 37800
rect 9490 37680 9496 37732
rect 9548 37720 9554 37732
rect 14366 37720 14372 37732
rect 9548 37692 14372 37720
rect 9548 37680 9554 37692
rect 14366 37680 14372 37692
rect 14424 37680 14430 37732
rect 16850 37612 16856 37664
rect 16908 37652 16914 37664
rect 17221 37655 17279 37661
rect 17221 37652 17233 37655
rect 16908 37624 17233 37652
rect 16908 37612 16914 37624
rect 17221 37621 17233 37624
rect 17267 37621 17279 37655
rect 17221 37615 17279 37621
rect 18506 37612 18512 37664
rect 18564 37652 18570 37664
rect 19242 37652 19248 37664
rect 18564 37624 19248 37652
rect 18564 37612 18570 37624
rect 19242 37612 19248 37624
rect 19300 37612 19306 37664
rect 19524 37652 19552 37812
rect 19601 37809 19659 37815
rect 20180 37800 20208 37828
rect 20438 37816 20444 37868
rect 20496 37856 20502 37868
rect 20533 37859 20591 37865
rect 20533 37856 20545 37859
rect 20496 37828 20545 37856
rect 20496 37816 20502 37828
rect 20533 37825 20545 37828
rect 20579 37825 20591 37859
rect 22830 37856 22836 37868
rect 22791 37828 22836 37856
rect 20533 37819 20591 37825
rect 22830 37816 22836 37828
rect 22888 37816 22894 37868
rect 23014 37816 23020 37868
rect 23072 37856 23078 37868
rect 23109 37859 23167 37865
rect 23109 37856 23121 37859
rect 23072 37828 23121 37856
rect 23072 37816 23078 37828
rect 23109 37825 23121 37828
rect 23155 37825 23167 37859
rect 23109 37819 23167 37825
rect 23198 37816 23204 37868
rect 23256 37856 23262 37868
rect 23753 37859 23811 37865
rect 23753 37856 23765 37859
rect 23256 37828 23765 37856
rect 23256 37816 23262 37828
rect 23753 37825 23765 37828
rect 23799 37825 23811 37859
rect 24946 37856 24952 37868
rect 24907 37828 24952 37856
rect 23753 37819 23811 37825
rect 24946 37816 24952 37828
rect 25004 37816 25010 37868
rect 25501 37859 25559 37865
rect 25501 37825 25513 37859
rect 25547 37856 25559 37859
rect 26970 37856 26976 37868
rect 25547 37828 26976 37856
rect 25547 37825 25559 37828
rect 25501 37819 25559 37825
rect 26970 37816 26976 37828
rect 27028 37816 27034 37868
rect 27154 37856 27160 37868
rect 27115 37828 27160 37856
rect 27154 37816 27160 37828
rect 27212 37816 27218 37868
rect 27249 37859 27307 37865
rect 27249 37825 27261 37859
rect 27295 37825 27307 37859
rect 27522 37856 27528 37868
rect 27483 37828 27528 37856
rect 27249 37819 27307 37825
rect 19819 37791 19877 37797
rect 19819 37788 19831 37791
rect 19720 37760 19831 37788
rect 19610 37680 19616 37732
rect 19668 37720 19674 37732
rect 19720 37720 19748 37760
rect 19819 37757 19831 37760
rect 19865 37757 19877 37791
rect 19819 37751 19877 37757
rect 20162 37748 20168 37800
rect 20220 37748 20226 37800
rect 22738 37748 22744 37800
rect 22796 37788 22802 37800
rect 22925 37791 22983 37797
rect 22925 37788 22937 37791
rect 22796 37760 22937 37788
rect 22796 37748 22802 37760
rect 22925 37757 22937 37760
rect 22971 37788 22983 37791
rect 25958 37788 25964 37800
rect 22971 37760 25964 37788
rect 22971 37757 22983 37760
rect 22925 37751 22983 37757
rect 25958 37748 25964 37760
rect 26016 37748 26022 37800
rect 27062 37748 27068 37800
rect 27120 37788 27126 37800
rect 27264 37788 27292 37819
rect 27522 37816 27528 37828
rect 27580 37816 27586 37868
rect 43622 37816 43628 37868
rect 43680 37856 43686 37868
rect 44085 37859 44143 37865
rect 44085 37856 44097 37859
rect 43680 37828 44097 37856
rect 43680 37816 43686 37828
rect 44085 37825 44097 37828
rect 44131 37856 44143 37859
rect 44266 37856 44272 37868
rect 44131 37828 44272 37856
rect 44131 37825 44143 37828
rect 44085 37819 44143 37825
rect 44266 37816 44272 37828
rect 44324 37816 44330 37868
rect 27120 37760 27292 37788
rect 27120 37748 27126 37760
rect 27338 37748 27344 37800
rect 27396 37788 27402 37800
rect 44453 37791 44511 37797
rect 44453 37788 44465 37791
rect 27396 37760 44465 37788
rect 27396 37748 27402 37760
rect 44453 37757 44465 37760
rect 44499 37788 44511 37791
rect 44910 37788 44916 37800
rect 44499 37760 44916 37788
rect 44499 37757 44511 37760
rect 44453 37751 44511 37757
rect 44910 37748 44916 37760
rect 44968 37748 44974 37800
rect 19978 37720 19984 37732
rect 19668 37692 19748 37720
rect 19939 37692 19984 37720
rect 19668 37680 19674 37692
rect 19978 37680 19984 37692
rect 20036 37680 20042 37732
rect 20898 37652 20904 37664
rect 19524 37624 20904 37652
rect 20898 37612 20904 37624
rect 20956 37612 20962 37664
rect 21266 37612 21272 37664
rect 21324 37652 21330 37664
rect 22833 37655 22891 37661
rect 22833 37652 22845 37655
rect 21324 37624 22845 37652
rect 21324 37612 21330 37624
rect 22833 37621 22845 37624
rect 22879 37652 22891 37655
rect 23198 37652 23204 37664
rect 22879 37624 23204 37652
rect 22879 37621 22891 37624
rect 22833 37615 22891 37621
rect 23198 37612 23204 37624
rect 23256 37612 23262 37664
rect 23290 37612 23296 37664
rect 23348 37652 23354 37664
rect 23348 37624 23393 37652
rect 23348 37612 23354 37624
rect 23566 37612 23572 37664
rect 23624 37652 23630 37664
rect 23845 37655 23903 37661
rect 23845 37652 23857 37655
rect 23624 37624 23857 37652
rect 23624 37612 23630 37624
rect 23845 37621 23857 37624
rect 23891 37621 23903 37655
rect 27430 37652 27436 37664
rect 27391 37624 27436 37652
rect 23845 37615 23903 37621
rect 27430 37612 27436 37624
rect 27488 37612 27494 37664
rect 47762 37652 47768 37664
rect 47723 37624 47768 37652
rect 47762 37612 47768 37624
rect 47820 37612 47826 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 15930 37448 15936 37460
rect 15891 37420 15936 37448
rect 15930 37408 15936 37420
rect 15988 37408 15994 37460
rect 16482 37448 16488 37460
rect 16395 37420 16488 37448
rect 16482 37408 16488 37420
rect 16540 37448 16546 37460
rect 16540 37420 17908 37448
rect 16540 37408 16546 37420
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 2041 37207 2099 37213
rect 15562 37204 15568 37256
rect 15620 37244 15626 37256
rect 15657 37247 15715 37253
rect 15657 37244 15669 37247
rect 15620 37216 15669 37244
rect 15620 37204 15626 37216
rect 15657 37213 15669 37216
rect 15703 37213 15715 37247
rect 15657 37207 15715 37213
rect 15749 37247 15807 37253
rect 15749 37213 15761 37247
rect 15795 37244 15807 37247
rect 15930 37244 15936 37256
rect 15795 37216 15936 37244
rect 15795 37213 15807 37216
rect 15749 37207 15807 37213
rect 15930 37204 15936 37216
rect 15988 37204 15994 37256
rect 16022 37204 16028 37256
rect 16080 37244 16086 37256
rect 16500 37244 16528 37408
rect 17880 37380 17908 37420
rect 19334 37408 19340 37460
rect 19392 37448 19398 37460
rect 19610 37448 19616 37460
rect 19392 37420 19616 37448
rect 19392 37408 19398 37420
rect 19610 37408 19616 37420
rect 19668 37408 19674 37460
rect 20898 37448 20904 37460
rect 20859 37420 20904 37448
rect 20898 37408 20904 37420
rect 20956 37408 20962 37460
rect 23293 37451 23351 37457
rect 23293 37417 23305 37451
rect 23339 37417 23351 37451
rect 24946 37448 24952 37460
rect 24907 37420 24952 37448
rect 23293 37411 23351 37417
rect 19352 37380 19380 37408
rect 17880 37352 19380 37380
rect 20809 37383 20867 37389
rect 20809 37349 20821 37383
rect 20855 37380 20867 37383
rect 23308 37380 23336 37411
rect 24946 37408 24952 37420
rect 25004 37408 25010 37460
rect 26881 37451 26939 37457
rect 26881 37417 26893 37451
rect 26927 37448 26939 37451
rect 27154 37448 27160 37460
rect 26927 37420 27160 37448
rect 26927 37417 26939 37420
rect 26881 37411 26939 37417
rect 27154 37408 27160 37420
rect 27212 37408 27218 37460
rect 44266 37448 44272 37460
rect 44227 37420 44272 37448
rect 44266 37408 44272 37420
rect 44324 37408 44330 37460
rect 24857 37383 24915 37389
rect 20855 37352 22094 37380
rect 23308 37352 24808 37380
rect 20855 37349 20867 37352
rect 20809 37343 20867 37349
rect 16850 37312 16856 37324
rect 16811 37284 16856 37312
rect 16850 37272 16856 37284
rect 16908 37272 16914 37324
rect 18966 37272 18972 37324
rect 19024 37312 19030 37324
rect 20162 37312 20168 37324
rect 19024 37284 20168 37312
rect 19024 37272 19030 37284
rect 20162 37272 20168 37284
rect 20220 37272 20226 37324
rect 20993 37315 21051 37321
rect 20993 37281 21005 37315
rect 21039 37312 21051 37315
rect 21266 37312 21272 37324
rect 21039 37284 21272 37312
rect 21039 37281 21051 37284
rect 20993 37275 21051 37281
rect 21266 37272 21272 37284
rect 21324 37272 21330 37324
rect 22066 37312 22094 37352
rect 24780 37312 24808 37352
rect 24857 37349 24869 37383
rect 24903 37380 24915 37383
rect 25498 37380 25504 37392
rect 24903 37352 25504 37380
rect 24903 37349 24915 37352
rect 24857 37343 24915 37349
rect 25498 37340 25504 37352
rect 25556 37340 25562 37392
rect 26970 37340 26976 37392
rect 27028 37380 27034 37392
rect 28810 37380 28816 37392
rect 27028 37352 28816 37380
rect 27028 37340 27034 37352
rect 28810 37340 28816 37352
rect 28868 37340 28874 37392
rect 25590 37312 25596 37324
rect 22066 37284 23428 37312
rect 24780 37284 25596 37312
rect 23400 37256 23428 37284
rect 25590 37272 25596 37284
rect 25648 37272 25654 37324
rect 26513 37315 26571 37321
rect 26513 37281 26525 37315
rect 26559 37312 26571 37315
rect 26559 37284 27568 37312
rect 26559 37281 26571 37284
rect 26513 37275 26571 37281
rect 16080 37216 16528 37244
rect 16577 37247 16635 37253
rect 16080 37204 16086 37216
rect 16577 37213 16589 37247
rect 16623 37213 16635 37247
rect 19242 37244 19248 37256
rect 19203 37216 19248 37244
rect 16577 37207 16635 37213
rect 16592 37176 16620 37207
rect 19242 37204 19248 37216
rect 19300 37204 19306 37256
rect 19702 37204 19708 37256
rect 19760 37244 19766 37256
rect 20714 37244 20720 37256
rect 19760 37216 20720 37244
rect 19760 37204 19766 37216
rect 20714 37204 20720 37216
rect 20772 37204 20778 37256
rect 22833 37247 22891 37253
rect 22833 37213 22845 37247
rect 22879 37213 22891 37247
rect 23198 37244 23204 37256
rect 23159 37216 23204 37244
rect 22833 37207 22891 37213
rect 16758 37176 16764 37188
rect 16592 37148 16764 37176
rect 16758 37136 16764 37148
rect 16816 37136 16822 37188
rect 19337 37179 19395 37185
rect 19337 37176 19349 37179
rect 18078 37148 19349 37176
rect 19337 37145 19349 37148
rect 19383 37145 19395 37179
rect 19337 37139 19395 37145
rect 19794 37136 19800 37188
rect 19852 37136 19858 37188
rect 22848 37176 22876 37207
rect 23198 37204 23204 37216
rect 23256 37204 23262 37256
rect 23382 37204 23388 37256
rect 23440 37244 23446 37256
rect 26697 37247 26755 37253
rect 23440 37216 23533 37244
rect 23440 37204 23446 37216
rect 26697 37213 26709 37247
rect 26743 37244 26755 37247
rect 27338 37244 27344 37256
rect 26743 37216 27344 37244
rect 26743 37213 26755 37216
rect 26697 37207 26755 37213
rect 27338 37204 27344 37216
rect 27396 37204 27402 37256
rect 27540 37253 27568 37284
rect 27525 37247 27583 37253
rect 27525 37213 27537 37247
rect 27571 37244 27583 37247
rect 27890 37244 27896 37256
rect 27571 37216 27896 37244
rect 27571 37213 27583 37216
rect 27525 37207 27583 37213
rect 27890 37204 27896 37216
rect 27948 37244 27954 37256
rect 28350 37244 28356 37256
rect 27948 37216 28356 37244
rect 27948 37204 27954 37216
rect 28350 37204 28356 37216
rect 28408 37204 28414 37256
rect 28828 37253 28856 37340
rect 31754 37272 31760 37324
rect 31812 37312 31818 37324
rect 45373 37315 45431 37321
rect 45373 37312 45385 37315
rect 31812 37284 45385 37312
rect 31812 37272 31818 37284
rect 45373 37281 45385 37284
rect 45419 37312 45431 37315
rect 45462 37312 45468 37324
rect 45419 37284 45468 37312
rect 45419 37281 45431 37284
rect 45373 37275 45431 37281
rect 45462 37272 45468 37284
rect 45520 37272 45526 37324
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 28813 37247 28871 37253
rect 28813 37213 28825 37247
rect 28859 37213 28871 37247
rect 28813 37207 28871 37213
rect 29454 37204 29460 37256
rect 29512 37244 29518 37256
rect 44082 37244 44088 37256
rect 29512 37216 44088 37244
rect 29512 37204 29518 37216
rect 44082 37204 44088 37216
rect 44140 37204 44146 37256
rect 44266 37204 44272 37256
rect 44324 37244 44330 37256
rect 45097 37247 45155 37253
rect 45097 37244 45109 37247
rect 44324 37216 45109 37244
rect 44324 37204 44330 37216
rect 45097 37213 45109 37216
rect 45143 37213 45155 37247
rect 45097 37207 45155 37213
rect 46293 37247 46351 37253
rect 46293 37213 46305 37247
rect 46339 37213 46351 37247
rect 46293 37207 46351 37213
rect 22848 37148 24072 37176
rect 15473 37111 15531 37117
rect 15473 37077 15485 37111
rect 15519 37108 15531 37111
rect 15838 37108 15844 37120
rect 15519 37080 15844 37108
rect 15519 37077 15531 37080
rect 15473 37071 15531 37077
rect 15838 37068 15844 37080
rect 15896 37068 15902 37120
rect 18325 37111 18383 37117
rect 18325 37077 18337 37111
rect 18371 37108 18383 37111
rect 18414 37108 18420 37120
rect 18371 37080 18420 37108
rect 18371 37077 18383 37080
rect 18325 37071 18383 37077
rect 18414 37068 18420 37080
rect 18472 37068 18478 37120
rect 19812 37108 19840 37136
rect 22554 37108 22560 37120
rect 19812 37080 22560 37108
rect 22554 37068 22560 37080
rect 22612 37108 22618 37120
rect 23017 37111 23075 37117
rect 23017 37108 23029 37111
rect 22612 37080 23029 37108
rect 22612 37068 22618 37080
rect 23017 37077 23029 37080
rect 23063 37077 23075 37111
rect 24044 37108 24072 37148
rect 24118 37136 24124 37188
rect 24176 37176 24182 37188
rect 24489 37179 24547 37185
rect 24489 37176 24501 37179
rect 24176 37148 24501 37176
rect 24176 37136 24182 37148
rect 24489 37145 24501 37148
rect 24535 37145 24547 37179
rect 24489 37139 24547 37145
rect 24210 37108 24216 37120
rect 24044 37080 24216 37108
rect 23017 37071 23075 37077
rect 24210 37068 24216 37080
rect 24268 37108 24274 37120
rect 24946 37108 24952 37120
rect 24268 37080 24952 37108
rect 24268 37068 24274 37080
rect 24946 37068 24952 37080
rect 25004 37068 25010 37120
rect 27706 37108 27712 37120
rect 27667 37080 27712 37108
rect 27706 37068 27712 37080
rect 27764 37068 27770 37120
rect 28905 37111 28963 37117
rect 28905 37077 28917 37111
rect 28951 37108 28963 37111
rect 29178 37108 29184 37120
rect 28951 37080 29184 37108
rect 28951 37077 28963 37080
rect 28905 37071 28963 37077
rect 29178 37068 29184 37080
rect 29236 37068 29242 37120
rect 46308 37108 46336 37207
rect 46477 37179 46535 37185
rect 46477 37145 46489 37179
rect 46523 37176 46535 37179
rect 47670 37176 47676 37188
rect 46523 37148 47676 37176
rect 46523 37145 46535 37148
rect 46477 37139 46535 37145
rect 47670 37136 47676 37148
rect 47728 37136 47734 37188
rect 47762 37108 47768 37120
rect 46308 37080 47768 37108
rect 47762 37068 47768 37080
rect 47820 37068 47826 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 18138 36904 18144 36916
rect 18099 36876 18144 36904
rect 18138 36864 18144 36876
rect 18196 36864 18202 36916
rect 22186 36864 22192 36916
rect 22244 36904 22250 36916
rect 22649 36907 22707 36913
rect 22649 36904 22661 36907
rect 22244 36876 22661 36904
rect 22244 36864 22250 36876
rect 22649 36873 22661 36876
rect 22695 36873 22707 36907
rect 24118 36904 24124 36916
rect 24079 36876 24124 36904
rect 22649 36867 22707 36873
rect 24118 36864 24124 36876
rect 24176 36864 24182 36916
rect 27062 36904 27068 36916
rect 27023 36876 27068 36904
rect 27062 36864 27068 36876
rect 27120 36864 27126 36916
rect 27249 36907 27307 36913
rect 27249 36873 27261 36907
rect 27295 36904 27307 36907
rect 27706 36904 27712 36916
rect 27295 36876 27712 36904
rect 27295 36873 27307 36876
rect 27249 36867 27307 36873
rect 27706 36864 27712 36876
rect 27764 36864 27770 36916
rect 47670 36904 47676 36916
rect 47631 36876 47676 36904
rect 47670 36864 47676 36876
rect 47728 36864 47734 36916
rect 16761 36839 16819 36845
rect 16761 36836 16773 36839
rect 15410 36808 16773 36836
rect 16761 36805 16773 36808
rect 16807 36805 16819 36839
rect 16761 36799 16819 36805
rect 19426 36796 19432 36848
rect 19484 36836 19490 36848
rect 23198 36836 23204 36848
rect 19484 36808 23204 36836
rect 19484 36796 19490 36808
rect 23198 36796 23204 36808
rect 23256 36796 23262 36848
rect 23750 36836 23756 36848
rect 23711 36808 23756 36836
rect 23750 36796 23756 36808
rect 23808 36796 23814 36848
rect 23969 36839 24027 36845
rect 23969 36805 23981 36839
rect 24015 36836 24027 36839
rect 25038 36836 25044 36848
rect 24015 36808 25044 36836
rect 24015 36805 24027 36808
rect 23969 36799 24027 36805
rect 25038 36796 25044 36808
rect 25096 36796 25102 36848
rect 28994 36836 29000 36848
rect 25148 36808 29000 36836
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 16669 36771 16727 36777
rect 16669 36737 16681 36771
rect 16715 36768 16727 36771
rect 17773 36771 17831 36777
rect 16715 36740 17080 36768
rect 16715 36737 16727 36740
rect 16669 36731 16727 36737
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 13906 36700 13912 36712
rect 13867 36672 13912 36700
rect 13906 36660 13912 36672
rect 13964 36660 13970 36712
rect 14185 36703 14243 36709
rect 14185 36669 14197 36703
rect 14231 36700 14243 36703
rect 15654 36700 15660 36712
rect 14231 36672 15660 36700
rect 14231 36669 14243 36672
rect 14185 36663 14243 36669
rect 15654 36660 15660 36672
rect 15712 36660 15718 36712
rect 17052 36632 17080 36740
rect 17773 36737 17785 36771
rect 17819 36768 17831 36771
rect 18414 36768 18420 36780
rect 17819 36740 18420 36768
rect 17819 36737 17831 36740
rect 17773 36731 17831 36737
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 22830 36768 22836 36780
rect 22791 36740 22836 36768
rect 22830 36728 22836 36740
rect 22888 36728 22894 36780
rect 23014 36768 23020 36780
rect 22975 36740 23020 36768
rect 23014 36728 23020 36740
rect 23072 36728 23078 36780
rect 23109 36771 23167 36777
rect 23109 36737 23121 36771
rect 23155 36768 23167 36771
rect 24118 36768 24124 36780
rect 23155 36740 24124 36768
rect 23155 36737 23167 36740
rect 23109 36731 23167 36737
rect 24118 36728 24124 36740
rect 24176 36728 24182 36780
rect 24946 36768 24952 36780
rect 24907 36740 24952 36768
rect 24946 36728 24952 36740
rect 25004 36728 25010 36780
rect 17865 36703 17923 36709
rect 17865 36669 17877 36703
rect 17911 36700 17923 36703
rect 18138 36700 18144 36712
rect 17911 36672 18144 36700
rect 17911 36669 17923 36672
rect 17865 36663 17923 36669
rect 18138 36660 18144 36672
rect 18196 36660 18202 36712
rect 19334 36660 19340 36712
rect 19392 36700 19398 36712
rect 24854 36700 24860 36712
rect 19392 36672 24860 36700
rect 19392 36660 19398 36672
rect 24854 36660 24860 36672
rect 24912 36660 24918 36712
rect 18046 36632 18052 36644
rect 17052 36604 18052 36632
rect 18046 36592 18052 36604
rect 18104 36632 18110 36644
rect 19242 36632 19248 36644
rect 18104 36604 19248 36632
rect 18104 36592 18110 36604
rect 19242 36592 19248 36604
rect 19300 36592 19306 36644
rect 20714 36592 20720 36644
rect 20772 36632 20778 36644
rect 25148 36632 25176 36808
rect 28994 36796 29000 36808
rect 29052 36796 29058 36848
rect 29178 36796 29184 36848
rect 29236 36796 29242 36848
rect 44082 36796 44088 36848
rect 44140 36836 44146 36848
rect 47026 36836 47032 36848
rect 44140 36808 47032 36836
rect 44140 36796 44146 36808
rect 47026 36796 47032 36808
rect 47084 36796 47090 36848
rect 26786 36728 26792 36780
rect 26844 36768 26850 36780
rect 27190 36771 27248 36777
rect 27190 36768 27202 36771
rect 26844 36740 27202 36768
rect 26844 36728 26850 36740
rect 27190 36737 27202 36740
rect 27236 36737 27248 36771
rect 27190 36731 27248 36737
rect 27614 36728 27620 36780
rect 27672 36768 27678 36780
rect 28445 36771 28503 36777
rect 28445 36768 28457 36771
rect 27672 36740 28457 36768
rect 27672 36728 27678 36740
rect 28445 36737 28457 36740
rect 28491 36737 28503 36771
rect 28445 36731 28503 36737
rect 47210 36728 47216 36780
rect 47268 36768 47274 36780
rect 47581 36771 47639 36777
rect 47581 36768 47593 36771
rect 47268 36740 47593 36768
rect 47268 36728 47274 36740
rect 47581 36737 47593 36740
rect 47627 36737 47639 36771
rect 47581 36731 47639 36737
rect 27709 36703 27767 36709
rect 27709 36669 27721 36703
rect 27755 36700 27767 36703
rect 27890 36700 27896 36712
rect 27755 36672 27896 36700
rect 27755 36669 27767 36672
rect 27709 36663 27767 36669
rect 27890 36660 27896 36672
rect 27948 36660 27954 36712
rect 28721 36703 28779 36709
rect 28721 36669 28733 36703
rect 28767 36700 28779 36703
rect 29270 36700 29276 36712
rect 28767 36672 29276 36700
rect 28767 36669 28779 36672
rect 28721 36663 28779 36669
rect 29270 36660 29276 36672
rect 29328 36660 29334 36712
rect 47486 36660 47492 36712
rect 47544 36700 47550 36712
rect 47670 36700 47676 36712
rect 47544 36672 47676 36700
rect 47544 36660 47550 36672
rect 47670 36660 47676 36672
rect 47728 36660 47734 36712
rect 20772 36604 25176 36632
rect 20772 36592 20778 36604
rect 15657 36567 15715 36573
rect 15657 36533 15669 36567
rect 15703 36564 15715 36567
rect 15930 36564 15936 36576
rect 15703 36536 15936 36564
rect 15703 36533 15715 36536
rect 15657 36527 15715 36533
rect 15930 36524 15936 36536
rect 15988 36564 15994 36576
rect 16206 36564 16212 36576
rect 15988 36536 16212 36564
rect 15988 36524 15994 36536
rect 16206 36524 16212 36536
rect 16264 36524 16270 36576
rect 22554 36524 22560 36576
rect 22612 36564 22618 36576
rect 23290 36564 23296 36576
rect 22612 36536 23296 36564
rect 22612 36524 22618 36536
rect 23290 36524 23296 36536
rect 23348 36524 23354 36576
rect 23382 36524 23388 36576
rect 23440 36564 23446 36576
rect 23937 36567 23995 36573
rect 23937 36564 23949 36567
rect 23440 36536 23949 36564
rect 23440 36524 23446 36536
rect 23937 36533 23949 36536
rect 23983 36533 23995 36567
rect 23937 36527 23995 36533
rect 25133 36567 25191 36573
rect 25133 36533 25145 36567
rect 25179 36564 25191 36567
rect 25222 36564 25228 36576
rect 25179 36536 25228 36564
rect 25179 36533 25191 36536
rect 25133 36527 25191 36533
rect 25222 36524 25228 36536
rect 25280 36524 25286 36576
rect 25682 36524 25688 36576
rect 25740 36564 25746 36576
rect 27617 36567 27675 36573
rect 27617 36564 27629 36567
rect 25740 36536 27629 36564
rect 25740 36524 25746 36536
rect 27617 36533 27629 36536
rect 27663 36533 27675 36567
rect 27617 36527 27675 36533
rect 28810 36524 28816 36576
rect 28868 36564 28874 36576
rect 30193 36567 30251 36573
rect 30193 36564 30205 36567
rect 28868 36536 30205 36564
rect 28868 36524 28874 36536
rect 30193 36533 30205 36536
rect 30239 36533 30251 36567
rect 30193 36527 30251 36533
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 15654 36360 15660 36372
rect 15615 36332 15660 36360
rect 15654 36320 15660 36332
rect 15712 36320 15718 36372
rect 22830 36360 22836 36372
rect 22791 36332 22836 36360
rect 22830 36320 22836 36332
rect 22888 36320 22894 36372
rect 25038 36360 25044 36372
rect 24999 36332 25044 36360
rect 25038 36320 25044 36332
rect 25096 36320 25102 36372
rect 25498 36360 25504 36372
rect 25459 36332 25504 36360
rect 25498 36320 25504 36332
rect 25556 36320 25562 36372
rect 27065 36363 27123 36369
rect 27065 36329 27077 36363
rect 27111 36360 27123 36363
rect 27982 36360 27988 36372
rect 27111 36332 27988 36360
rect 27111 36329 27123 36332
rect 27065 36323 27123 36329
rect 27982 36320 27988 36332
rect 28040 36320 28046 36372
rect 15197 36295 15255 36301
rect 15197 36261 15209 36295
rect 15243 36292 15255 36295
rect 16025 36295 16083 36301
rect 16025 36292 16037 36295
rect 15243 36264 16037 36292
rect 15243 36261 15255 36264
rect 15197 36255 15255 36261
rect 16025 36261 16037 36264
rect 16071 36261 16083 36295
rect 26878 36292 26884 36304
rect 16025 36255 16083 36261
rect 23032 36264 26884 36292
rect 14918 36224 14924 36236
rect 14879 36196 14924 36224
rect 14918 36184 14924 36196
rect 14976 36184 14982 36236
rect 16206 36224 16212 36236
rect 15672 36196 16212 36224
rect 2130 36156 2136 36168
rect 2091 36128 2136 36156
rect 2130 36116 2136 36128
rect 2188 36116 2194 36168
rect 14829 36159 14887 36165
rect 14829 36125 14841 36159
rect 14875 36156 14887 36159
rect 15672 36156 15700 36196
rect 16206 36184 16212 36196
rect 16264 36184 16270 36236
rect 15838 36156 15844 36168
rect 14875 36128 15700 36156
rect 15799 36128 15844 36156
rect 14875 36125 14887 36128
rect 14829 36119 14887 36125
rect 15838 36116 15844 36128
rect 15896 36116 15902 36168
rect 16114 36156 16120 36168
rect 16075 36128 16120 36156
rect 16114 36116 16120 36128
rect 16172 36116 16178 36168
rect 20162 36116 20168 36168
rect 20220 36156 20226 36168
rect 20533 36159 20591 36165
rect 20533 36156 20545 36159
rect 20220 36128 20545 36156
rect 20220 36116 20226 36128
rect 20533 36125 20545 36128
rect 20579 36125 20591 36159
rect 20533 36119 20591 36125
rect 22005 36159 22063 36165
rect 22005 36125 22017 36159
rect 22051 36156 22063 36159
rect 22554 36156 22560 36168
rect 22051 36128 22560 36156
rect 22051 36125 22063 36128
rect 22005 36119 22063 36125
rect 22554 36116 22560 36128
rect 22612 36116 22618 36168
rect 23032 36165 23060 36264
rect 23566 36224 23572 36236
rect 23400 36196 23572 36224
rect 23017 36159 23075 36165
rect 23017 36125 23029 36159
rect 23063 36125 23075 36159
rect 23017 36119 23075 36125
rect 23201 36159 23259 36165
rect 23201 36125 23213 36159
rect 23247 36156 23259 36159
rect 23400 36156 23428 36196
rect 23566 36184 23572 36196
rect 23624 36224 23630 36236
rect 24872 36233 24900 36264
rect 26878 36252 26884 36264
rect 26936 36252 26942 36304
rect 24765 36227 24823 36233
rect 24765 36224 24777 36227
rect 23624 36196 24777 36224
rect 23624 36184 23630 36196
rect 24765 36193 24777 36196
rect 24811 36193 24823 36227
rect 24765 36187 24823 36193
rect 24857 36227 24915 36233
rect 24857 36193 24869 36227
rect 24903 36193 24915 36227
rect 25958 36224 25964 36236
rect 24857 36187 24915 36193
rect 24964 36196 25820 36224
rect 25919 36196 25964 36224
rect 23247 36128 23428 36156
rect 23477 36159 23535 36165
rect 23247 36125 23259 36128
rect 23201 36119 23259 36125
rect 23477 36125 23489 36159
rect 23523 36156 23535 36159
rect 23842 36156 23848 36168
rect 23523 36128 23848 36156
rect 23523 36125 23535 36128
rect 23477 36119 23535 36125
rect 23842 36116 23848 36128
rect 23900 36116 23906 36168
rect 24397 36159 24455 36165
rect 24397 36125 24409 36159
rect 24443 36156 24455 36159
rect 24964 36156 24992 36196
rect 24443 36128 24992 36156
rect 24443 36125 24455 36128
rect 24397 36119 24455 36125
rect 25498 36116 25504 36168
rect 25556 36156 25562 36168
rect 25682 36156 25688 36168
rect 25556 36128 25688 36156
rect 25556 36116 25562 36128
rect 25682 36116 25688 36128
rect 25740 36116 25746 36168
rect 25792 36165 25820 36196
rect 25958 36184 25964 36196
rect 26016 36184 26022 36236
rect 28810 36224 28816 36236
rect 27080 36196 28816 36224
rect 25777 36159 25835 36165
rect 25777 36125 25789 36159
rect 25823 36156 25835 36159
rect 25866 36156 25872 36168
rect 25823 36128 25872 36156
rect 25823 36125 25835 36128
rect 25777 36119 25835 36125
rect 25866 36116 25872 36128
rect 25924 36116 25930 36168
rect 26053 36159 26111 36165
rect 26053 36125 26065 36159
rect 26099 36125 26111 36159
rect 26970 36156 26976 36168
rect 26931 36128 26976 36156
rect 26053 36119 26111 36125
rect 13906 36048 13912 36100
rect 13964 36088 13970 36100
rect 16758 36088 16764 36100
rect 13964 36060 16764 36088
rect 13964 36048 13970 36060
rect 16758 36048 16764 36060
rect 16816 36048 16822 36100
rect 22186 36088 22192 36100
rect 22147 36060 22192 36088
rect 22186 36048 22192 36060
rect 22244 36048 22250 36100
rect 23106 36088 23112 36100
rect 23067 36060 23112 36088
rect 23106 36048 23112 36060
rect 23164 36048 23170 36100
rect 23290 36048 23296 36100
rect 23348 36097 23354 36100
rect 23348 36091 23377 36097
rect 23365 36057 23377 36091
rect 23348 36051 23377 36057
rect 23348 36048 23354 36051
rect 24762 36048 24768 36100
rect 24820 36088 24826 36100
rect 26068 36088 26096 36119
rect 26970 36116 26976 36128
rect 27028 36116 27034 36168
rect 27080 36165 27108 36196
rect 27065 36159 27123 36165
rect 27065 36125 27077 36159
rect 27111 36125 27123 36159
rect 27065 36119 27123 36125
rect 27706 36116 27712 36168
rect 27764 36156 27770 36168
rect 28000 36165 28028 36196
rect 28810 36184 28816 36196
rect 28868 36184 28874 36236
rect 27893 36159 27951 36165
rect 27893 36156 27905 36159
rect 27764 36128 27905 36156
rect 27764 36116 27770 36128
rect 27893 36125 27905 36128
rect 27939 36125 27951 36159
rect 27893 36119 27951 36125
rect 27985 36159 28043 36165
rect 27985 36125 27997 36159
rect 28031 36125 28043 36159
rect 27985 36119 28043 36125
rect 28169 36159 28227 36165
rect 28169 36125 28181 36159
rect 28215 36125 28227 36159
rect 28169 36119 28227 36125
rect 24820 36060 26096 36088
rect 24820 36048 24826 36060
rect 26694 36048 26700 36100
rect 26752 36088 26758 36100
rect 26789 36091 26847 36097
rect 26789 36088 26801 36091
rect 26752 36060 26801 36088
rect 26752 36048 26758 36060
rect 26789 36057 26801 36060
rect 26835 36057 26847 36091
rect 26789 36051 26847 36057
rect 26878 36048 26884 36100
rect 26936 36088 26942 36100
rect 28184 36088 28212 36119
rect 28258 36116 28264 36168
rect 28316 36156 28322 36168
rect 28316 36128 28361 36156
rect 28316 36116 28322 36128
rect 26936 36060 28212 36088
rect 26936 36048 26942 36060
rect 15194 35980 15200 36032
rect 15252 36020 15258 36032
rect 16114 36020 16120 36032
rect 15252 35992 16120 36020
rect 15252 35980 15258 35992
rect 16114 35980 16120 35992
rect 16172 35980 16178 36032
rect 20625 36023 20683 36029
rect 20625 35989 20637 36023
rect 20671 36020 20683 36023
rect 20898 36020 20904 36032
rect 20671 35992 20904 36020
rect 20671 35989 20683 35992
rect 20625 35983 20683 35989
rect 20898 35980 20904 35992
rect 20956 35980 20962 36032
rect 22370 36020 22376 36032
rect 22331 35992 22376 36020
rect 22370 35980 22376 35992
rect 22428 35980 22434 36032
rect 26234 35980 26240 36032
rect 26292 36020 26298 36032
rect 27249 36023 27307 36029
rect 27249 36020 27261 36023
rect 26292 35992 27261 36020
rect 26292 35980 26298 35992
rect 27249 35989 27261 35992
rect 27295 35989 27307 36023
rect 27249 35983 27307 35989
rect 27709 36023 27767 36029
rect 27709 35989 27721 36023
rect 27755 36020 27767 36023
rect 28534 36020 28540 36032
rect 27755 35992 28540 36020
rect 27755 35989 27767 35992
rect 27709 35983 27767 35989
rect 28534 35980 28540 35992
rect 28592 35980 28598 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 20806 35816 20812 35828
rect 19536 35788 20812 35816
rect 16758 35708 16764 35760
rect 16816 35748 16822 35760
rect 19536 35748 19564 35788
rect 20806 35776 20812 35788
rect 20864 35776 20870 35828
rect 23382 35816 23388 35828
rect 23343 35788 23388 35816
rect 23382 35776 23388 35788
rect 23440 35776 23446 35828
rect 24118 35816 24124 35828
rect 24079 35788 24124 35816
rect 24118 35776 24124 35788
rect 24176 35776 24182 35828
rect 26329 35819 26387 35825
rect 26329 35785 26341 35819
rect 26375 35816 26387 35819
rect 26878 35816 26884 35828
rect 26375 35788 26884 35816
rect 26375 35785 26387 35788
rect 26329 35779 26387 35785
rect 16816 35720 19564 35748
rect 16816 35708 16822 35720
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 17129 35683 17187 35689
rect 17129 35649 17141 35683
rect 17175 35649 17187 35683
rect 17129 35643 17187 35649
rect 17957 35683 18015 35689
rect 17957 35649 17969 35683
rect 18003 35680 18015 35683
rect 18506 35680 18512 35692
rect 18003 35652 18512 35680
rect 18003 35649 18015 35652
rect 17957 35643 18015 35649
rect 14182 35504 14188 35556
rect 14240 35544 14246 35556
rect 17144 35544 17172 35643
rect 18506 35640 18512 35652
rect 18564 35640 18570 35692
rect 19536 35689 19564 35720
rect 22186 35708 22192 35760
rect 22244 35748 22250 35760
rect 22925 35751 22983 35757
rect 22925 35748 22937 35751
rect 22244 35720 22937 35748
rect 22244 35708 22250 35720
rect 22925 35717 22937 35720
rect 22971 35748 22983 35751
rect 23566 35748 23572 35760
rect 22971 35720 23572 35748
rect 22971 35717 22983 35720
rect 22925 35711 22983 35717
rect 23566 35708 23572 35720
rect 23624 35708 23630 35760
rect 26344 35748 26372 35779
rect 26878 35776 26884 35788
rect 26936 35776 26942 35828
rect 27338 35816 27344 35828
rect 27299 35788 27344 35816
rect 27338 35776 27344 35788
rect 27396 35776 27402 35828
rect 28994 35776 29000 35828
rect 29052 35776 29058 35828
rect 29270 35816 29276 35828
rect 29231 35788 29276 35816
rect 29270 35776 29276 35788
rect 29328 35776 29334 35828
rect 29362 35776 29368 35828
rect 29420 35816 29426 35828
rect 47854 35816 47860 35828
rect 29420 35788 47860 35816
rect 29420 35776 29426 35788
rect 47854 35776 47860 35788
rect 47912 35776 47918 35828
rect 23952 35720 26372 35748
rect 29012 35748 29040 35776
rect 29638 35748 29644 35760
rect 29012 35720 29644 35748
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35649 19579 35683
rect 19521 35643 19579 35649
rect 20898 35640 20904 35692
rect 20956 35640 20962 35692
rect 22278 35680 22284 35692
rect 22239 35652 22284 35680
rect 22278 35640 22284 35652
rect 22336 35640 22342 35692
rect 22738 35640 22744 35692
rect 22796 35680 22802 35692
rect 23201 35683 23259 35689
rect 23201 35680 23213 35683
rect 22796 35652 23213 35680
rect 22796 35640 22802 35652
rect 23201 35649 23213 35652
rect 23247 35649 23259 35683
rect 23201 35643 23259 35649
rect 23474 35640 23480 35692
rect 23532 35680 23538 35692
rect 23952 35689 23980 35720
rect 29638 35708 29644 35720
rect 29696 35748 29702 35760
rect 30009 35751 30067 35757
rect 30009 35748 30021 35751
rect 29696 35720 30021 35748
rect 29696 35708 29702 35720
rect 30009 35717 30021 35720
rect 30055 35717 30067 35751
rect 30009 35711 30067 35717
rect 23845 35683 23903 35689
rect 23845 35680 23857 35683
rect 23532 35652 23857 35680
rect 23532 35640 23538 35652
rect 23845 35649 23857 35652
rect 23891 35649 23903 35683
rect 23845 35643 23903 35649
rect 23937 35683 23995 35689
rect 23937 35649 23949 35683
rect 23983 35649 23995 35683
rect 24762 35680 24768 35692
rect 23937 35643 23995 35649
rect 24044 35652 24624 35680
rect 24723 35652 24768 35680
rect 18138 35612 18144 35624
rect 18099 35584 18144 35612
rect 18138 35572 18144 35584
rect 18196 35572 18202 35624
rect 18233 35615 18291 35621
rect 18233 35581 18245 35615
rect 18279 35612 18291 35615
rect 18414 35612 18420 35624
rect 18279 35584 18420 35612
rect 18279 35581 18291 35584
rect 18233 35575 18291 35581
rect 18414 35572 18420 35584
rect 18472 35572 18478 35624
rect 19794 35612 19800 35624
rect 19755 35584 19800 35612
rect 19794 35572 19800 35584
rect 19852 35572 19858 35624
rect 20254 35572 20260 35624
rect 20312 35612 20318 35624
rect 22296 35612 22324 35640
rect 23017 35615 23075 35621
rect 23017 35612 23029 35615
rect 20312 35584 22094 35612
rect 22296 35584 23029 35612
rect 20312 35572 20318 35584
rect 18046 35544 18052 35556
rect 14240 35516 18052 35544
rect 14240 35504 14246 35516
rect 18046 35504 18052 35516
rect 18104 35504 18110 35556
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 2038 35476 2044 35488
rect 1443 35448 2044 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 2038 35436 2044 35448
rect 2096 35436 2102 35488
rect 17221 35479 17279 35485
rect 17221 35445 17233 35479
rect 17267 35476 17279 35479
rect 17494 35476 17500 35488
rect 17267 35448 17500 35476
rect 17267 35445 17279 35448
rect 17221 35439 17279 35445
rect 17494 35436 17500 35448
rect 17552 35436 17558 35488
rect 17678 35436 17684 35488
rect 17736 35476 17742 35488
rect 17773 35479 17831 35485
rect 17773 35476 17785 35479
rect 17736 35448 17785 35476
rect 17736 35436 17742 35448
rect 17773 35445 17785 35448
rect 17819 35445 17831 35479
rect 18156 35476 18184 35572
rect 22066 35544 22094 35584
rect 23017 35581 23029 35584
rect 23063 35581 23075 35615
rect 23860 35612 23888 35643
rect 24044 35612 24072 35652
rect 23860 35584 24072 35612
rect 24121 35615 24179 35621
rect 23017 35575 23075 35581
rect 24121 35581 24133 35615
rect 24167 35581 24179 35615
rect 24596 35612 24624 35652
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 25498 35680 25504 35692
rect 25459 35652 25504 35680
rect 25498 35640 25504 35652
rect 25556 35640 25562 35692
rect 26234 35680 26240 35692
rect 26195 35652 26240 35680
rect 26234 35640 26240 35652
rect 26292 35640 26298 35692
rect 26418 35680 26424 35692
rect 26379 35652 26424 35680
rect 26418 35640 26424 35652
rect 26476 35680 26482 35692
rect 26973 35683 27031 35689
rect 26973 35680 26985 35683
rect 26476 35652 26985 35680
rect 26476 35640 26482 35652
rect 26973 35649 26985 35652
rect 27019 35649 27031 35683
rect 28534 35680 28540 35692
rect 28495 35652 28540 35680
rect 26973 35643 27031 35649
rect 28534 35640 28540 35652
rect 28592 35640 28598 35692
rect 28721 35683 28779 35689
rect 28721 35649 28733 35683
rect 28767 35680 28779 35683
rect 28994 35680 29000 35692
rect 28767 35652 29000 35680
rect 28767 35649 28779 35652
rect 28721 35643 28779 35649
rect 28994 35640 29000 35652
rect 29052 35640 29058 35692
rect 29089 35683 29147 35689
rect 29089 35649 29101 35683
rect 29135 35680 29147 35683
rect 29178 35680 29184 35692
rect 29135 35652 29184 35680
rect 29135 35649 29147 35652
rect 29089 35643 29147 35649
rect 29178 35640 29184 35652
rect 29236 35640 29242 35692
rect 29825 35683 29883 35689
rect 29825 35649 29837 35683
rect 29871 35680 29883 35683
rect 29914 35680 29920 35692
rect 29871 35652 29920 35680
rect 29871 35649 29883 35652
rect 29825 35643 29883 35649
rect 29914 35640 29920 35652
rect 29972 35640 29978 35692
rect 30101 35683 30159 35689
rect 30101 35649 30113 35683
rect 30147 35649 30159 35683
rect 30101 35643 30159 35649
rect 24670 35612 24676 35624
rect 24583 35584 24676 35612
rect 24121 35575 24179 35581
rect 24136 35544 24164 35575
rect 24670 35572 24676 35584
rect 24728 35612 24734 35624
rect 27062 35612 27068 35624
rect 24728 35584 26188 35612
rect 27023 35584 27068 35612
rect 24728 35572 24734 35584
rect 25685 35547 25743 35553
rect 25685 35544 25697 35547
rect 22066 35516 25697 35544
rect 25685 35513 25697 35516
rect 25731 35544 25743 35547
rect 26050 35544 26056 35556
rect 25731 35516 26056 35544
rect 25731 35513 25743 35516
rect 25685 35507 25743 35513
rect 26050 35504 26056 35516
rect 26108 35504 26114 35556
rect 26160 35544 26188 35584
rect 27062 35572 27068 35584
rect 27120 35572 27126 35624
rect 28810 35612 28816 35624
rect 28771 35584 28816 35612
rect 28810 35572 28816 35584
rect 28868 35572 28874 35624
rect 28902 35572 28908 35624
rect 28960 35612 28966 35624
rect 28960 35584 29005 35612
rect 28960 35572 28966 35584
rect 30116 35544 30144 35643
rect 30190 35640 30196 35692
rect 30248 35680 30254 35692
rect 30248 35652 30293 35680
rect 30248 35640 30254 35652
rect 26160 35516 30144 35544
rect 21082 35476 21088 35488
rect 18156 35448 21088 35476
rect 17773 35439 17831 35445
rect 21082 35436 21088 35448
rect 21140 35436 21146 35488
rect 21266 35476 21272 35488
rect 21227 35448 21272 35476
rect 21266 35436 21272 35448
rect 21324 35436 21330 35488
rect 22373 35479 22431 35485
rect 22373 35445 22385 35479
rect 22419 35476 22431 35479
rect 22462 35476 22468 35488
rect 22419 35448 22468 35476
rect 22419 35445 22431 35448
rect 22373 35439 22431 35445
rect 22462 35436 22468 35448
rect 22520 35436 22526 35488
rect 23014 35476 23020 35488
rect 22975 35448 23020 35476
rect 23014 35436 23020 35448
rect 23072 35436 23078 35488
rect 24854 35476 24860 35488
rect 24767 35448 24860 35476
rect 24854 35436 24860 35448
rect 24912 35476 24918 35488
rect 26234 35476 26240 35488
rect 24912 35448 26240 35476
rect 24912 35436 24918 35448
rect 26234 35436 26240 35448
rect 26292 35436 26298 35488
rect 26694 35436 26700 35488
rect 26752 35476 26758 35488
rect 26973 35479 27031 35485
rect 26973 35476 26985 35479
rect 26752 35448 26985 35476
rect 26752 35436 26758 35448
rect 26973 35445 26985 35448
rect 27019 35445 27031 35479
rect 26973 35439 27031 35445
rect 30377 35479 30435 35485
rect 30377 35445 30389 35479
rect 30423 35476 30435 35479
rect 30926 35476 30932 35488
rect 30423 35448 30932 35476
rect 30423 35445 30435 35448
rect 30377 35439 30435 35445
rect 30926 35436 30932 35448
rect 30984 35436 30990 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 19794 35232 19800 35284
rect 19852 35272 19858 35284
rect 20625 35275 20683 35281
rect 20625 35272 20637 35275
rect 19852 35244 20637 35272
rect 19852 35232 19858 35244
rect 20625 35241 20637 35244
rect 20671 35241 20683 35275
rect 21082 35272 21088 35284
rect 21043 35244 21088 35272
rect 20625 35235 20683 35241
rect 21082 35232 21088 35244
rect 21140 35272 21146 35284
rect 22370 35272 22376 35284
rect 21140 35244 22232 35272
rect 22331 35244 22376 35272
rect 21140 35232 21146 35244
rect 18598 35164 18604 35216
rect 18656 35204 18662 35216
rect 22204 35204 22232 35244
rect 22370 35232 22376 35244
rect 22428 35232 22434 35284
rect 30006 35272 30012 35284
rect 26068 35244 30012 35272
rect 26068 35204 26096 35244
rect 30006 35232 30012 35244
rect 30064 35232 30070 35284
rect 18656 35176 20392 35204
rect 22204 35176 26096 35204
rect 26145 35207 26203 35213
rect 18656 35164 18662 35176
rect 16758 35136 16764 35148
rect 16719 35108 16764 35136
rect 16758 35096 16764 35108
rect 16816 35096 16822 35148
rect 19426 35028 19432 35080
rect 19484 35068 19490 35080
rect 19877 35071 19935 35077
rect 19484 35066 19840 35068
rect 19877 35066 19889 35071
rect 19484 35040 19889 35066
rect 19484 35028 19490 35040
rect 19812 35038 19889 35040
rect 19877 35037 19889 35038
rect 19923 35037 19935 35071
rect 19877 35031 19935 35037
rect 20073 35069 20131 35075
rect 20073 35035 20085 35069
rect 20119 35035 20131 35069
rect 20073 35029 20131 35035
rect 20165 35071 20223 35077
rect 20165 35037 20177 35071
rect 20211 35037 20223 35071
rect 20165 35031 20223 35037
rect 20257 35071 20315 35077
rect 20257 35037 20269 35071
rect 20303 35068 20315 35071
rect 20364 35068 20392 35176
rect 26145 35173 26157 35207
rect 26191 35204 26203 35207
rect 27525 35207 27583 35213
rect 27525 35204 27537 35207
rect 26191 35176 27537 35204
rect 26191 35173 26203 35176
rect 26145 35167 26203 35173
rect 27525 35173 27537 35176
rect 27571 35173 27583 35207
rect 27525 35167 27583 35173
rect 21174 35096 21180 35148
rect 21232 35136 21238 35148
rect 21232 35108 21277 35136
rect 21232 35096 21238 35108
rect 21450 35096 21456 35148
rect 21508 35136 21514 35148
rect 22005 35139 22063 35145
rect 22005 35136 22017 35139
rect 21508 35108 22017 35136
rect 21508 35096 21514 35108
rect 22005 35105 22017 35108
rect 22051 35105 22063 35139
rect 22462 35136 22468 35148
rect 22423 35108 22468 35136
rect 22005 35099 22063 35105
rect 22462 35096 22468 35108
rect 22520 35136 22526 35148
rect 25682 35136 25688 35148
rect 22520 35108 25688 35136
rect 22520 35096 22526 35108
rect 25682 35096 25688 35108
rect 25740 35136 25746 35148
rect 26418 35136 26424 35148
rect 25740 35108 26424 35136
rect 25740 35096 25746 35108
rect 26418 35096 26424 35108
rect 26476 35136 26482 35148
rect 26789 35139 26847 35145
rect 26789 35136 26801 35139
rect 26476 35108 26801 35136
rect 26476 35096 26482 35108
rect 26789 35105 26801 35108
rect 26835 35105 26847 35139
rect 26970 35136 26976 35148
rect 26931 35108 26976 35136
rect 26789 35099 26847 35105
rect 26970 35096 26976 35108
rect 27028 35096 27034 35148
rect 27338 35096 27344 35148
rect 27396 35136 27402 35148
rect 27396 35108 27660 35136
rect 27396 35096 27402 35108
rect 20303 35040 20392 35068
rect 20452 35071 20510 35077
rect 20303 35037 20315 35040
rect 20257 35031 20315 35037
rect 20452 35037 20464 35071
rect 20498 35068 20510 35071
rect 20714 35068 20720 35080
rect 20498 35040 20720 35068
rect 20498 35037 20510 35040
rect 20452 35031 20510 35037
rect 17034 35000 17040 35012
rect 16995 34972 17040 35000
rect 17034 34960 17040 34972
rect 17092 34960 17098 35012
rect 17494 34960 17500 35012
rect 17552 34960 17558 35012
rect 18340 34972 18644 35000
rect 15010 34892 15016 34944
rect 15068 34932 15074 34944
rect 15562 34932 15568 34944
rect 15068 34904 15568 34932
rect 15068 34892 15074 34904
rect 15562 34892 15568 34904
rect 15620 34932 15626 34944
rect 18340 34932 18368 34972
rect 18506 34932 18512 34944
rect 15620 34904 18368 34932
rect 18467 34904 18512 34932
rect 15620 34892 15626 34904
rect 18506 34892 18512 34904
rect 18564 34892 18570 34944
rect 18616 34932 18644 34972
rect 19978 34960 19984 35012
rect 20036 35000 20042 35012
rect 20088 35000 20116 35029
rect 20036 34972 20116 35000
rect 20180 35000 20208 35031
rect 20714 35028 20720 35040
rect 20772 35028 20778 35080
rect 21266 35068 21272 35080
rect 21008 35040 21272 35068
rect 21008 35000 21036 35040
rect 21266 35028 21272 35040
rect 21324 35068 21330 35080
rect 21361 35071 21419 35077
rect 21361 35068 21373 35071
rect 21324 35040 21373 35068
rect 21324 35028 21330 35040
rect 21361 35037 21373 35040
rect 21407 35068 21419 35071
rect 22189 35071 22247 35077
rect 22189 35068 22201 35071
rect 21407 35040 22201 35068
rect 21407 35037 21419 35040
rect 21361 35031 21419 35037
rect 22189 35037 22201 35040
rect 22235 35037 22247 35071
rect 22189 35031 22247 35037
rect 23750 35028 23756 35080
rect 23808 35068 23814 35080
rect 24394 35068 24400 35080
rect 23808 35040 24400 35068
rect 23808 35028 23814 35040
rect 24394 35028 24400 35040
rect 24452 35028 24458 35080
rect 25774 35068 25780 35080
rect 25735 35040 25780 35068
rect 25774 35028 25780 35040
rect 25832 35028 25838 35080
rect 25866 35028 25872 35080
rect 25924 35068 25930 35080
rect 25961 35071 26019 35077
rect 25961 35068 25973 35071
rect 25924 35040 25973 35068
rect 25924 35028 25930 35040
rect 25961 35037 25973 35040
rect 26007 35037 26019 35071
rect 25961 35031 26019 35037
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35037 26295 35071
rect 26694 35068 26700 35080
rect 26655 35040 26700 35068
rect 26237 35031 26295 35037
rect 20180 34972 21036 35000
rect 21085 35003 21143 35009
rect 20036 34960 20042 34972
rect 21085 34969 21097 35003
rect 21131 35000 21143 35003
rect 22370 35000 22376 35012
rect 21131 34972 22376 35000
rect 21131 34969 21143 34972
rect 21085 34963 21143 34969
rect 22370 34960 22376 34972
rect 22428 34960 22434 35012
rect 24118 34960 24124 35012
rect 24176 35000 24182 35012
rect 26252 35000 26280 35031
rect 26694 35028 26700 35040
rect 26752 35028 26758 35080
rect 27632 35077 27660 35108
rect 27706 35096 27712 35148
rect 27764 35136 27770 35148
rect 30377 35139 30435 35145
rect 30377 35136 30389 35139
rect 27764 35108 30389 35136
rect 27764 35096 27770 35108
rect 30377 35105 30389 35108
rect 30423 35136 30435 35139
rect 32122 35136 32128 35148
rect 30423 35108 32128 35136
rect 30423 35105 30435 35108
rect 30377 35099 30435 35105
rect 32122 35096 32128 35108
rect 32180 35096 32186 35148
rect 27433 35071 27491 35077
rect 27433 35037 27445 35071
rect 27479 35037 27491 35071
rect 27433 35031 27491 35037
rect 27617 35071 27675 35077
rect 27617 35037 27629 35071
rect 27663 35037 27675 35071
rect 48130 35068 48136 35080
rect 48091 35040 48136 35068
rect 27617 35031 27675 35037
rect 24176 34972 26280 35000
rect 26973 35003 27031 35009
rect 24176 34960 24182 34972
rect 26973 34969 26985 35003
rect 27019 35000 27031 35003
rect 27448 35000 27476 35031
rect 48130 35028 48136 35040
rect 48188 35028 48194 35080
rect 27019 34972 27476 35000
rect 30653 35003 30711 35009
rect 27019 34969 27031 34972
rect 26973 34963 27031 34969
rect 30653 34969 30665 35003
rect 30699 35000 30711 35003
rect 30742 35000 30748 35012
rect 30699 34972 30748 35000
rect 30699 34969 30711 34972
rect 30653 34963 30711 34969
rect 30742 34960 30748 34972
rect 30800 34960 30806 35012
rect 32214 35000 32220 35012
rect 31878 34972 32220 35000
rect 32214 34960 32220 34972
rect 32272 34960 32278 35012
rect 20254 34932 20260 34944
rect 18616 34904 20260 34932
rect 20254 34892 20260 34904
rect 20312 34892 20318 34944
rect 20438 34892 20444 34944
rect 20496 34932 20502 34944
rect 21174 34932 21180 34944
rect 20496 34904 21180 34932
rect 20496 34892 20502 34904
rect 21174 34892 21180 34904
rect 21232 34892 21238 34944
rect 21545 34935 21603 34941
rect 21545 34901 21557 34935
rect 21591 34932 21603 34935
rect 21726 34932 21732 34944
rect 21591 34904 21732 34932
rect 21591 34901 21603 34904
rect 21545 34895 21603 34901
rect 21726 34892 21732 34904
rect 21784 34892 21790 34944
rect 23106 34892 23112 34944
rect 23164 34932 23170 34944
rect 24581 34935 24639 34941
rect 24581 34932 24593 34935
rect 23164 34904 24593 34932
rect 23164 34892 23170 34904
rect 24581 34901 24593 34904
rect 24627 34932 24639 34935
rect 26878 34932 26884 34944
rect 24627 34904 26884 34932
rect 24627 34901 24639 34904
rect 24581 34895 24639 34901
rect 26878 34892 26884 34904
rect 26936 34892 26942 34944
rect 29914 34892 29920 34944
rect 29972 34932 29978 34944
rect 32125 34935 32183 34941
rect 32125 34932 32137 34935
rect 29972 34904 32137 34932
rect 29972 34892 29978 34904
rect 32125 34901 32137 34904
rect 32171 34901 32183 34935
rect 32125 34895 32183 34901
rect 47118 34892 47124 34944
rect 47176 34932 47182 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47176 34904 47961 34932
rect 47176 34892 47182 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 10318 34688 10324 34740
rect 10376 34728 10382 34740
rect 10376 34700 16988 34728
rect 10376 34688 10382 34700
rect 14277 34663 14335 34669
rect 14277 34629 14289 34663
rect 14323 34660 14335 34663
rect 15470 34660 15476 34672
rect 14323 34632 15476 34660
rect 14323 34629 14335 34632
rect 14277 34623 14335 34629
rect 15470 34620 15476 34632
rect 15528 34620 15534 34672
rect 16960 34660 16988 34700
rect 17034 34688 17040 34740
rect 17092 34728 17098 34740
rect 17957 34731 18015 34737
rect 17957 34728 17969 34731
rect 17092 34700 17969 34728
rect 17092 34688 17098 34700
rect 17957 34697 17969 34700
rect 18003 34697 18015 34731
rect 17957 34691 18015 34697
rect 20806 34688 20812 34740
rect 20864 34728 20870 34740
rect 22833 34731 22891 34737
rect 22833 34728 22845 34731
rect 20864 34700 22845 34728
rect 20864 34688 20870 34700
rect 22833 34697 22845 34700
rect 22879 34697 22891 34731
rect 22833 34691 22891 34697
rect 23385 34731 23443 34737
rect 23385 34697 23397 34731
rect 23431 34728 23443 34731
rect 24029 34731 24087 34737
rect 24029 34728 24041 34731
rect 23431 34700 24041 34728
rect 23431 34697 23443 34700
rect 23385 34691 23443 34697
rect 24029 34697 24041 34700
rect 24075 34697 24087 34731
rect 25866 34728 25872 34740
rect 25827 34700 25872 34728
rect 24029 34691 24087 34697
rect 18414 34660 18420 34672
rect 16960 34632 17632 34660
rect 18375 34632 18420 34660
rect 14182 34592 14188 34604
rect 14143 34564 14188 34592
rect 14182 34552 14188 34564
rect 14240 34552 14246 34604
rect 15010 34592 15016 34604
rect 14971 34564 15016 34592
rect 15010 34552 15016 34564
rect 15068 34552 15074 34604
rect 15102 34552 15108 34604
rect 15160 34592 15166 34604
rect 15381 34595 15439 34601
rect 15160 34564 15205 34592
rect 15160 34552 15166 34564
rect 15381 34561 15393 34595
rect 15427 34592 15439 34595
rect 16022 34592 16028 34604
rect 15427 34564 16028 34592
rect 15427 34561 15439 34564
rect 15381 34555 15439 34561
rect 16022 34552 16028 34564
rect 16080 34552 16086 34604
rect 17218 34592 17224 34604
rect 17179 34564 17224 34592
rect 17218 34552 17224 34564
rect 17276 34552 17282 34604
rect 17310 34552 17316 34604
rect 17368 34592 17374 34604
rect 17604 34601 17632 34632
rect 18414 34620 18420 34632
rect 18472 34620 18478 34672
rect 19426 34620 19432 34672
rect 19484 34660 19490 34672
rect 20714 34660 20720 34672
rect 19484 34632 20720 34660
rect 19484 34620 19490 34632
rect 20714 34620 20720 34632
rect 20772 34620 20778 34672
rect 20898 34620 20904 34672
rect 20956 34660 20962 34672
rect 22741 34663 22799 34669
rect 22741 34660 22753 34663
rect 20956 34632 22753 34660
rect 20956 34620 20962 34632
rect 22741 34629 22753 34632
rect 22787 34629 22799 34663
rect 24044 34660 24072 34691
rect 25866 34688 25872 34700
rect 25924 34688 25930 34740
rect 29362 34728 29368 34740
rect 26068 34700 29368 34728
rect 26068 34660 26096 34700
rect 29362 34688 29368 34700
rect 29420 34688 29426 34740
rect 30742 34728 30748 34740
rect 30703 34700 30748 34728
rect 30742 34688 30748 34700
rect 30800 34688 30806 34740
rect 32214 34728 32220 34740
rect 32175 34700 32220 34728
rect 32214 34688 32220 34700
rect 32272 34688 32278 34740
rect 26970 34660 26976 34672
rect 24044 34632 26096 34660
rect 26160 34632 26976 34660
rect 22741 34623 22799 34629
rect 17405 34595 17463 34601
rect 17405 34592 17417 34595
rect 17368 34564 17417 34592
rect 17368 34552 17374 34564
rect 17405 34561 17417 34564
rect 17451 34561 17463 34595
rect 17405 34555 17463 34561
rect 17589 34595 17647 34601
rect 17589 34561 17601 34595
rect 17635 34561 17647 34595
rect 17770 34592 17776 34604
rect 17731 34564 17776 34592
rect 17589 34555 17647 34561
rect 17770 34552 17776 34564
rect 17828 34552 17834 34604
rect 18506 34552 18512 34604
rect 18564 34592 18570 34604
rect 18601 34595 18659 34601
rect 18601 34592 18613 34595
rect 18564 34564 18613 34592
rect 18564 34552 18570 34564
rect 18601 34561 18613 34564
rect 18647 34561 18659 34595
rect 18601 34555 18659 34561
rect 19613 34595 19671 34601
rect 19613 34561 19625 34595
rect 19659 34592 19671 34595
rect 20254 34592 20260 34604
rect 19659 34564 20260 34592
rect 19659 34561 19671 34564
rect 19613 34555 19671 34561
rect 15286 34524 15292 34536
rect 15247 34496 15292 34524
rect 15286 34484 15292 34496
rect 15344 34484 15350 34536
rect 17497 34527 17555 34533
rect 17497 34493 17509 34527
rect 17543 34524 17555 34527
rect 18616 34524 18644 34555
rect 20254 34552 20260 34564
rect 20312 34552 20318 34604
rect 20349 34595 20407 34601
rect 20349 34561 20361 34595
rect 20395 34592 20407 34595
rect 20806 34592 20812 34604
rect 20395 34564 20812 34592
rect 20395 34561 20407 34564
rect 20349 34555 20407 34561
rect 20806 34552 20812 34564
rect 20864 34552 20870 34604
rect 21174 34552 21180 34604
rect 21232 34592 21238 34604
rect 21821 34595 21879 34601
rect 21821 34592 21833 34595
rect 21232 34564 21833 34592
rect 21232 34552 21238 34564
rect 21821 34561 21833 34564
rect 21867 34561 21879 34595
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21821 34555 21879 34561
rect 21928 34564 22017 34592
rect 20625 34527 20683 34533
rect 20625 34524 20637 34527
rect 17543 34496 18644 34524
rect 19352 34496 20637 34524
rect 17543 34493 17555 34496
rect 17497 34487 17555 34493
rect 17586 34416 17592 34468
rect 17644 34456 17650 34468
rect 19352 34456 19380 34496
rect 20625 34493 20637 34496
rect 20671 34524 20683 34527
rect 20990 34524 20996 34536
rect 20671 34496 20996 34524
rect 20671 34493 20683 34496
rect 20625 34487 20683 34493
rect 20990 34484 20996 34496
rect 21048 34484 21054 34536
rect 21082 34484 21088 34536
rect 21140 34524 21146 34536
rect 21928 34524 21956 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22189 34595 22247 34601
rect 22189 34561 22201 34595
rect 22235 34592 22247 34595
rect 22278 34592 22284 34604
rect 22235 34564 22284 34592
rect 22235 34561 22247 34564
rect 22189 34555 22247 34561
rect 22278 34552 22284 34564
rect 22336 34552 22342 34604
rect 26050 34592 26056 34604
rect 26011 34564 26056 34592
rect 26050 34552 26056 34564
rect 26108 34552 26114 34604
rect 26160 34601 26188 34632
rect 26970 34620 26976 34632
rect 27028 34620 27034 34672
rect 30834 34620 30840 34672
rect 30892 34660 30898 34672
rect 31113 34663 31171 34669
rect 31113 34660 31125 34663
rect 30892 34632 31125 34660
rect 30892 34620 30898 34632
rect 31113 34629 31125 34632
rect 31159 34629 31171 34663
rect 31113 34623 31171 34629
rect 26145 34595 26203 34601
rect 26145 34561 26157 34595
rect 26191 34561 26203 34595
rect 26145 34555 26203 34561
rect 26234 34552 26240 34604
rect 26292 34592 26298 34604
rect 26421 34595 26479 34601
rect 26421 34592 26433 34595
rect 26292 34564 26433 34592
rect 26292 34552 26298 34564
rect 26421 34561 26433 34564
rect 26467 34561 26479 34595
rect 29914 34592 29920 34604
rect 29827 34564 29920 34592
rect 26421 34555 26479 34561
rect 29914 34552 29920 34564
rect 29972 34592 29978 34604
rect 30098 34592 30104 34604
rect 29972 34564 30104 34592
rect 29972 34552 29978 34564
rect 30098 34552 30104 34564
rect 30156 34552 30162 34604
rect 30926 34592 30932 34604
rect 30887 34564 30932 34592
rect 30926 34552 30932 34564
rect 30984 34552 30990 34604
rect 31205 34595 31263 34601
rect 31205 34561 31217 34595
rect 31251 34561 31263 34595
rect 31205 34555 31263 34561
rect 32125 34595 32183 34601
rect 32125 34561 32137 34595
rect 32171 34592 32183 34595
rect 32858 34592 32864 34604
rect 32171 34564 32864 34592
rect 32171 34561 32183 34564
rect 32125 34555 32183 34561
rect 21140 34496 21956 34524
rect 21140 34484 21146 34496
rect 23658 34484 23664 34536
rect 23716 34524 23722 34536
rect 24121 34527 24179 34533
rect 24121 34524 24133 34527
rect 23716 34496 24133 34524
rect 23716 34484 23722 34496
rect 24121 34493 24133 34496
rect 24167 34493 24179 34527
rect 24121 34487 24179 34493
rect 24305 34527 24363 34533
rect 24305 34493 24317 34527
rect 24351 34524 24363 34527
rect 24762 34524 24768 34536
rect 24351 34496 24768 34524
rect 24351 34493 24363 34496
rect 24305 34487 24363 34493
rect 24762 34484 24768 34496
rect 24820 34524 24826 34536
rect 29822 34524 29828 34536
rect 24820 34496 24900 34524
rect 29783 34496 29828 34524
rect 24820 34484 24826 34496
rect 21450 34456 21456 34468
rect 17644 34428 19380 34456
rect 20640 34428 21456 34456
rect 17644 34416 17650 34428
rect 14550 34348 14556 34400
rect 14608 34388 14614 34400
rect 14829 34391 14887 34397
rect 14829 34388 14841 34391
rect 14608 34360 14841 34388
rect 14608 34348 14614 34360
rect 14829 34357 14841 34360
rect 14875 34357 14887 34391
rect 18782 34388 18788 34400
rect 18743 34360 18788 34388
rect 14829 34351 14887 34357
rect 18782 34348 18788 34360
rect 18840 34348 18846 34400
rect 19426 34348 19432 34400
rect 19484 34388 19490 34400
rect 19797 34391 19855 34397
rect 19797 34388 19809 34391
rect 19484 34360 19809 34388
rect 19484 34348 19490 34360
rect 19797 34357 19809 34360
rect 19843 34388 19855 34391
rect 19978 34388 19984 34400
rect 19843 34360 19984 34388
rect 19843 34357 19855 34360
rect 19797 34351 19855 34357
rect 19978 34348 19984 34360
rect 20036 34348 20042 34400
rect 20640 34397 20668 34428
rect 21450 34416 21456 34428
rect 21508 34416 21514 34468
rect 20625 34391 20683 34397
rect 20625 34357 20637 34391
rect 20671 34357 20683 34391
rect 20625 34351 20683 34357
rect 20714 34348 20720 34400
rect 20772 34388 20778 34400
rect 20901 34391 20959 34397
rect 20901 34388 20913 34391
rect 20772 34360 20913 34388
rect 20772 34348 20778 34360
rect 20901 34357 20913 34360
rect 20947 34357 20959 34391
rect 20901 34351 20959 34357
rect 20990 34348 20996 34400
rect 21048 34388 21054 34400
rect 21542 34388 21548 34400
rect 21048 34360 21548 34388
rect 21048 34348 21054 34360
rect 21542 34348 21548 34360
rect 21600 34348 21606 34400
rect 23474 34348 23480 34400
rect 23532 34388 23538 34400
rect 23661 34391 23719 34397
rect 23661 34388 23673 34391
rect 23532 34360 23673 34388
rect 23532 34348 23538 34360
rect 23661 34357 23673 34360
rect 23707 34357 23719 34391
rect 24872 34388 24900 34496
rect 29822 34484 29828 34496
rect 29880 34484 29886 34536
rect 25038 34416 25044 34468
rect 25096 34456 25102 34468
rect 29178 34456 29184 34468
rect 25096 34428 29184 34456
rect 25096 34416 25102 34428
rect 29178 34416 29184 34428
rect 29236 34416 29242 34468
rect 30285 34459 30343 34465
rect 30285 34425 30297 34459
rect 30331 34456 30343 34459
rect 31220 34456 31248 34555
rect 32858 34552 32864 34564
rect 32916 34552 32922 34604
rect 48130 34592 48136 34604
rect 48091 34564 48136 34592
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 30331 34428 31248 34456
rect 30331 34425 30343 34428
rect 30285 34419 30343 34425
rect 25130 34388 25136 34400
rect 24872 34360 25136 34388
rect 23661 34351 23719 34357
rect 25130 34348 25136 34360
rect 25188 34348 25194 34400
rect 26329 34391 26387 34397
rect 26329 34357 26341 34391
rect 26375 34388 26387 34391
rect 26418 34388 26424 34400
rect 26375 34360 26424 34388
rect 26375 34357 26387 34360
rect 26329 34351 26387 34357
rect 26418 34348 26424 34360
rect 26476 34348 26482 34400
rect 47854 34348 47860 34400
rect 47912 34388 47918 34400
rect 47949 34391 48007 34397
rect 47949 34388 47961 34391
rect 47912 34360 47961 34388
rect 47912 34348 47918 34360
rect 47949 34357 47961 34360
rect 47995 34357 48007 34391
rect 47949 34351 48007 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 15010 34144 15016 34196
rect 15068 34184 15074 34196
rect 15068 34156 16620 34184
rect 15068 34144 15074 34156
rect 13906 34008 13912 34060
rect 13964 34048 13970 34060
rect 14093 34051 14151 34057
rect 14093 34048 14105 34051
rect 13964 34020 14105 34048
rect 13964 34008 13970 34020
rect 14093 34017 14105 34020
rect 14139 34017 14151 34051
rect 14093 34011 14151 34017
rect 14918 34008 14924 34060
rect 14976 34048 14982 34060
rect 16592 34048 16620 34156
rect 17034 34144 17040 34196
rect 17092 34184 17098 34196
rect 17586 34184 17592 34196
rect 17092 34156 17592 34184
rect 17092 34144 17098 34156
rect 17586 34144 17592 34156
rect 17644 34144 17650 34196
rect 17770 34144 17776 34196
rect 17828 34184 17834 34196
rect 20625 34187 20683 34193
rect 20625 34184 20637 34187
rect 17828 34156 20637 34184
rect 17828 34144 17834 34156
rect 20625 34153 20637 34156
rect 20671 34184 20683 34187
rect 25038 34184 25044 34196
rect 20671 34156 25044 34184
rect 20671 34153 20683 34156
rect 20625 34147 20683 34153
rect 25038 34144 25044 34156
rect 25096 34144 25102 34196
rect 25332 34156 26832 34184
rect 17218 34076 17224 34128
rect 17276 34116 17282 34128
rect 17865 34119 17923 34125
rect 17865 34116 17877 34119
rect 17276 34088 17877 34116
rect 17276 34076 17282 34088
rect 17865 34085 17877 34088
rect 17911 34085 17923 34119
rect 25332 34116 25360 34156
rect 17865 34079 17923 34085
rect 17972 34088 25360 34116
rect 26804 34116 26832 34156
rect 26970 34144 26976 34196
rect 27028 34184 27034 34196
rect 27249 34187 27307 34193
rect 27249 34184 27261 34187
rect 27028 34156 27261 34184
rect 27028 34144 27034 34156
rect 27249 34153 27261 34156
rect 27295 34153 27307 34187
rect 27249 34147 27307 34153
rect 27338 34144 27344 34196
rect 27396 34184 27402 34196
rect 48041 34187 48099 34193
rect 48041 34184 48053 34187
rect 27396 34156 48053 34184
rect 27396 34144 27402 34156
rect 48041 34153 48053 34156
rect 48087 34153 48099 34187
rect 48041 34147 48099 34153
rect 28810 34116 28816 34128
rect 26804 34088 28816 34116
rect 17972 34048 18000 34088
rect 28810 34076 28816 34088
rect 28868 34076 28874 34128
rect 14976 34020 16528 34048
rect 16592 34020 18000 34048
rect 21177 34051 21235 34057
rect 14976 34008 14982 34020
rect 1578 33980 1584 33992
rect 1539 33952 1584 33980
rect 1578 33940 1584 33952
rect 1636 33940 1642 33992
rect 15470 33940 15476 33992
rect 15528 33940 15534 33992
rect 16500 33989 16528 34020
rect 17328 33989 17356 34020
rect 21177 34017 21189 34051
rect 21223 34048 21235 34051
rect 21726 34048 21732 34060
rect 21223 34020 21732 34048
rect 21223 34017 21235 34020
rect 21177 34011 21235 34017
rect 21726 34008 21732 34020
rect 21784 34008 21790 34060
rect 25406 34048 25412 34060
rect 22112 34020 25412 34048
rect 16301 33983 16359 33989
rect 16301 33949 16313 33983
rect 16347 33949 16359 33983
rect 16301 33943 16359 33949
rect 16485 33983 16543 33989
rect 16485 33949 16497 33983
rect 16531 33949 16543 33983
rect 16485 33943 16543 33949
rect 17313 33983 17371 33989
rect 17313 33949 17325 33983
rect 17359 33949 17371 33983
rect 17678 33980 17684 33992
rect 17639 33952 17684 33980
rect 17313 33943 17371 33949
rect 14366 33912 14372 33924
rect 14327 33884 14372 33912
rect 14366 33872 14372 33884
rect 14424 33872 14430 33924
rect 16316 33912 16344 33943
rect 17678 33940 17684 33952
rect 17736 33940 17742 33992
rect 20441 33983 20499 33989
rect 20441 33949 20453 33983
rect 20487 33980 20499 33983
rect 20530 33980 20536 33992
rect 20487 33952 20536 33980
rect 20487 33949 20499 33952
rect 20441 33943 20499 33949
rect 20530 33940 20536 33952
rect 20588 33940 20594 33992
rect 20714 33940 20720 33992
rect 20772 33980 20778 33992
rect 21453 33983 21511 33989
rect 21453 33980 21465 33983
rect 20772 33952 21465 33980
rect 20772 33940 20778 33952
rect 21453 33949 21465 33952
rect 21499 33949 21511 33983
rect 21453 33943 21511 33949
rect 15672 33884 16344 33912
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 1946 33844 1952 33856
rect 1443 33816 1952 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 1946 33804 1952 33816
rect 2004 33804 2010 33856
rect 13906 33804 13912 33856
rect 13964 33844 13970 33856
rect 15672 33844 15700 33884
rect 18506 33872 18512 33924
rect 18564 33912 18570 33924
rect 22112 33912 22140 34020
rect 23201 33983 23259 33989
rect 23201 33949 23213 33983
rect 23247 33980 23259 33983
rect 23474 33980 23480 33992
rect 23247 33952 23480 33980
rect 23247 33949 23259 33952
rect 23201 33943 23259 33949
rect 23474 33940 23480 33952
rect 23532 33940 23538 33992
rect 23676 33989 23704 34020
rect 25406 34008 25412 34020
rect 25464 34008 25470 34060
rect 27614 34048 27620 34060
rect 25516 34020 27620 34048
rect 23661 33983 23719 33989
rect 23661 33949 23673 33983
rect 23707 33949 23719 33983
rect 24394 33980 24400 33992
rect 24355 33952 24400 33980
rect 23661 33943 23719 33949
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 25516 33989 25544 34020
rect 27614 34008 27620 34020
rect 27672 34008 27678 34060
rect 25501 33983 25559 33989
rect 25501 33949 25513 33983
rect 25547 33949 25559 33983
rect 25501 33943 25559 33949
rect 18564 33884 22140 33912
rect 18564 33872 18570 33884
rect 22186 33872 22192 33924
rect 22244 33912 22250 33924
rect 25516 33912 25544 33943
rect 27706 33940 27712 33992
rect 27764 33980 27770 33992
rect 27801 33983 27859 33989
rect 27801 33980 27813 33983
rect 27764 33952 27813 33980
rect 27764 33940 27770 33952
rect 27801 33949 27813 33952
rect 27847 33949 27859 33983
rect 30377 33983 30435 33989
rect 27801 33943 27859 33949
rect 30024 33952 30328 33980
rect 25774 33912 25780 33924
rect 22244 33884 25544 33912
rect 25735 33884 25780 33912
rect 22244 33872 22250 33884
rect 25774 33872 25780 33884
rect 25832 33872 25838 33924
rect 26326 33872 26332 33924
rect 26384 33872 26390 33924
rect 30024 33912 30052 33952
rect 27816 33884 30052 33912
rect 15838 33844 15844 33856
rect 13964 33816 15700 33844
rect 15799 33816 15844 33844
rect 13964 33804 13970 33816
rect 15838 33804 15844 33816
rect 15896 33804 15902 33856
rect 16390 33844 16396 33856
rect 16351 33816 16396 33844
rect 16390 33804 16396 33816
rect 16448 33804 16454 33856
rect 22462 33804 22468 33856
rect 22520 33844 22526 33856
rect 23017 33847 23075 33853
rect 23017 33844 23029 33847
rect 22520 33816 23029 33844
rect 22520 33804 22526 33816
rect 23017 33813 23029 33816
rect 23063 33813 23075 33847
rect 23750 33844 23756 33856
rect 23711 33816 23756 33844
rect 23017 33807 23075 33813
rect 23750 33804 23756 33816
rect 23808 33804 23814 33856
rect 24578 33844 24584 33856
rect 24539 33816 24584 33844
rect 24578 33804 24584 33816
rect 24636 33844 24642 33856
rect 27816 33844 27844 33884
rect 30098 33872 30104 33924
rect 30156 33912 30162 33924
rect 30193 33915 30251 33921
rect 30193 33912 30205 33915
rect 30156 33884 30205 33912
rect 30156 33872 30162 33884
rect 30193 33881 30205 33884
rect 30239 33881 30251 33915
rect 30300 33912 30328 33952
rect 30377 33949 30389 33983
rect 30423 33980 30435 33983
rect 31021 33983 31079 33989
rect 31021 33980 31033 33983
rect 30423 33952 31033 33980
rect 30423 33949 30435 33952
rect 30377 33943 30435 33949
rect 31021 33949 31033 33952
rect 31067 33980 31079 33983
rect 31754 33980 31760 33992
rect 31067 33952 31760 33980
rect 31067 33949 31079 33952
rect 31021 33943 31079 33949
rect 31754 33940 31760 33952
rect 31812 33940 31818 33992
rect 30834 33912 30840 33924
rect 30300 33884 30840 33912
rect 30193 33875 30251 33881
rect 30834 33872 30840 33884
rect 30892 33872 30898 33924
rect 47946 33912 47952 33924
rect 47907 33884 47952 33912
rect 47946 33872 47952 33884
rect 48004 33872 48010 33924
rect 27982 33844 27988 33856
rect 24636 33816 27844 33844
rect 27943 33816 27988 33844
rect 24636 33804 24642 33816
rect 27982 33804 27988 33816
rect 28040 33804 28046 33856
rect 29362 33804 29368 33856
rect 29420 33844 29426 33856
rect 30561 33847 30619 33853
rect 30561 33844 30573 33847
rect 29420 33816 30573 33844
rect 29420 33804 29426 33816
rect 30561 33813 30573 33816
rect 30607 33813 30619 33847
rect 31110 33844 31116 33856
rect 31071 33816 31116 33844
rect 30561 33807 30619 33813
rect 31110 33804 31116 33816
rect 31168 33804 31174 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 13906 33640 13912 33652
rect 13867 33612 13912 33640
rect 13906 33600 13912 33612
rect 13964 33600 13970 33652
rect 14366 33640 14372 33652
rect 14327 33612 14372 33640
rect 14366 33600 14372 33612
rect 14424 33600 14430 33652
rect 15838 33600 15844 33652
rect 15896 33640 15902 33652
rect 18325 33643 18383 33649
rect 15896 33612 18184 33640
rect 15896 33600 15902 33612
rect 16390 33572 16396 33584
rect 14752 33544 16396 33572
rect 13633 33507 13691 33513
rect 13633 33473 13645 33507
rect 13679 33504 13691 33507
rect 14366 33504 14372 33516
rect 13679 33476 14372 33504
rect 13679 33473 13691 33476
rect 13633 33467 13691 33473
rect 14366 33464 14372 33476
rect 14424 33464 14430 33516
rect 14550 33504 14556 33516
rect 14511 33476 14556 33504
rect 14550 33464 14556 33476
rect 14608 33464 14614 33516
rect 14752 33513 14780 33544
rect 16390 33532 16396 33544
rect 16448 33532 16454 33584
rect 14737 33507 14795 33513
rect 14737 33473 14749 33507
rect 14783 33473 14795 33507
rect 14737 33467 14795 33473
rect 14829 33507 14887 33513
rect 14829 33473 14841 33507
rect 14875 33504 14887 33507
rect 15194 33504 15200 33516
rect 14875 33476 15200 33504
rect 14875 33473 14887 33476
rect 14829 33467 14887 33473
rect 15194 33464 15200 33476
rect 15252 33464 15258 33516
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33504 15899 33507
rect 16850 33504 16856 33516
rect 15887 33476 16436 33504
rect 16811 33476 16856 33504
rect 15887 33473 15899 33476
rect 15841 33467 15899 33473
rect 16408 33448 16436 33476
rect 16850 33464 16856 33476
rect 16908 33464 16914 33516
rect 17862 33504 17868 33516
rect 16960 33476 17264 33504
rect 17823 33476 17868 33504
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 1854 33436 1860 33448
rect 1719 33408 1860 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 1854 33396 1860 33408
rect 1912 33396 1918 33448
rect 13906 33436 13912 33448
rect 13867 33408 13912 33436
rect 13906 33396 13912 33408
rect 13964 33396 13970 33448
rect 14918 33396 14924 33448
rect 14976 33436 14982 33448
rect 16025 33439 16083 33445
rect 16025 33436 16037 33439
rect 14976 33408 16037 33436
rect 14976 33396 14982 33408
rect 16025 33405 16037 33408
rect 16071 33405 16083 33439
rect 16025 33399 16083 33405
rect 16117 33439 16175 33445
rect 16117 33405 16129 33439
rect 16163 33436 16175 33439
rect 16206 33436 16212 33448
rect 16163 33408 16212 33436
rect 16163 33405 16175 33408
rect 16117 33399 16175 33405
rect 16206 33396 16212 33408
rect 16264 33396 16270 33448
rect 16390 33396 16396 33448
rect 16448 33396 16454 33448
rect 16482 33396 16488 33448
rect 16540 33436 16546 33448
rect 16960 33436 16988 33476
rect 16540 33408 16988 33436
rect 17129 33439 17187 33445
rect 16540 33396 16546 33408
rect 17129 33405 17141 33439
rect 17175 33405 17187 33439
rect 17236 33436 17264 33476
rect 17862 33464 17868 33476
rect 17920 33464 17926 33516
rect 18156 33513 18184 33612
rect 18325 33609 18337 33643
rect 18371 33640 18383 33643
rect 20438 33640 20444 33652
rect 18371 33612 20444 33640
rect 18371 33609 18383 33612
rect 18325 33603 18383 33609
rect 20438 33600 20444 33612
rect 20496 33600 20502 33652
rect 20530 33600 20536 33652
rect 20588 33640 20594 33652
rect 24302 33640 24308 33652
rect 20588 33612 24308 33640
rect 20588 33600 20594 33612
rect 24302 33600 24308 33612
rect 24360 33600 24366 33652
rect 25406 33600 25412 33652
rect 25464 33640 25470 33652
rect 26142 33640 26148 33652
rect 25464 33612 26148 33640
rect 25464 33600 25470 33612
rect 26142 33600 26148 33612
rect 26200 33600 26206 33652
rect 26326 33640 26332 33652
rect 26287 33612 26332 33640
rect 26326 33600 26332 33612
rect 26384 33600 26390 33652
rect 27614 33640 27620 33652
rect 27575 33612 27620 33640
rect 27614 33600 27620 33612
rect 27672 33600 27678 33652
rect 28810 33640 28816 33652
rect 28771 33612 28816 33640
rect 28810 33600 28816 33612
rect 28868 33600 28874 33652
rect 21085 33575 21143 33581
rect 21085 33541 21097 33575
rect 21131 33572 21143 33575
rect 22002 33572 22008 33584
rect 21131 33544 22008 33572
rect 21131 33541 21143 33544
rect 21085 33535 21143 33541
rect 22002 33532 22008 33544
rect 22060 33532 22066 33584
rect 22462 33572 22468 33584
rect 22423 33544 22468 33572
rect 22462 33532 22468 33544
rect 22520 33532 22526 33584
rect 23750 33572 23756 33584
rect 23690 33544 23756 33572
rect 23750 33532 23756 33544
rect 23808 33532 23814 33584
rect 24949 33575 25007 33581
rect 24949 33541 24961 33575
rect 24995 33572 25007 33575
rect 27338 33572 27344 33584
rect 24995 33544 27344 33572
rect 24995 33541 25007 33544
rect 24949 33535 25007 33541
rect 18141 33507 18199 33513
rect 18141 33473 18153 33507
rect 18187 33473 18199 33507
rect 22186 33504 22192 33516
rect 22147 33476 22192 33504
rect 18141 33467 18199 33473
rect 22186 33464 22192 33476
rect 22244 33464 22250 33516
rect 25608 33513 25636 33544
rect 27338 33532 27344 33544
rect 27396 33532 27402 33584
rect 29822 33572 29828 33584
rect 29564 33544 29828 33572
rect 25593 33507 25651 33513
rect 25593 33473 25605 33507
rect 25639 33473 25651 33507
rect 25593 33467 25651 33473
rect 26142 33464 26148 33516
rect 26200 33504 26206 33516
rect 26237 33507 26295 33513
rect 26237 33504 26249 33507
rect 26200 33476 26249 33504
rect 26200 33464 26206 33476
rect 26237 33473 26249 33476
rect 26283 33504 26295 33507
rect 26970 33504 26976 33516
rect 26283 33476 26976 33504
rect 26283 33473 26295 33476
rect 26237 33467 26295 33473
rect 26970 33464 26976 33476
rect 27028 33464 27034 33516
rect 27525 33507 27583 33513
rect 27525 33473 27537 33507
rect 27571 33504 27583 33507
rect 27798 33504 27804 33516
rect 27571 33476 27804 33504
rect 27571 33473 27583 33476
rect 27525 33467 27583 33473
rect 27798 33464 27804 33476
rect 27856 33464 27862 33516
rect 28169 33507 28227 33513
rect 28169 33473 28181 33507
rect 28215 33473 28227 33507
rect 28169 33467 28227 33473
rect 28316 33507 28374 33513
rect 28316 33473 28328 33507
rect 28362 33504 28374 33507
rect 29362 33504 29368 33516
rect 28362 33476 29368 33504
rect 28362 33473 28374 33476
rect 28316 33467 28374 33473
rect 18049 33439 18107 33445
rect 17236 33408 17908 33436
rect 17129 33399 17187 33405
rect 15657 33371 15715 33377
rect 15657 33337 15669 33371
rect 15703 33368 15715 33371
rect 17144 33368 17172 33399
rect 15703 33340 17172 33368
rect 15703 33337 15715 33340
rect 15657 33331 15715 33337
rect 13725 33303 13783 33309
rect 13725 33269 13737 33303
rect 13771 33300 13783 33303
rect 15010 33300 15016 33312
rect 13771 33272 15016 33300
rect 13771 33269 13783 33272
rect 13725 33263 13783 33269
rect 15010 33260 15016 33272
rect 15068 33260 15074 33312
rect 17034 33300 17040 33312
rect 16995 33272 17040 33300
rect 17034 33260 17040 33272
rect 17092 33260 17098 33312
rect 17126 33260 17132 33312
rect 17184 33300 17190 33312
rect 17880 33309 17908 33408
rect 18049 33405 18061 33439
rect 18095 33436 18107 33439
rect 18782 33436 18788 33448
rect 18095 33408 18788 33436
rect 18095 33405 18107 33408
rect 18049 33399 18107 33405
rect 18782 33396 18788 33408
rect 18840 33436 18846 33448
rect 28184 33436 28212 33467
rect 29362 33464 29368 33476
rect 29420 33464 29426 33516
rect 18840 33408 28212 33436
rect 28537 33439 28595 33445
rect 18840 33396 18846 33408
rect 28537 33405 28549 33439
rect 28583 33436 28595 33439
rect 29564 33436 29592 33544
rect 29822 33532 29828 33544
rect 29880 33532 29886 33584
rect 30006 33532 30012 33584
rect 30064 33572 30070 33584
rect 30101 33575 30159 33581
rect 30101 33572 30113 33575
rect 30064 33544 30113 33572
rect 30064 33532 30070 33544
rect 30101 33541 30113 33544
rect 30147 33541 30159 33575
rect 30101 33535 30159 33541
rect 29641 33507 29699 33513
rect 29641 33473 29653 33507
rect 29687 33504 29699 33507
rect 29730 33504 29736 33516
rect 29687 33476 29736 33504
rect 29687 33473 29699 33476
rect 29641 33467 29699 33473
rect 29730 33464 29736 33476
rect 29788 33464 29794 33516
rect 28583 33408 29592 33436
rect 28583 33405 28595 33408
rect 28537 33399 28595 33405
rect 25314 33328 25320 33380
rect 25372 33368 25378 33380
rect 25590 33368 25596 33380
rect 25372 33340 25596 33368
rect 25372 33328 25378 33340
rect 25590 33328 25596 33340
rect 25648 33368 25654 33380
rect 25685 33371 25743 33377
rect 25685 33368 25697 33371
rect 25648 33340 25697 33368
rect 25648 33328 25654 33340
rect 25685 33337 25697 33340
rect 25731 33337 25743 33371
rect 25685 33331 25743 33337
rect 28445 33371 28503 33377
rect 28445 33337 28457 33371
rect 28491 33368 28503 33371
rect 29457 33371 29515 33377
rect 29457 33368 29469 33371
rect 28491 33340 29469 33368
rect 28491 33337 28503 33340
rect 28445 33331 28503 33337
rect 29457 33337 29469 33340
rect 29503 33368 29515 33371
rect 29546 33368 29552 33380
rect 29503 33340 29552 33368
rect 29503 33337 29515 33340
rect 29457 33331 29515 33337
rect 29546 33328 29552 33340
rect 29604 33328 29610 33380
rect 30116 33368 30144 33535
rect 33134 33532 33140 33584
rect 33192 33532 33198 33584
rect 30561 33507 30619 33513
rect 30561 33473 30573 33507
rect 30607 33504 30619 33507
rect 31110 33504 31116 33516
rect 30607 33476 31116 33504
rect 30607 33473 30619 33476
rect 30561 33467 30619 33473
rect 31110 33464 31116 33476
rect 31168 33464 31174 33516
rect 32122 33504 32128 33516
rect 32083 33476 32128 33504
rect 32122 33464 32128 33476
rect 32180 33464 32186 33516
rect 47029 33507 47087 33513
rect 47029 33473 47041 33507
rect 47075 33473 47087 33507
rect 47029 33467 47087 33473
rect 47581 33507 47639 33513
rect 47581 33473 47593 33507
rect 47627 33504 47639 33507
rect 48222 33504 48228 33516
rect 47627 33476 48228 33504
rect 47627 33473 47639 33476
rect 47581 33467 47639 33473
rect 30834 33436 30840 33448
rect 30795 33408 30840 33436
rect 30834 33396 30840 33408
rect 30892 33396 30898 33448
rect 30929 33439 30987 33445
rect 30929 33405 30941 33439
rect 30975 33405 30987 33439
rect 32398 33436 32404 33448
rect 32359 33408 32404 33436
rect 30929 33399 30987 33405
rect 30944 33368 30972 33399
rect 32398 33396 32404 33408
rect 32456 33396 32462 33448
rect 47044 33436 47072 33467
rect 48222 33464 48228 33476
rect 48280 33464 48286 33516
rect 48041 33439 48099 33445
rect 48041 33436 48053 33439
rect 47044 33408 48053 33436
rect 48041 33405 48053 33408
rect 48087 33405 48099 33439
rect 48041 33399 48099 33405
rect 30116 33340 30972 33368
rect 17405 33303 17463 33309
rect 17405 33300 17417 33303
rect 17184 33272 17417 33300
rect 17184 33260 17190 33272
rect 17405 33269 17417 33272
rect 17451 33269 17463 33303
rect 17405 33263 17463 33269
rect 17865 33303 17923 33309
rect 17865 33269 17877 33303
rect 17911 33269 17923 33303
rect 17865 33263 17923 33269
rect 20898 33260 20904 33312
rect 20956 33300 20962 33312
rect 21177 33303 21235 33309
rect 21177 33300 21189 33303
rect 20956 33272 21189 33300
rect 20956 33260 20962 33272
rect 21177 33269 21189 33272
rect 21223 33269 21235 33303
rect 23934 33300 23940 33312
rect 23895 33272 23940 33300
rect 21177 33263 21235 33269
rect 23934 33260 23940 33272
rect 23992 33260 23998 33312
rect 25041 33303 25099 33309
rect 25041 33269 25053 33303
rect 25087 33300 25099 33303
rect 25406 33300 25412 33312
rect 25087 33272 25412 33300
rect 25087 33269 25099 33272
rect 25041 33263 25099 33269
rect 25406 33260 25412 33272
rect 25464 33260 25470 33312
rect 29178 33260 29184 33312
rect 29236 33300 29242 33312
rect 30653 33303 30711 33309
rect 30653 33300 30665 33303
rect 29236 33272 30665 33300
rect 29236 33260 29242 33272
rect 30653 33269 30665 33272
rect 30699 33269 30711 33303
rect 30653 33263 30711 33269
rect 31021 33303 31079 33309
rect 31021 33269 31033 33303
rect 31067 33300 31079 33303
rect 31478 33300 31484 33312
rect 31067 33272 31484 33300
rect 31067 33269 31079 33272
rect 31021 33263 31079 33269
rect 31478 33260 31484 33272
rect 31536 33260 31542 33312
rect 31754 33260 31760 33312
rect 31812 33300 31818 33312
rect 33873 33303 33931 33309
rect 33873 33300 33885 33303
rect 31812 33272 33885 33300
rect 31812 33260 31818 33272
rect 33873 33269 33885 33272
rect 33919 33269 33931 33303
rect 33873 33263 33931 33269
rect 46845 33303 46903 33309
rect 46845 33269 46857 33303
rect 46891 33300 46903 33303
rect 47210 33300 47216 33312
rect 46891 33272 47216 33300
rect 46891 33269 46903 33272
rect 46845 33263 46903 33269
rect 47210 33260 47216 33272
rect 47268 33260 47274 33312
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1946 33096 1952 33108
rect 1907 33068 1952 33096
rect 1946 33056 1952 33068
rect 2004 33056 2010 33108
rect 14366 33056 14372 33108
rect 14424 33096 14430 33108
rect 14461 33099 14519 33105
rect 14461 33096 14473 33099
rect 14424 33068 14473 33096
rect 14424 33056 14430 33068
rect 14461 33065 14473 33068
rect 14507 33096 14519 33099
rect 15289 33099 15347 33105
rect 15289 33096 15301 33099
rect 14507 33068 15301 33096
rect 14507 33065 14519 33068
rect 14461 33059 14519 33065
rect 15289 33065 15301 33068
rect 15335 33065 15347 33099
rect 15289 33059 15347 33065
rect 16485 33099 16543 33105
rect 16485 33065 16497 33099
rect 16531 33065 16543 33099
rect 16485 33059 16543 33065
rect 16669 33099 16727 33105
rect 16669 33065 16681 33099
rect 16715 33096 16727 33099
rect 17862 33096 17868 33108
rect 16715 33068 17868 33096
rect 16715 33065 16727 33068
rect 16669 33059 16727 33065
rect 14829 33031 14887 33037
rect 14829 32997 14841 33031
rect 14875 33028 14887 33031
rect 14918 33028 14924 33040
rect 14875 33000 14924 33028
rect 14875 32997 14887 33000
rect 14829 32991 14887 32997
rect 14918 32988 14924 33000
rect 14976 32988 14982 33040
rect 16500 33028 16528 33059
rect 17862 33056 17868 33068
rect 17920 33056 17926 33108
rect 20990 33096 20996 33108
rect 20088 33068 20996 33096
rect 17218 33028 17224 33040
rect 16500 33000 17224 33028
rect 17218 32988 17224 33000
rect 17276 32988 17282 33040
rect 17310 32988 17316 33040
rect 17368 33028 17374 33040
rect 20088 33028 20116 33068
rect 20990 33056 20996 33068
rect 21048 33056 21054 33108
rect 22094 33056 22100 33108
rect 22152 33096 22158 33108
rect 26053 33099 26111 33105
rect 26053 33096 26065 33099
rect 22152 33068 26065 33096
rect 22152 33056 22158 33068
rect 26053 33065 26065 33068
rect 26099 33065 26111 33099
rect 26053 33059 26111 33065
rect 23658 33028 23664 33040
rect 17368 33000 20116 33028
rect 23619 33000 23664 33028
rect 17368 32988 17374 33000
rect 23658 32988 23664 33000
rect 23716 32988 23722 33040
rect 2317 32963 2375 32969
rect 2317 32929 2329 32963
rect 2363 32960 2375 32963
rect 2363 32932 3004 32960
rect 2363 32929 2375 32932
rect 2317 32923 2375 32929
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32892 1915 32895
rect 1946 32892 1952 32904
rect 1903 32864 1952 32892
rect 1903 32861 1915 32864
rect 1857 32855 1915 32861
rect 1946 32852 1952 32864
rect 2004 32852 2010 32904
rect 2976 32901 3004 32932
rect 13906 32920 13912 32972
rect 13964 32960 13970 32972
rect 14553 32963 14611 32969
rect 14553 32960 14565 32963
rect 13964 32932 14565 32960
rect 13964 32920 13970 32932
rect 14553 32929 14565 32932
rect 14599 32960 14611 32963
rect 15102 32960 15108 32972
rect 14599 32932 15108 32960
rect 14599 32929 14611 32932
rect 14553 32923 14611 32929
rect 15102 32920 15108 32932
rect 15160 32960 15166 32972
rect 23385 32963 23443 32969
rect 15160 32932 15608 32960
rect 15160 32920 15166 32932
rect 2961 32895 3019 32901
rect 2961 32861 2973 32895
rect 3007 32861 3019 32895
rect 14458 32892 14464 32904
rect 14371 32864 14464 32892
rect 2961 32855 3019 32861
rect 14458 32852 14464 32864
rect 14516 32892 14522 32904
rect 15010 32892 15016 32904
rect 14516 32864 15016 32892
rect 14516 32852 14522 32864
rect 15010 32852 15016 32864
rect 15068 32892 15074 32904
rect 15289 32895 15347 32901
rect 15289 32892 15301 32895
rect 15068 32864 15301 32892
rect 15068 32852 15074 32864
rect 15289 32861 15301 32864
rect 15335 32861 15347 32895
rect 15470 32892 15476 32904
rect 15431 32864 15476 32892
rect 15289 32855 15347 32861
rect 15470 32852 15476 32864
rect 15528 32852 15534 32904
rect 15580 32901 15608 32932
rect 16500 32932 23336 32960
rect 15565 32895 15623 32901
rect 15565 32861 15577 32895
rect 15611 32892 15623 32895
rect 15838 32892 15844 32904
rect 15611 32864 15844 32892
rect 15611 32861 15623 32864
rect 15565 32855 15623 32861
rect 15838 32852 15844 32864
rect 15896 32852 15902 32904
rect 16390 32892 16396 32904
rect 16351 32864 16396 32892
rect 16390 32852 16396 32864
rect 16448 32852 16454 32904
rect 16500 32901 16528 32932
rect 16485 32895 16543 32901
rect 16485 32861 16497 32895
rect 16531 32861 16543 32895
rect 17126 32892 17132 32904
rect 17087 32864 17132 32892
rect 16485 32855 16543 32861
rect 17126 32852 17132 32864
rect 17184 32852 17190 32904
rect 17310 32892 17316 32904
rect 17271 32864 17316 32892
rect 17310 32852 17316 32864
rect 17368 32852 17374 32904
rect 17405 32895 17463 32901
rect 17405 32861 17417 32895
rect 17451 32861 17463 32895
rect 17405 32855 17463 32861
rect 16206 32824 16212 32836
rect 16167 32796 16212 32824
rect 16206 32784 16212 32796
rect 16264 32784 16270 32836
rect 2222 32716 2228 32768
rect 2280 32756 2286 32768
rect 2777 32759 2835 32765
rect 2777 32756 2789 32759
rect 2280 32728 2789 32756
rect 2280 32716 2286 32728
rect 2777 32725 2789 32728
rect 2823 32725 2835 32759
rect 2777 32719 2835 32725
rect 15749 32759 15807 32765
rect 15749 32725 15761 32759
rect 15795 32756 15807 32759
rect 16850 32756 16856 32768
rect 15795 32728 16856 32756
rect 15795 32725 15807 32728
rect 15749 32719 15807 32725
rect 16850 32716 16856 32728
rect 16908 32716 16914 32768
rect 17310 32716 17316 32768
rect 17368 32756 17374 32768
rect 17420 32756 17448 32855
rect 17494 32852 17500 32904
rect 17552 32892 17558 32904
rect 17681 32895 17739 32901
rect 17552 32864 17597 32892
rect 17552 32852 17558 32864
rect 17681 32861 17693 32895
rect 17727 32892 17739 32895
rect 17770 32892 17776 32904
rect 17727 32864 17776 32892
rect 17727 32861 17739 32864
rect 17681 32855 17739 32861
rect 17770 32852 17776 32864
rect 17828 32852 17834 32904
rect 18506 32892 18512 32904
rect 18467 32864 18512 32892
rect 18506 32852 18512 32864
rect 18564 32852 18570 32904
rect 19978 32892 19984 32904
rect 19939 32864 19984 32892
rect 19978 32852 19984 32864
rect 20036 32852 20042 32904
rect 22186 32892 22192 32904
rect 22147 32864 22192 32892
rect 22186 32852 22192 32864
rect 22244 32852 22250 32904
rect 23308 32901 23336 32932
rect 23385 32929 23397 32963
rect 23431 32960 23443 32963
rect 23474 32960 23480 32972
rect 23431 32932 23480 32960
rect 23431 32929 23443 32932
rect 23385 32923 23443 32929
rect 23474 32920 23480 32932
rect 23532 32920 23538 32972
rect 23293 32895 23351 32901
rect 23293 32861 23305 32895
rect 23339 32892 23351 32895
rect 23934 32892 23940 32904
rect 23339 32864 23940 32892
rect 23339 32861 23351 32864
rect 23293 32855 23351 32861
rect 23934 32852 23940 32864
rect 23992 32852 23998 32904
rect 26068 32892 26096 33059
rect 29270 33056 29276 33108
rect 29328 33096 29334 33108
rect 32217 33099 32275 33105
rect 29328 33068 32076 33096
rect 29328 33056 29334 33068
rect 26418 32988 26424 33040
rect 26476 33028 26482 33040
rect 31938 33028 31944 33040
rect 26476 33000 31944 33028
rect 26476 32988 26482 33000
rect 31938 32988 31944 33000
rect 31996 32988 32002 33040
rect 29822 32920 29828 32972
rect 29880 32960 29886 32972
rect 29917 32963 29975 32969
rect 29917 32960 29929 32963
rect 29880 32932 29929 32960
rect 29880 32920 29886 32932
rect 29917 32929 29929 32932
rect 29963 32929 29975 32963
rect 29917 32923 29975 32929
rect 31754 32920 31760 32972
rect 31812 32960 31818 32972
rect 31812 32932 31857 32960
rect 31812 32920 31818 32932
rect 32048 32904 32076 33068
rect 32217 33065 32229 33099
rect 32263 33096 32275 33099
rect 32398 33096 32404 33108
rect 32263 33068 32404 33096
rect 32263 33065 32275 33068
rect 32217 33059 32275 33065
rect 32398 33056 32404 33068
rect 32456 33056 32462 33108
rect 32953 33099 33011 33105
rect 32953 33065 32965 33099
rect 32999 33096 33011 33099
rect 33134 33096 33140 33108
rect 32999 33068 33140 33096
rect 32999 33065 33011 33068
rect 32953 33059 33011 33065
rect 33134 33056 33140 33068
rect 33192 33056 33198 33108
rect 47118 32960 47124 32972
rect 47079 32932 47124 32960
rect 47118 32920 47124 32932
rect 47176 32920 47182 32972
rect 47670 32960 47676 32972
rect 47631 32932 47676 32960
rect 47670 32920 47676 32932
rect 47728 32920 47734 32972
rect 27065 32895 27123 32901
rect 27065 32892 27077 32895
rect 26068 32864 27077 32892
rect 27065 32861 27077 32864
rect 27111 32861 27123 32895
rect 27065 32855 27123 32861
rect 29641 32895 29699 32901
rect 29641 32861 29653 32895
rect 29687 32892 29699 32895
rect 29730 32892 29736 32904
rect 29687 32864 29736 32892
rect 29687 32861 29699 32864
rect 29641 32855 29699 32861
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 31478 32892 31484 32904
rect 31439 32864 31484 32892
rect 31478 32852 31484 32864
rect 31536 32852 31542 32904
rect 31665 32895 31723 32901
rect 31665 32861 31677 32895
rect 31711 32861 31723 32895
rect 31665 32855 31723 32861
rect 20254 32824 20260 32836
rect 20215 32796 20260 32824
rect 20254 32784 20260 32796
rect 20312 32784 20318 32836
rect 22281 32827 22339 32833
rect 22281 32824 22293 32827
rect 21482 32796 22293 32824
rect 22281 32793 22293 32796
rect 22327 32793 22339 32827
rect 24762 32824 24768 32836
rect 24723 32796 24768 32824
rect 22281 32787 22339 32793
rect 24762 32784 24768 32796
rect 24820 32784 24826 32836
rect 27249 32827 27307 32833
rect 27249 32793 27261 32827
rect 27295 32824 27307 32827
rect 27798 32824 27804 32836
rect 27295 32796 27804 32824
rect 27295 32793 27307 32796
rect 27249 32787 27307 32793
rect 27798 32784 27804 32796
rect 27856 32784 27862 32836
rect 31570 32824 31576 32836
rect 28000 32796 31576 32824
rect 28000 32768 28028 32796
rect 31570 32784 31576 32796
rect 31628 32824 31634 32836
rect 31680 32824 31708 32855
rect 31846 32852 31852 32904
rect 31904 32892 31910 32904
rect 31904 32864 31949 32892
rect 31904 32852 31910 32864
rect 32030 32852 32036 32904
rect 32088 32892 32094 32904
rect 32858 32892 32864 32904
rect 32088 32864 32133 32892
rect 32819 32864 32864 32892
rect 32088 32852 32094 32864
rect 32858 32852 32864 32864
rect 32916 32852 32922 32904
rect 46290 32852 46296 32904
rect 46348 32892 46354 32904
rect 46569 32895 46627 32901
rect 46569 32892 46581 32895
rect 46348 32864 46581 32892
rect 46348 32852 46354 32864
rect 46569 32861 46581 32864
rect 46615 32861 46627 32895
rect 46569 32855 46627 32861
rect 31628 32796 31708 32824
rect 31628 32784 31634 32796
rect 47210 32784 47216 32836
rect 47268 32824 47274 32836
rect 47268 32796 47313 32824
rect 47268 32784 47274 32796
rect 17368 32728 17448 32756
rect 17368 32716 17374 32728
rect 17770 32716 17776 32768
rect 17828 32756 17834 32768
rect 17865 32759 17923 32765
rect 17865 32756 17877 32759
rect 17828 32728 17877 32756
rect 17828 32716 17834 32728
rect 17865 32725 17877 32728
rect 17911 32725 17923 32759
rect 17865 32719 17923 32725
rect 18506 32716 18512 32768
rect 18564 32756 18570 32768
rect 18601 32759 18659 32765
rect 18601 32756 18613 32759
rect 18564 32728 18613 32756
rect 18564 32716 18570 32728
rect 18601 32725 18613 32728
rect 18647 32725 18659 32759
rect 18601 32719 18659 32725
rect 21082 32716 21088 32768
rect 21140 32756 21146 32768
rect 21729 32759 21787 32765
rect 21729 32756 21741 32759
rect 21140 32728 21741 32756
rect 21140 32716 21146 32728
rect 21729 32725 21741 32728
rect 21775 32725 21787 32759
rect 21729 32719 21787 32725
rect 21818 32716 21824 32768
rect 21876 32756 21882 32768
rect 27982 32756 27988 32768
rect 21876 32728 27988 32756
rect 21876 32716 21882 32728
rect 27982 32716 27988 32728
rect 28040 32716 28046 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 15470 32512 15476 32564
rect 15528 32552 15534 32564
rect 17037 32555 17095 32561
rect 17037 32552 17049 32555
rect 15528 32524 17049 32552
rect 15528 32512 15534 32524
rect 17037 32521 17049 32524
rect 17083 32521 17095 32555
rect 17310 32552 17316 32564
rect 17037 32515 17095 32521
rect 17144 32524 17316 32552
rect 2222 32484 2228 32496
rect 2183 32456 2228 32484
rect 2222 32444 2228 32456
rect 2280 32444 2286 32496
rect 16390 32444 16396 32496
rect 16448 32484 16454 32496
rect 16853 32487 16911 32493
rect 16853 32484 16865 32487
rect 16448 32456 16865 32484
rect 16448 32444 16454 32456
rect 16853 32453 16865 32456
rect 16899 32484 16911 32487
rect 17144 32484 17172 32524
rect 17310 32512 17316 32524
rect 17368 32552 17374 32564
rect 19245 32555 19303 32561
rect 19245 32552 19257 32555
rect 17368 32524 19257 32552
rect 17368 32512 17374 32524
rect 19245 32521 19257 32524
rect 19291 32521 19303 32555
rect 19245 32515 19303 32521
rect 20254 32512 20260 32564
rect 20312 32552 20318 32564
rect 21269 32555 21327 32561
rect 21269 32552 21281 32555
rect 20312 32524 21281 32552
rect 20312 32512 20318 32524
rect 21269 32521 21281 32524
rect 21315 32521 21327 32555
rect 21269 32515 21327 32521
rect 24210 32512 24216 32564
rect 24268 32561 24274 32564
rect 24268 32555 24287 32561
rect 24275 32521 24287 32555
rect 24394 32552 24400 32564
rect 24355 32524 24400 32552
rect 24268 32515 24287 32521
rect 24268 32512 24274 32515
rect 24394 32512 24400 32524
rect 24452 32512 24458 32564
rect 27614 32512 27620 32564
rect 27672 32512 27678 32564
rect 29546 32552 29552 32564
rect 29507 32524 29552 32552
rect 29546 32512 29552 32524
rect 29604 32512 29610 32564
rect 31938 32512 31944 32564
rect 31996 32552 32002 32564
rect 48041 32555 48099 32561
rect 48041 32552 48053 32555
rect 31996 32524 48053 32552
rect 31996 32512 32002 32524
rect 48041 32521 48053 32524
rect 48087 32521 48099 32555
rect 48041 32515 48099 32521
rect 16899 32456 17172 32484
rect 16899 32453 16911 32456
rect 16853 32447 16911 32453
rect 17494 32444 17500 32496
rect 17552 32444 17558 32496
rect 17770 32484 17776 32496
rect 17731 32456 17776 32484
rect 17770 32444 17776 32456
rect 17828 32444 17834 32496
rect 18506 32444 18512 32496
rect 18564 32444 18570 32496
rect 20806 32444 20812 32496
rect 20864 32444 20870 32496
rect 20990 32444 20996 32496
rect 21048 32484 21054 32496
rect 21818 32484 21824 32496
rect 21048 32456 21824 32484
rect 21048 32444 21054 32456
rect 2038 32416 2044 32428
rect 1999 32388 2044 32416
rect 2038 32376 2044 32388
rect 2096 32376 2102 32428
rect 16206 32376 16212 32428
rect 16264 32416 16270 32428
rect 16669 32419 16727 32425
rect 16669 32416 16681 32419
rect 16264 32388 16681 32416
rect 16264 32376 16270 32388
rect 16669 32385 16681 32388
rect 16715 32385 16727 32419
rect 17512 32416 17540 32444
rect 16669 32379 16727 32385
rect 16776 32388 17540 32416
rect 3881 32351 3939 32357
rect 3881 32317 3893 32351
rect 3927 32348 3939 32351
rect 4706 32348 4712 32360
rect 3927 32320 4712 32348
rect 3927 32317 3939 32320
rect 3881 32311 3939 32317
rect 4706 32308 4712 32320
rect 4764 32308 4770 32360
rect 16574 32308 16580 32360
rect 16632 32348 16638 32360
rect 16776 32348 16804 32388
rect 20346 32376 20352 32428
rect 20404 32416 20410 32428
rect 20533 32419 20591 32425
rect 20533 32416 20545 32419
rect 20404 32388 20545 32416
rect 20404 32376 20410 32388
rect 20533 32385 20545 32388
rect 20579 32385 20591 32419
rect 20533 32379 20591 32385
rect 20717 32419 20775 32425
rect 20717 32385 20729 32419
rect 20763 32385 20775 32419
rect 20824 32416 20852 32444
rect 21082 32416 21088 32428
rect 20824 32388 21088 32416
rect 20717 32379 20775 32385
rect 16632 32320 16804 32348
rect 17497 32351 17555 32357
rect 16632 32308 16638 32320
rect 17497 32317 17509 32351
rect 17543 32317 17555 32351
rect 17497 32311 17555 32317
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1581 32215 1639 32221
rect 1581 32212 1593 32215
rect 1452 32184 1593 32212
rect 1452 32172 1458 32184
rect 1581 32181 1593 32184
rect 1627 32181 1639 32215
rect 17512 32212 17540 32311
rect 19702 32308 19708 32360
rect 19760 32348 19766 32360
rect 20732 32348 20760 32379
rect 21082 32376 21088 32388
rect 21140 32376 21146 32428
rect 19760 32320 20760 32348
rect 19760 32308 19766 32320
rect 17862 32212 17868 32224
rect 17512 32184 17868 32212
rect 1581 32175 1639 32181
rect 17862 32172 17868 32184
rect 17920 32172 17926 32224
rect 20732 32212 20760 32320
rect 20809 32351 20867 32357
rect 20809 32317 20821 32351
rect 20855 32317 20867 32351
rect 20809 32311 20867 32317
rect 20901 32351 20959 32357
rect 20901 32317 20913 32351
rect 20947 32348 20959 32351
rect 21192 32348 21220 32456
rect 21818 32444 21824 32456
rect 21876 32444 21882 32496
rect 23106 32444 23112 32496
rect 23164 32484 23170 32496
rect 24029 32487 24087 32493
rect 24029 32484 24041 32487
rect 23164 32456 24041 32484
rect 23164 32444 23170 32456
rect 24029 32453 24041 32456
rect 24075 32484 24087 32487
rect 25406 32484 25412 32496
rect 24075 32456 25412 32484
rect 24075 32453 24087 32456
rect 24029 32447 24087 32453
rect 25406 32444 25412 32456
rect 25464 32444 25470 32496
rect 27632 32484 27660 32512
rect 26988 32456 27660 32484
rect 24946 32416 24952 32428
rect 24907 32388 24952 32416
rect 24946 32376 24952 32388
rect 25004 32376 25010 32428
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32416 25835 32419
rect 26050 32416 26056 32428
rect 25823 32388 26056 32416
rect 25823 32385 25835 32388
rect 25777 32379 25835 32385
rect 26050 32376 26056 32388
rect 26108 32416 26114 32428
rect 26694 32416 26700 32428
rect 26108 32388 26700 32416
rect 26108 32376 26114 32388
rect 26694 32376 26700 32388
rect 26752 32376 26758 32428
rect 26988 32425 27016 32456
rect 28258 32444 28264 32496
rect 28316 32444 28322 32496
rect 29181 32487 29239 32493
rect 29181 32453 29193 32487
rect 29227 32484 29239 32487
rect 29914 32484 29920 32496
rect 29227 32456 29920 32484
rect 29227 32453 29239 32456
rect 29181 32447 29239 32453
rect 29914 32444 29920 32456
rect 29972 32484 29978 32496
rect 29972 32456 30144 32484
rect 29972 32444 29978 32456
rect 26973 32419 27031 32425
rect 26973 32385 26985 32419
rect 27019 32385 27031 32419
rect 29365 32419 29423 32425
rect 29365 32416 29377 32419
rect 26973 32379 27031 32385
rect 28736 32388 29377 32416
rect 28736 32360 28764 32388
rect 29365 32385 29377 32388
rect 29411 32385 29423 32419
rect 29365 32379 29423 32385
rect 29822 32376 29828 32428
rect 29880 32416 29886 32428
rect 30116 32425 30144 32456
rect 32858 32444 32864 32496
rect 32916 32444 32922 32496
rect 30009 32419 30067 32425
rect 30009 32416 30021 32419
rect 29880 32388 30021 32416
rect 29880 32376 29886 32388
rect 30009 32385 30021 32388
rect 30055 32385 30067 32419
rect 30009 32379 30067 32385
rect 30101 32419 30159 32425
rect 30101 32385 30113 32419
rect 30147 32385 30159 32419
rect 32122 32416 32128 32428
rect 32083 32388 32128 32416
rect 30101 32379 30159 32385
rect 32122 32376 32128 32388
rect 32180 32376 32186 32428
rect 46658 32376 46664 32428
rect 46716 32416 46722 32428
rect 46845 32419 46903 32425
rect 46845 32416 46857 32419
rect 46716 32388 46857 32416
rect 46716 32376 46722 32388
rect 46845 32385 46857 32388
rect 46891 32416 46903 32419
rect 47578 32416 47584 32428
rect 46891 32388 47584 32416
rect 46891 32385 46903 32388
rect 46845 32379 46903 32385
rect 47578 32376 47584 32388
rect 47636 32376 47642 32428
rect 47946 32416 47952 32428
rect 47907 32388 47952 32416
rect 47946 32376 47952 32388
rect 48004 32376 48010 32428
rect 25682 32348 25688 32360
rect 20947 32320 21220 32348
rect 25643 32320 25688 32348
rect 20947 32317 20959 32320
rect 20901 32311 20959 32317
rect 20824 32280 20852 32311
rect 25682 32308 25688 32320
rect 25740 32308 25746 32360
rect 26786 32308 26792 32360
rect 26844 32348 26850 32360
rect 27249 32351 27307 32357
rect 27249 32348 27261 32351
rect 26844 32320 27261 32348
rect 26844 32308 26850 32320
rect 27249 32317 27261 32320
rect 27295 32317 27307 32351
rect 28718 32348 28724 32360
rect 28631 32320 28724 32348
rect 27249 32311 27307 32317
rect 28718 32308 28724 32320
rect 28776 32308 28782 32360
rect 32398 32348 32404 32360
rect 32359 32320 32404 32348
rect 32398 32308 32404 32320
rect 32456 32308 32462 32360
rect 20990 32280 20996 32292
rect 20824 32252 20996 32280
rect 20990 32240 20996 32252
rect 21048 32240 21054 32292
rect 24946 32280 24952 32292
rect 24228 32252 24952 32280
rect 24118 32212 24124 32224
rect 20732 32184 24124 32212
rect 24118 32172 24124 32184
rect 24176 32172 24182 32224
rect 24228 32221 24256 32252
rect 24946 32240 24952 32252
rect 25004 32240 25010 32292
rect 25130 32280 25136 32292
rect 25091 32252 25136 32280
rect 25130 32240 25136 32252
rect 25188 32240 25194 32292
rect 28350 32240 28356 32292
rect 28408 32280 28414 32292
rect 29178 32280 29184 32292
rect 28408 32252 29184 32280
rect 28408 32240 28414 32252
rect 29178 32240 29184 32252
rect 29236 32240 29242 32292
rect 24213 32215 24271 32221
rect 24213 32181 24225 32215
rect 24259 32181 24271 32215
rect 24213 32175 24271 32181
rect 25774 32172 25780 32224
rect 25832 32212 25838 32224
rect 26145 32215 26203 32221
rect 26145 32212 26157 32215
rect 25832 32184 26157 32212
rect 25832 32172 25838 32184
rect 26145 32181 26157 32184
rect 26191 32181 26203 32215
rect 26145 32175 26203 32181
rect 26234 32172 26240 32224
rect 26292 32212 26298 32224
rect 27706 32212 27712 32224
rect 26292 32184 27712 32212
rect 26292 32172 26298 32184
rect 27706 32172 27712 32184
rect 27764 32212 27770 32224
rect 28534 32212 28540 32224
rect 27764 32184 28540 32212
rect 27764 32172 27770 32184
rect 28534 32172 28540 32184
rect 28592 32172 28598 32224
rect 30098 32212 30104 32224
rect 30059 32184 30104 32212
rect 30098 32172 30104 32184
rect 30156 32172 30162 32224
rect 30374 32212 30380 32224
rect 30335 32184 30380 32212
rect 30374 32172 30380 32184
rect 30432 32172 30438 32224
rect 31754 32172 31760 32224
rect 31812 32212 31818 32224
rect 33873 32215 33931 32221
rect 33873 32212 33885 32215
rect 31812 32184 33885 32212
rect 31812 32172 31818 32184
rect 33873 32181 33885 32184
rect 33919 32181 33931 32215
rect 33873 32175 33931 32181
rect 46474 32172 46480 32224
rect 46532 32212 46538 32224
rect 46937 32215 46995 32221
rect 46937 32212 46949 32215
rect 46532 32184 46949 32212
rect 46532 32172 46538 32184
rect 46937 32181 46949 32184
rect 46983 32181 46995 32215
rect 46937 32175 46995 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 15194 31968 15200 32020
rect 15252 32008 15258 32020
rect 15252 31980 17632 32008
rect 15252 31968 15258 31980
rect 17037 31943 17095 31949
rect 17037 31909 17049 31943
rect 17083 31940 17095 31943
rect 17494 31940 17500 31952
rect 17083 31912 17500 31940
rect 17083 31909 17095 31912
rect 17037 31903 17095 31909
rect 17494 31900 17500 31912
rect 17552 31900 17558 31952
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 14369 31875 14427 31881
rect 14369 31841 14381 31875
rect 14415 31872 14427 31875
rect 14458 31872 14464 31884
rect 14415 31844 14464 31872
rect 14415 31841 14427 31844
rect 14369 31835 14427 31841
rect 14458 31832 14464 31844
rect 14516 31832 14522 31884
rect 14550 31832 14556 31884
rect 14608 31872 14614 31884
rect 14645 31875 14703 31881
rect 14645 31872 14657 31875
rect 14608 31844 14657 31872
rect 14608 31832 14614 31844
rect 14645 31841 14657 31844
rect 14691 31841 14703 31875
rect 15841 31875 15899 31881
rect 15841 31872 15853 31875
rect 14645 31835 14703 31841
rect 14844 31844 15853 31872
rect 14277 31807 14335 31813
rect 14277 31773 14289 31807
rect 14323 31804 14335 31807
rect 14844 31804 14872 31844
rect 15841 31841 15853 31844
rect 15887 31841 15899 31875
rect 15841 31835 15899 31841
rect 16850 31832 16856 31884
rect 16908 31872 16914 31884
rect 16908 31844 17264 31872
rect 16908 31832 16914 31844
rect 17236 31816 17264 31844
rect 14323 31776 14872 31804
rect 14323 31773 14335 31776
rect 14277 31767 14335 31773
rect 14384 31748 14412 31776
rect 15562 31764 15568 31816
rect 15620 31804 15626 31816
rect 15657 31807 15715 31813
rect 15657 31804 15669 31807
rect 15620 31776 15669 31804
rect 15620 31764 15626 31776
rect 15657 31773 15669 31776
rect 15703 31804 15715 31807
rect 16482 31804 16488 31816
rect 15703 31776 16488 31804
rect 15703 31773 15715 31776
rect 15657 31767 15715 31773
rect 16482 31764 16488 31776
rect 16540 31764 16546 31816
rect 16942 31764 16948 31816
rect 17000 31804 17006 31816
rect 17037 31807 17095 31813
rect 17037 31804 17049 31807
rect 17000 31776 17049 31804
rect 17000 31764 17006 31776
rect 17037 31773 17049 31776
rect 17083 31773 17095 31807
rect 17037 31767 17095 31773
rect 17218 31764 17224 31816
rect 17276 31804 17282 31816
rect 17276 31776 17321 31804
rect 17276 31764 17282 31776
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 14366 31696 14372 31748
rect 14424 31696 14430 31748
rect 17604 31736 17632 31980
rect 17862 31968 17868 32020
rect 17920 32008 17926 32020
rect 19889 32011 19947 32017
rect 19889 32008 19901 32011
rect 17920 31980 19901 32008
rect 17920 31968 17926 31980
rect 19889 31977 19901 31980
rect 19935 32008 19947 32011
rect 19978 32008 19984 32020
rect 19935 31980 19984 32008
rect 19935 31977 19947 31980
rect 19889 31971 19947 31977
rect 19978 31968 19984 31980
rect 20036 31968 20042 32020
rect 23293 32011 23351 32017
rect 20088 31980 22094 32008
rect 17678 31900 17684 31952
rect 17736 31940 17742 31952
rect 20088 31940 20116 31980
rect 20898 31940 20904 31952
rect 17736 31912 20116 31940
rect 20456 31912 20904 31940
rect 17736 31900 17742 31912
rect 18414 31872 18420 31884
rect 17696 31844 18420 31872
rect 17696 31813 17724 31844
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 17681 31807 17739 31813
rect 17681 31773 17693 31807
rect 17727 31773 17739 31807
rect 17681 31767 17739 31773
rect 17773 31807 17831 31813
rect 17773 31773 17785 31807
rect 17819 31804 17831 31807
rect 17954 31804 17960 31816
rect 17819 31776 17960 31804
rect 17819 31773 17831 31776
rect 17773 31767 17831 31773
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 19702 31804 19708 31816
rect 18064 31776 19708 31804
rect 18064 31736 18092 31776
rect 19702 31764 19708 31776
rect 19760 31764 19766 31816
rect 19797 31807 19855 31813
rect 19797 31773 19809 31807
rect 19843 31804 19855 31807
rect 20456 31804 20484 31912
rect 20898 31900 20904 31912
rect 20956 31900 20962 31952
rect 20990 31900 20996 31952
rect 21048 31940 21054 31952
rect 21048 31912 21093 31940
rect 21048 31900 21054 31912
rect 20533 31875 20591 31881
rect 20533 31841 20545 31875
rect 20579 31841 20591 31875
rect 20533 31835 20591 31841
rect 19843 31776 20484 31804
rect 19843 31773 19855 31776
rect 19797 31767 19855 31773
rect 17604 31708 18092 31736
rect 20548 31736 20576 31835
rect 20625 31807 20683 31813
rect 20625 31773 20637 31807
rect 20671 31804 20683 31807
rect 20806 31804 20812 31816
rect 20671 31776 20812 31804
rect 20671 31773 20683 31776
rect 20625 31767 20683 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 22066 31804 22094 31980
rect 23293 31977 23305 32011
rect 23339 31977 23351 32011
rect 23474 32008 23480 32020
rect 23435 31980 23480 32008
rect 23293 31971 23351 31977
rect 23308 31940 23336 31971
rect 23474 31968 23480 31980
rect 23532 31968 23538 32020
rect 24854 32008 24860 32020
rect 24228 31980 24860 32008
rect 24228 31952 24256 31980
rect 24854 31968 24860 31980
rect 24912 31968 24918 32020
rect 24946 31968 24952 32020
rect 25004 32008 25010 32020
rect 25777 32011 25835 32017
rect 25777 32008 25789 32011
rect 25004 31980 25789 32008
rect 25004 31968 25010 31980
rect 25777 31977 25789 31980
rect 25823 31977 25835 32011
rect 26786 32008 26792 32020
rect 26747 31980 26792 32008
rect 25777 31971 25835 31977
rect 26786 31968 26792 31980
rect 26844 31968 26850 32020
rect 28813 32011 28871 32017
rect 26896 31980 28672 32008
rect 23566 31940 23572 31952
rect 23308 31912 23572 31940
rect 23566 31900 23572 31912
rect 23624 31940 23630 31952
rect 24210 31940 24216 31952
rect 23624 31912 24216 31940
rect 23624 31900 23630 31912
rect 24210 31900 24216 31912
rect 24268 31900 24274 31952
rect 24394 31900 24400 31952
rect 24452 31940 24458 31952
rect 26896 31940 26924 31980
rect 27801 31943 27859 31949
rect 27801 31940 27813 31943
rect 24452 31912 26924 31940
rect 27172 31912 27813 31940
rect 24452 31900 24458 31912
rect 24765 31875 24823 31881
rect 24765 31841 24777 31875
rect 24811 31872 24823 31875
rect 25498 31872 25504 31884
rect 24811 31844 25504 31872
rect 24811 31841 24823 31844
rect 24765 31835 24823 31841
rect 25498 31832 25504 31844
rect 25556 31872 25562 31884
rect 26142 31872 26148 31884
rect 25556 31844 26148 31872
rect 25556 31832 25562 31844
rect 26142 31832 26148 31844
rect 26200 31832 26206 31884
rect 27172 31813 27200 31912
rect 27801 31909 27813 31912
rect 27847 31909 27859 31943
rect 28350 31940 28356 31952
rect 27801 31903 27859 31909
rect 28184 31912 28356 31940
rect 27246 31832 27252 31884
rect 27304 31872 27310 31884
rect 27304 31844 27349 31872
rect 27304 31832 27310 31844
rect 24949 31807 25007 31813
rect 22066 31776 23244 31804
rect 23216 31770 23244 31776
rect 23339 31773 23397 31779
rect 23339 31770 23351 31773
rect 20898 31736 20904 31748
rect 20548 31708 20904 31736
rect 20898 31696 20904 31708
rect 20956 31696 20962 31748
rect 23106 31736 23112 31748
rect 23067 31708 23112 31736
rect 23106 31696 23112 31708
rect 23164 31696 23170 31748
rect 23216 31742 23351 31770
rect 23339 31739 23351 31742
rect 23385 31739 23397 31773
rect 24949 31773 24961 31807
rect 24995 31804 25007 31807
rect 25685 31807 25743 31813
rect 25685 31804 25697 31807
rect 24995 31776 25697 31804
rect 24995 31773 25007 31776
rect 24949 31767 25007 31773
rect 25685 31773 25697 31776
rect 25731 31773 25743 31807
rect 25685 31767 25743 31773
rect 26973 31807 27031 31813
rect 26973 31773 26985 31807
rect 27019 31804 27031 31807
rect 27125 31807 27200 31813
rect 27019 31776 27053 31804
rect 27019 31773 27031 31776
rect 26973 31767 27031 31773
rect 27125 31773 27137 31807
rect 27171 31776 27200 31807
rect 27338 31804 27344 31816
rect 27251 31776 27344 31804
rect 27171 31773 27183 31776
rect 27125 31767 27183 31773
rect 23339 31733 23397 31739
rect 24854 31696 24860 31748
rect 24912 31736 24918 31748
rect 24964 31736 24992 31767
rect 25225 31739 25283 31745
rect 25225 31736 25237 31739
rect 24912 31708 24992 31736
rect 25056 31708 25237 31736
rect 24912 31696 24918 31708
rect 20162 31628 20168 31680
rect 20220 31668 20226 31680
rect 22186 31668 22192 31680
rect 20220 31640 22192 31668
rect 20220 31628 20226 31640
rect 22186 31628 22192 31640
rect 22244 31668 22250 31680
rect 22554 31668 22560 31680
rect 22244 31640 22560 31668
rect 22244 31628 22250 31640
rect 22554 31628 22560 31640
rect 22612 31628 22618 31680
rect 24946 31628 24952 31680
rect 25004 31668 25010 31680
rect 25056 31668 25084 31708
rect 25225 31705 25237 31708
rect 25271 31705 25283 31739
rect 25225 31699 25283 31705
rect 25004 31640 25084 31668
rect 25004 31628 25010 31640
rect 25130 31628 25136 31680
rect 25188 31668 25194 31680
rect 25406 31668 25412 31680
rect 25188 31640 25412 31668
rect 25188 31628 25194 31640
rect 25406 31628 25412 31640
rect 25464 31628 25470 31680
rect 25700 31668 25728 31767
rect 26988 31736 27016 31767
rect 27338 31764 27344 31776
rect 27396 31804 27402 31816
rect 27522 31804 27528 31816
rect 27396 31776 27528 31804
rect 27396 31764 27402 31776
rect 27522 31764 27528 31776
rect 27580 31764 27586 31816
rect 27982 31804 27988 31816
rect 27943 31776 27988 31804
rect 27982 31764 27988 31776
rect 28040 31764 28046 31816
rect 28077 31807 28135 31813
rect 28077 31773 28089 31807
rect 28123 31804 28135 31807
rect 28184 31804 28212 31912
rect 28350 31900 28356 31912
rect 28408 31900 28414 31952
rect 28644 31940 28672 31980
rect 28813 31977 28825 32011
rect 28859 32008 28871 32011
rect 29178 32008 29184 32020
rect 28859 31980 29184 32008
rect 28859 31977 28871 31980
rect 28813 31971 28871 31977
rect 29178 31968 29184 31980
rect 29236 31968 29242 32020
rect 30282 32008 30288 32020
rect 30243 31980 30288 32008
rect 30282 31968 30288 31980
rect 30340 31968 30346 32020
rect 32217 32011 32275 32017
rect 32217 31977 32229 32011
rect 32263 32008 32275 32011
rect 32398 32008 32404 32020
rect 32263 31980 32404 32008
rect 32263 31977 32275 31980
rect 32217 31971 32275 31977
rect 32398 31968 32404 31980
rect 32456 31968 32462 32020
rect 32858 32008 32864 32020
rect 32819 31980 32864 32008
rect 32858 31968 32864 31980
rect 32916 31968 32922 32020
rect 30561 31943 30619 31949
rect 28644 31912 30512 31940
rect 28261 31875 28319 31881
rect 28261 31841 28273 31875
rect 28307 31872 28319 31875
rect 28534 31872 28540 31884
rect 28307 31844 28540 31872
rect 28307 31841 28319 31844
rect 28261 31835 28319 31841
rect 28534 31832 28540 31844
rect 28592 31832 28598 31884
rect 28718 31832 28724 31884
rect 28776 31872 28782 31884
rect 28776 31844 29040 31872
rect 28776 31832 28782 31844
rect 28123 31776 28212 31804
rect 28353 31807 28411 31813
rect 28123 31773 28135 31776
rect 28077 31767 28135 31773
rect 28353 31773 28365 31807
rect 28399 31804 28411 31807
rect 28736 31804 28764 31832
rect 28399 31776 28764 31804
rect 28399 31773 28411 31776
rect 28353 31767 28411 31773
rect 28810 31764 28816 31816
rect 28868 31804 28874 31816
rect 29012 31813 29040 31844
rect 28997 31807 29055 31813
rect 28868 31776 28913 31804
rect 28868 31764 28874 31776
rect 28997 31773 29009 31807
rect 29043 31773 29055 31807
rect 28997 31767 29055 31773
rect 29822 31764 29828 31816
rect 29880 31804 29886 31816
rect 30006 31804 30012 31816
rect 29880 31776 30012 31804
rect 29880 31764 29886 31776
rect 30006 31764 30012 31776
rect 30064 31764 30070 31816
rect 30285 31807 30343 31813
rect 30285 31773 30297 31807
rect 30331 31804 30343 31807
rect 30484 31804 30512 31912
rect 30561 31909 30573 31943
rect 30607 31909 30619 31943
rect 40402 31940 40408 31952
rect 30561 31903 30619 31909
rect 31864 31912 40408 31940
rect 30331 31776 30512 31804
rect 30576 31804 30604 31903
rect 31754 31872 31760 31884
rect 31715 31844 31760 31872
rect 31754 31832 31760 31844
rect 31812 31832 31818 31884
rect 31864 31881 31892 31912
rect 40402 31900 40408 31912
rect 40460 31900 40466 31952
rect 31849 31875 31907 31881
rect 31849 31841 31861 31875
rect 31895 31841 31907 31875
rect 46290 31872 46296 31884
rect 46251 31844 46296 31872
rect 31849 31835 31907 31841
rect 46290 31832 46296 31844
rect 46348 31832 46354 31884
rect 46474 31872 46480 31884
rect 46435 31844 46480 31872
rect 46474 31832 46480 31844
rect 46532 31832 46538 31884
rect 48130 31872 48136 31884
rect 48091 31844 48136 31872
rect 48130 31832 48136 31844
rect 48188 31832 48194 31884
rect 31481 31807 31539 31813
rect 31481 31804 31493 31807
rect 30576 31776 31493 31804
rect 30331 31773 30343 31776
rect 30285 31767 30343 31773
rect 31481 31773 31493 31776
rect 31527 31773 31539 31807
rect 31481 31767 31539 31773
rect 31570 31764 31576 31816
rect 31628 31804 31634 31816
rect 31665 31807 31723 31813
rect 31665 31804 31677 31807
rect 31628 31776 31677 31804
rect 31628 31764 31634 31776
rect 31665 31773 31677 31776
rect 31711 31773 31723 31807
rect 32030 31804 32036 31816
rect 31991 31776 32036 31804
rect 31665 31767 31723 31773
rect 32030 31764 32036 31776
rect 32088 31764 32094 31816
rect 32122 31764 32128 31816
rect 32180 31804 32186 31816
rect 32766 31804 32772 31816
rect 32180 31776 32772 31804
rect 32180 31764 32186 31776
rect 32766 31764 32772 31776
rect 32824 31764 32830 31816
rect 28626 31736 28632 31748
rect 26988 31708 28632 31736
rect 28626 31696 28632 31708
rect 28684 31696 28690 31748
rect 28828 31736 28856 31764
rect 30374 31736 30380 31748
rect 28828 31708 30380 31736
rect 30374 31696 30380 31708
rect 30432 31696 30438 31748
rect 27522 31668 27528 31680
rect 25700 31640 27528 31668
rect 27522 31628 27528 31640
rect 27580 31628 27586 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 2225 31467 2283 31473
rect 2225 31464 2237 31467
rect 1636 31436 2237 31464
rect 1636 31424 1642 31436
rect 2225 31433 2237 31436
rect 2271 31433 2283 31467
rect 15562 31464 15568 31476
rect 15523 31436 15568 31464
rect 2225 31427 2283 31433
rect 15562 31424 15568 31436
rect 15620 31424 15626 31476
rect 24118 31424 24124 31476
rect 24176 31464 24182 31476
rect 24765 31467 24823 31473
rect 24765 31464 24777 31467
rect 24176 31436 24777 31464
rect 24176 31424 24182 31436
rect 24765 31433 24777 31436
rect 24811 31433 24823 31467
rect 24765 31427 24823 31433
rect 1946 31356 1952 31408
rect 2004 31396 2010 31408
rect 3053 31399 3111 31405
rect 3053 31396 3065 31399
rect 2004 31368 3065 31396
rect 2004 31356 2010 31368
rect 3053 31365 3065 31368
rect 3099 31365 3111 31399
rect 4706 31396 4712 31408
rect 4667 31368 4712 31396
rect 3053 31359 3111 31365
rect 4706 31356 4712 31368
rect 4764 31356 4770 31408
rect 15654 31396 15660 31408
rect 15318 31368 15660 31396
rect 15654 31356 15660 31368
rect 15712 31356 15718 31408
rect 20714 31396 20720 31408
rect 20675 31368 20720 31396
rect 20714 31356 20720 31368
rect 20772 31356 20778 31408
rect 24780 31396 24808 31427
rect 28626 31424 28632 31476
rect 28684 31464 28690 31476
rect 28905 31467 28963 31473
rect 28905 31464 28917 31467
rect 28684 31436 28917 31464
rect 28684 31424 28690 31436
rect 28905 31433 28917 31436
rect 28951 31433 28963 31467
rect 30098 31464 30104 31476
rect 28905 31427 28963 31433
rect 29656 31436 30104 31464
rect 24780 31368 26004 31396
rect 2133 31331 2191 31337
rect 2133 31297 2145 31331
rect 2179 31328 2191 31331
rect 2314 31328 2320 31340
rect 2179 31300 2320 31328
rect 2179 31297 2191 31300
rect 2133 31291 2191 31297
rect 2314 31288 2320 31300
rect 2372 31288 2378 31340
rect 17034 31328 17040 31340
rect 16995 31300 17040 31328
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 17865 31331 17923 31337
rect 17865 31297 17877 31331
rect 17911 31328 17923 31331
rect 18322 31328 18328 31340
rect 17911 31300 18328 31328
rect 17911 31297 17923 31300
rect 17865 31291 17923 31297
rect 18322 31288 18328 31300
rect 18380 31288 18386 31340
rect 20073 31331 20131 31337
rect 20073 31297 20085 31331
rect 20119 31328 20131 31331
rect 20162 31328 20168 31340
rect 20119 31300 20168 31328
rect 20119 31297 20131 31300
rect 20073 31291 20131 31297
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 20901 31331 20959 31337
rect 20901 31297 20913 31331
rect 20947 31328 20959 31331
rect 20990 31328 20996 31340
rect 20947 31300 20996 31328
rect 20947 31297 20959 31300
rect 20901 31291 20959 31297
rect 20990 31288 20996 31300
rect 21048 31288 21054 31340
rect 23566 31328 23572 31340
rect 23527 31300 23572 31328
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 24578 31328 24584 31340
rect 24539 31300 24584 31328
rect 24578 31288 24584 31300
rect 24636 31288 24642 31340
rect 25774 31328 25780 31340
rect 25735 31300 25780 31328
rect 25774 31288 25780 31300
rect 25832 31288 25838 31340
rect 25976 31337 26004 31368
rect 25961 31331 26019 31337
rect 25961 31297 25973 31331
rect 26007 31297 26019 31331
rect 25961 31291 26019 31297
rect 27430 31288 27436 31340
rect 27488 31328 27494 31340
rect 27525 31331 27583 31337
rect 27525 31328 27537 31331
rect 27488 31300 27537 31328
rect 27488 31288 27494 31300
rect 27525 31297 27537 31300
rect 27571 31297 27583 31331
rect 28626 31328 28632 31340
rect 28587 31300 28632 31328
rect 27525 31291 27583 31297
rect 28626 31288 28632 31300
rect 28684 31288 28690 31340
rect 28721 31331 28779 31337
rect 28721 31297 28733 31331
rect 28767 31328 28779 31331
rect 28810 31328 28816 31340
rect 28767 31300 28816 31328
rect 28767 31297 28779 31300
rect 28721 31291 28779 31297
rect 28810 31288 28816 31300
rect 28868 31288 28874 31340
rect 29656 31337 29684 31436
rect 30098 31424 30104 31436
rect 30156 31424 30162 31476
rect 30374 31424 30380 31476
rect 30432 31464 30438 31476
rect 30561 31467 30619 31473
rect 30561 31464 30573 31467
rect 30432 31436 30573 31464
rect 30432 31424 30438 31436
rect 30561 31433 30573 31436
rect 30607 31433 30619 31467
rect 30561 31427 30619 31433
rect 29917 31399 29975 31405
rect 29917 31365 29929 31399
rect 29963 31396 29975 31399
rect 29963 31368 30696 31396
rect 29963 31365 29975 31368
rect 29917 31359 29975 31365
rect 29641 31331 29699 31337
rect 29641 31297 29653 31331
rect 29687 31297 29699 31331
rect 29641 31291 29699 31297
rect 29733 31331 29791 31337
rect 29733 31297 29745 31331
rect 29779 31328 29791 31331
rect 30006 31328 30012 31340
rect 29779 31300 30012 31328
rect 29779 31297 29791 31300
rect 29733 31291 29791 31297
rect 30006 31288 30012 31300
rect 30064 31288 30070 31340
rect 30668 31337 30696 31368
rect 30377 31331 30435 31337
rect 30377 31297 30389 31331
rect 30423 31297 30435 31331
rect 30377 31291 30435 31297
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31297 30711 31331
rect 32122 31328 32128 31340
rect 32083 31300 32128 31328
rect 30653 31291 30711 31297
rect 2866 31260 2872 31272
rect 2827 31232 2872 31260
rect 2866 31220 2872 31232
rect 2924 31220 2930 31272
rect 13817 31263 13875 31269
rect 13817 31229 13829 31263
rect 13863 31260 13875 31263
rect 14093 31263 14151 31269
rect 13863 31232 13952 31260
rect 13863 31229 13875 31232
rect 13817 31223 13875 31229
rect 13924 31124 13952 31232
rect 14093 31229 14105 31263
rect 14139 31260 14151 31263
rect 15102 31260 15108 31272
rect 14139 31232 15108 31260
rect 14139 31229 14151 31232
rect 14093 31223 14151 31229
rect 15102 31220 15108 31232
rect 15160 31220 15166 31272
rect 16850 31260 16856 31272
rect 16811 31232 16856 31260
rect 16850 31220 16856 31232
rect 16908 31220 16914 31272
rect 23198 31220 23204 31272
rect 23256 31260 23262 31272
rect 23293 31263 23351 31269
rect 23293 31260 23305 31263
rect 23256 31232 23305 31260
rect 23256 31220 23262 31232
rect 23293 31229 23305 31232
rect 23339 31229 23351 31263
rect 29914 31260 29920 31272
rect 29875 31232 29920 31260
rect 23293 31223 23351 31229
rect 29914 31220 29920 31232
rect 29972 31220 29978 31272
rect 17034 31192 17040 31204
rect 15120 31164 17040 31192
rect 15120 31124 15148 31164
rect 17034 31152 17040 31164
rect 17092 31152 17098 31204
rect 17144 31164 22094 31192
rect 13924 31096 15148 31124
rect 16390 31084 16396 31136
rect 16448 31124 16454 31136
rect 17144 31124 17172 31164
rect 16448 31096 17172 31124
rect 17221 31127 17279 31133
rect 16448 31084 16454 31096
rect 17221 31093 17233 31127
rect 17267 31124 17279 31127
rect 17310 31124 17316 31136
rect 17267 31096 17316 31124
rect 17267 31093 17279 31096
rect 17221 31087 17279 31093
rect 17310 31084 17316 31096
rect 17368 31084 17374 31136
rect 18046 31124 18052 31136
rect 18007 31096 18052 31124
rect 18046 31084 18052 31096
rect 18104 31084 18110 31136
rect 20162 31124 20168 31136
rect 20123 31096 20168 31124
rect 20162 31084 20168 31096
rect 20220 31084 20226 31136
rect 20438 31084 20444 31136
rect 20496 31124 20502 31136
rect 20898 31124 20904 31136
rect 20496 31096 20904 31124
rect 20496 31084 20502 31096
rect 20898 31084 20904 31096
rect 20956 31124 20962 31136
rect 21085 31127 21143 31133
rect 21085 31124 21097 31127
rect 20956 31096 21097 31124
rect 20956 31084 20962 31096
rect 21085 31093 21097 31096
rect 21131 31093 21143 31127
rect 22066 31124 22094 31164
rect 23750 31152 23756 31204
rect 23808 31192 23814 31204
rect 27982 31192 27988 31204
rect 23808 31164 27988 31192
rect 23808 31152 23814 31164
rect 27982 31152 27988 31164
rect 28040 31152 28046 31204
rect 28718 31152 28724 31204
rect 28776 31192 28782 31204
rect 30392 31192 30420 31291
rect 32122 31288 32128 31300
rect 32180 31288 32186 31340
rect 28776 31164 30420 31192
rect 28776 31152 28782 31164
rect 24670 31124 24676 31136
rect 22066 31096 24676 31124
rect 21085 31087 21143 31093
rect 24670 31084 24676 31096
rect 24728 31124 24734 31136
rect 25406 31124 25412 31136
rect 24728 31096 25412 31124
rect 24728 31084 24734 31096
rect 25406 31084 25412 31096
rect 25464 31084 25470 31136
rect 25682 31084 25688 31136
rect 25740 31124 25746 31136
rect 25777 31127 25835 31133
rect 25777 31124 25789 31127
rect 25740 31096 25789 31124
rect 25740 31084 25746 31096
rect 25777 31093 25789 31096
rect 25823 31093 25835 31127
rect 27706 31124 27712 31136
rect 27667 31096 27712 31124
rect 25777 31087 25835 31093
rect 27706 31084 27712 31096
rect 27764 31084 27770 31136
rect 30098 31084 30104 31136
rect 30156 31124 30162 31136
rect 30377 31127 30435 31133
rect 30377 31124 30389 31127
rect 30156 31096 30389 31124
rect 30156 31084 30162 31096
rect 30377 31093 30389 31096
rect 30423 31093 30435 31127
rect 32214 31124 32220 31136
rect 32175 31096 32220 31124
rect 30377 31087 30435 31093
rect 32214 31084 32220 31096
rect 32272 31084 32278 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 15102 30920 15108 30932
rect 15063 30892 15108 30920
rect 15102 30880 15108 30892
rect 15160 30880 15166 30932
rect 15654 30920 15660 30932
rect 15615 30892 15660 30920
rect 15654 30880 15660 30892
rect 15712 30880 15718 30932
rect 16666 30880 16672 30932
rect 16724 30920 16730 30932
rect 17126 30920 17132 30932
rect 16724 30892 17132 30920
rect 16724 30880 16730 30892
rect 17126 30880 17132 30892
rect 17184 30880 17190 30932
rect 17310 30920 17316 30932
rect 17271 30892 17316 30920
rect 17310 30880 17316 30892
rect 17368 30880 17374 30932
rect 18414 30880 18420 30932
rect 18472 30920 18478 30932
rect 18509 30923 18567 30929
rect 18509 30920 18521 30923
rect 18472 30892 18521 30920
rect 18472 30880 18478 30892
rect 18509 30889 18521 30892
rect 18555 30889 18567 30923
rect 18509 30883 18567 30889
rect 20898 30880 20904 30932
rect 20956 30920 20962 30932
rect 21821 30923 21879 30929
rect 21821 30920 21833 30923
rect 20956 30892 21833 30920
rect 20956 30880 20962 30892
rect 21821 30889 21833 30892
rect 21867 30889 21879 30923
rect 21821 30883 21879 30889
rect 24765 30923 24823 30929
rect 24765 30889 24777 30923
rect 24811 30920 24823 30923
rect 24854 30920 24860 30932
rect 24811 30892 24860 30920
rect 24811 30889 24823 30892
rect 24765 30883 24823 30889
rect 24854 30880 24860 30892
rect 24912 30880 24918 30932
rect 25406 30880 25412 30932
rect 25464 30920 25470 30932
rect 28905 30923 28963 30929
rect 28905 30920 28917 30923
rect 25464 30892 28917 30920
rect 25464 30880 25470 30892
rect 28905 30889 28917 30892
rect 28951 30889 28963 30923
rect 28905 30883 28963 30889
rect 29914 30880 29920 30932
rect 29972 30920 29978 30932
rect 32585 30923 32643 30929
rect 32585 30920 32597 30923
rect 29972 30892 32597 30920
rect 29972 30880 29978 30892
rect 32585 30889 32597 30892
rect 32631 30889 32643 30923
rect 32585 30883 32643 30889
rect 18046 30852 18052 30864
rect 15580 30824 18052 30852
rect 14366 30744 14372 30796
rect 14424 30784 14430 30796
rect 14424 30756 14596 30784
rect 14424 30744 14430 30756
rect 14458 30716 14464 30728
rect 14419 30688 14464 30716
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 14568 30725 14596 30756
rect 15010 30725 15016 30728
rect 14554 30719 14612 30725
rect 14554 30685 14566 30719
rect 14600 30685 14612 30719
rect 14554 30679 14612 30685
rect 14967 30719 15016 30725
rect 14967 30685 14979 30719
rect 15013 30685 15016 30719
rect 14967 30679 15016 30685
rect 15010 30676 15016 30679
rect 15068 30676 15074 30728
rect 15580 30725 15608 30824
rect 18046 30812 18052 30824
rect 18104 30812 18110 30864
rect 24578 30852 24584 30864
rect 23584 30824 24584 30852
rect 17034 30744 17040 30796
rect 17092 30784 17098 30796
rect 17862 30784 17868 30796
rect 17092 30756 17868 30784
rect 17092 30744 17098 30756
rect 17862 30744 17868 30756
rect 17920 30784 17926 30796
rect 19245 30787 19303 30793
rect 19245 30784 19257 30787
rect 17920 30756 19257 30784
rect 17920 30744 17926 30756
rect 19245 30753 19257 30756
rect 19291 30753 19303 30787
rect 19245 30747 19303 30753
rect 19521 30787 19579 30793
rect 19521 30753 19533 30787
rect 19567 30784 19579 30787
rect 20530 30784 20536 30796
rect 19567 30756 20536 30784
rect 19567 30753 19579 30756
rect 19521 30747 19579 30753
rect 20530 30744 20536 30756
rect 20588 30744 20594 30796
rect 20806 30744 20812 30796
rect 20864 30784 20870 30796
rect 21266 30784 21272 30796
rect 20864 30756 21272 30784
rect 20864 30744 20870 30756
rect 21266 30744 21272 30756
rect 21324 30784 21330 30796
rect 21913 30787 21971 30793
rect 21913 30784 21925 30787
rect 21324 30756 21925 30784
rect 21324 30744 21330 30756
rect 21913 30753 21925 30756
rect 21959 30753 21971 30787
rect 21913 30747 21971 30753
rect 15565 30719 15623 30725
rect 15565 30685 15577 30719
rect 15611 30685 15623 30719
rect 15565 30679 15623 30685
rect 17129 30719 17187 30725
rect 17129 30685 17141 30719
rect 17175 30685 17187 30719
rect 17129 30679 17187 30685
rect 17405 30719 17463 30725
rect 17405 30685 17417 30719
rect 17451 30716 17463 30719
rect 17494 30716 17500 30728
rect 17451 30688 17500 30716
rect 17451 30685 17463 30688
rect 17405 30679 17463 30685
rect 14737 30651 14795 30657
rect 14737 30617 14749 30651
rect 14783 30617 14795 30651
rect 14737 30611 14795 30617
rect 14829 30651 14887 30657
rect 14829 30617 14841 30651
rect 14875 30648 14887 30651
rect 16390 30648 16396 30660
rect 14875 30620 16396 30648
rect 14875 30617 14887 30620
rect 14829 30611 14887 30617
rect 14752 30580 14780 30611
rect 16390 30608 16396 30620
rect 16448 30608 16454 30660
rect 16298 30580 16304 30592
rect 14752 30552 16304 30580
rect 16298 30540 16304 30552
rect 16356 30540 16362 30592
rect 16574 30540 16580 30592
rect 16632 30580 16638 30592
rect 16945 30583 17003 30589
rect 16945 30580 16957 30583
rect 16632 30552 16957 30580
rect 16632 30540 16638 30552
rect 16945 30549 16957 30552
rect 16991 30549 17003 30583
rect 17144 30580 17172 30679
rect 17494 30676 17500 30688
rect 17552 30676 17558 30728
rect 18322 30716 18328 30728
rect 18235 30688 18328 30716
rect 18322 30676 18328 30688
rect 18380 30716 18386 30728
rect 18782 30716 18788 30728
rect 18380 30688 18788 30716
rect 18380 30676 18386 30688
rect 18782 30676 18788 30688
rect 18840 30676 18846 30728
rect 21634 30716 21640 30728
rect 21595 30688 21640 30716
rect 21634 30676 21640 30688
rect 21692 30676 21698 30728
rect 22554 30716 22560 30728
rect 22515 30688 22560 30716
rect 22554 30676 22560 30688
rect 22612 30676 22618 30728
rect 23584 30725 23612 30824
rect 24578 30812 24584 30824
rect 24636 30852 24642 30864
rect 24949 30855 25007 30861
rect 24949 30852 24961 30855
rect 24636 30824 24961 30852
rect 24636 30812 24642 30824
rect 24949 30821 24961 30824
rect 24995 30821 25007 30855
rect 24949 30815 25007 30821
rect 29638 30812 29644 30864
rect 29696 30852 29702 30864
rect 30006 30852 30012 30864
rect 29696 30824 30012 30852
rect 29696 30812 29702 30824
rect 30006 30812 30012 30824
rect 30064 30812 30070 30864
rect 23658 30744 23664 30796
rect 23716 30784 23722 30796
rect 25409 30787 25467 30793
rect 25409 30784 25421 30787
rect 23716 30756 25421 30784
rect 23716 30744 23722 30756
rect 25409 30753 25421 30756
rect 25455 30784 25467 30787
rect 27985 30787 28043 30793
rect 27985 30784 27997 30787
rect 25455 30756 27997 30784
rect 25455 30753 25467 30756
rect 25409 30747 25467 30753
rect 27985 30753 27997 30756
rect 28031 30784 28043 30787
rect 29546 30784 29552 30796
rect 28031 30756 29552 30784
rect 28031 30753 28043 30756
rect 27985 30747 28043 30753
rect 29546 30744 29552 30756
rect 29604 30784 29610 30796
rect 30837 30787 30895 30793
rect 30837 30784 30849 30787
rect 29604 30756 30849 30784
rect 29604 30744 29610 30756
rect 30837 30753 30849 30756
rect 30883 30753 30895 30787
rect 30837 30747 30895 30753
rect 43070 30744 43076 30796
rect 43128 30784 43134 30796
rect 47121 30787 47179 30793
rect 47121 30784 47133 30787
rect 43128 30756 47133 30784
rect 43128 30744 43134 30756
rect 47121 30753 47133 30756
rect 47167 30784 47179 30787
rect 47670 30784 47676 30796
rect 47167 30756 47676 30784
rect 47167 30753 47179 30756
rect 47121 30747 47179 30753
rect 47670 30744 47676 30756
rect 47728 30744 47734 30796
rect 23569 30719 23627 30725
rect 23569 30685 23581 30719
rect 23615 30685 23627 30719
rect 23569 30679 23627 30685
rect 24397 30719 24455 30725
rect 24397 30685 24409 30719
rect 24443 30685 24455 30719
rect 24397 30679 24455 30685
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30716 24823 30719
rect 24854 30716 24860 30728
rect 24811 30688 24860 30716
rect 24811 30685 24823 30688
rect 24765 30679 24823 30685
rect 20162 30608 20168 30660
rect 20220 30608 20226 30660
rect 22204 30620 22876 30648
rect 20806 30580 20812 30592
rect 17144 30552 20812 30580
rect 16945 30543 17003 30549
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 20990 30580 20996 30592
rect 20951 30552 20996 30580
rect 20990 30540 20996 30552
rect 21048 30540 21054 30592
rect 21450 30580 21456 30592
rect 21411 30552 21456 30580
rect 21450 30540 21456 30552
rect 21508 30540 21514 30592
rect 22094 30540 22100 30592
rect 22152 30580 22158 30592
rect 22204 30580 22232 30620
rect 22152 30552 22232 30580
rect 22649 30583 22707 30589
rect 22152 30540 22158 30552
rect 22649 30549 22661 30583
rect 22695 30580 22707 30583
rect 22738 30580 22744 30592
rect 22695 30552 22744 30580
rect 22695 30549 22707 30552
rect 22649 30543 22707 30549
rect 22738 30540 22744 30552
rect 22796 30540 22802 30592
rect 22848 30580 22876 30620
rect 23198 30608 23204 30660
rect 23256 30648 23262 30660
rect 24412 30648 24440 30679
rect 24854 30676 24860 30688
rect 24912 30716 24918 30728
rect 25314 30716 25320 30728
rect 24912 30688 25320 30716
rect 24912 30676 24918 30688
rect 25314 30676 25320 30688
rect 25372 30676 25378 30728
rect 27798 30716 27804 30728
rect 27759 30688 27804 30716
rect 27798 30676 27804 30688
rect 27856 30676 27862 30728
rect 28718 30716 28724 30728
rect 28679 30688 28724 30716
rect 28718 30676 28724 30688
rect 28776 30676 28782 30728
rect 29733 30719 29791 30725
rect 29733 30685 29745 30719
rect 29779 30685 29791 30719
rect 29733 30679 29791 30685
rect 23256 30620 24440 30648
rect 25685 30651 25743 30657
rect 23256 30608 23262 30620
rect 25685 30617 25697 30651
rect 25731 30617 25743 30651
rect 27062 30648 27068 30660
rect 26910 30620 27068 30648
rect 25685 30611 25743 30617
rect 23750 30580 23756 30592
rect 22848 30552 23756 30580
rect 23750 30540 23756 30552
rect 23808 30540 23814 30592
rect 25700 30580 25728 30611
rect 27062 30608 27068 30620
rect 27120 30608 27126 30660
rect 26326 30580 26332 30592
rect 25700 30552 26332 30580
rect 26326 30540 26332 30552
rect 26384 30540 26390 30592
rect 26694 30540 26700 30592
rect 26752 30580 26758 30592
rect 27157 30583 27215 30589
rect 27157 30580 27169 30583
rect 26752 30552 27169 30580
rect 26752 30540 26758 30552
rect 27157 30549 27169 30552
rect 27203 30549 27215 30583
rect 27157 30543 27215 30549
rect 29549 30583 29607 30589
rect 29549 30549 29561 30583
rect 29595 30580 29607 30583
rect 29638 30580 29644 30592
rect 29595 30552 29644 30580
rect 29595 30549 29607 30552
rect 29549 30543 29607 30549
rect 29638 30540 29644 30552
rect 29696 30540 29702 30592
rect 29748 30580 29776 30679
rect 29822 30676 29828 30728
rect 29880 30716 29886 30728
rect 30006 30716 30012 30728
rect 29880 30688 29925 30716
rect 29967 30688 30012 30716
rect 29880 30676 29886 30688
rect 30006 30676 30012 30688
rect 30064 30676 30070 30728
rect 30098 30676 30104 30728
rect 30156 30716 30162 30728
rect 30156 30688 30201 30716
rect 30156 30676 30162 30688
rect 32214 30676 32220 30728
rect 32272 30676 32278 30728
rect 31110 30648 31116 30660
rect 31071 30620 31116 30648
rect 31110 30608 31116 30620
rect 31168 30608 31174 30660
rect 45738 30608 45744 30660
rect 45796 30648 45802 30660
rect 46845 30651 46903 30657
rect 46845 30648 46857 30651
rect 45796 30620 46857 30648
rect 45796 30608 45802 30620
rect 46845 30617 46857 30620
rect 46891 30617 46903 30651
rect 46845 30611 46903 30617
rect 46937 30651 46995 30657
rect 46937 30617 46949 30651
rect 46983 30617 46995 30651
rect 46937 30611 46995 30617
rect 43346 30580 43352 30592
rect 29748 30552 43352 30580
rect 43346 30540 43352 30552
rect 43404 30540 43410 30592
rect 46952 30580 46980 30611
rect 48222 30580 48228 30592
rect 46952 30552 48228 30580
rect 48222 30540 48228 30552
rect 48280 30540 48286 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 14458 30336 14464 30388
rect 14516 30376 14522 30388
rect 14645 30379 14703 30385
rect 14645 30376 14657 30379
rect 14516 30348 14657 30376
rect 14516 30336 14522 30348
rect 14645 30345 14657 30348
rect 14691 30345 14703 30379
rect 14645 30339 14703 30345
rect 16850 30336 16856 30388
rect 16908 30376 16914 30388
rect 18417 30379 18475 30385
rect 18417 30376 18429 30379
rect 16908 30348 18429 30376
rect 16908 30336 16914 30348
rect 18417 30345 18429 30348
rect 18463 30345 18475 30379
rect 20438 30376 20444 30388
rect 18417 30339 18475 30345
rect 19904 30348 20444 30376
rect 17954 30268 17960 30320
rect 18012 30268 18018 30320
rect 19904 30308 19932 30348
rect 20438 30336 20444 30348
rect 20496 30336 20502 30388
rect 20530 30336 20536 30388
rect 20588 30376 20594 30388
rect 20625 30379 20683 30385
rect 20625 30376 20637 30379
rect 20588 30348 20637 30376
rect 20588 30336 20594 30348
rect 20625 30345 20637 30348
rect 20671 30345 20683 30379
rect 26050 30376 26056 30388
rect 20625 30339 20683 30345
rect 25848 30348 26056 30376
rect 20349 30311 20407 30317
rect 19536 30280 19932 30308
rect 19996 30280 20208 30308
rect 14550 30240 14556 30252
rect 14511 30212 14556 30240
rect 14550 30200 14556 30212
rect 14608 30200 14614 30252
rect 14734 30240 14740 30252
rect 14695 30212 14740 30240
rect 14734 30200 14740 30212
rect 14792 30200 14798 30252
rect 19536 30249 19564 30280
rect 19996 30249 20024 30280
rect 19337 30243 19395 30249
rect 19337 30209 19349 30243
rect 19383 30209 19395 30243
rect 19337 30203 19395 30209
rect 19521 30243 19579 30249
rect 19521 30209 19533 30243
rect 19567 30209 19579 30243
rect 19521 30203 19579 30209
rect 19981 30243 20039 30249
rect 19981 30209 19993 30243
rect 20027 30209 20039 30243
rect 19981 30203 20039 30209
rect 20074 30243 20132 30249
rect 20074 30209 20086 30243
rect 20120 30209 20132 30243
rect 20074 30203 20132 30209
rect 16669 30175 16727 30181
rect 16669 30141 16681 30175
rect 16715 30172 16727 30175
rect 16942 30172 16948 30184
rect 16715 30144 16804 30172
rect 16903 30144 16948 30172
rect 16715 30141 16727 30144
rect 16669 30135 16727 30141
rect 16776 30036 16804 30144
rect 16942 30132 16948 30144
rect 17000 30132 17006 30184
rect 17034 30036 17040 30048
rect 16776 30008 17040 30036
rect 17034 29996 17040 30008
rect 17092 29996 17098 30048
rect 19352 30036 19380 30203
rect 19429 30175 19487 30181
rect 19429 30141 19441 30175
rect 19475 30172 19487 30175
rect 20088 30172 20116 30203
rect 19475 30144 20116 30172
rect 19475 30141 19487 30144
rect 19429 30135 19487 30141
rect 20180 30104 20208 30280
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 20714 30308 20720 30320
rect 20395 30280 20720 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 20714 30268 20720 30280
rect 20772 30308 20778 30320
rect 20990 30308 20996 30320
rect 20772 30280 20996 30308
rect 20772 30268 20778 30280
rect 20990 30268 20996 30280
rect 21048 30308 21054 30320
rect 21048 30280 21312 30308
rect 21048 30268 21054 30280
rect 20530 30249 20536 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30209 20315 30243
rect 20257 30203 20315 30209
rect 20487 30243 20536 30249
rect 20487 30209 20499 30243
rect 20533 30209 20536 30243
rect 20487 30203 20536 30209
rect 20272 30172 20300 30203
rect 20530 30200 20536 30203
rect 20588 30200 20594 30252
rect 20806 30200 20812 30252
rect 20864 30240 20870 30252
rect 21085 30243 21143 30249
rect 21085 30240 21097 30243
rect 20864 30212 21097 30240
rect 20864 30200 20870 30212
rect 21085 30209 21097 30212
rect 21131 30240 21143 30243
rect 21174 30240 21180 30252
rect 21131 30212 21180 30240
rect 21131 30209 21143 30212
rect 21085 30203 21143 30209
rect 21174 30200 21180 30212
rect 21232 30200 21238 30252
rect 21284 30249 21312 30280
rect 22738 30268 22744 30320
rect 22796 30268 22802 30320
rect 24305 30311 24363 30317
rect 24305 30277 24317 30311
rect 24351 30308 24363 30311
rect 24578 30308 24584 30320
rect 24351 30280 24584 30308
rect 24351 30277 24363 30280
rect 24305 30271 24363 30277
rect 24578 30268 24584 30280
rect 24636 30268 24642 30320
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30209 21327 30243
rect 21269 30203 21327 30209
rect 24394 30200 24400 30252
rect 24452 30240 24458 30252
rect 24489 30243 24547 30249
rect 24489 30240 24501 30243
rect 24452 30212 24501 30240
rect 24452 30200 24458 30212
rect 24489 30209 24501 30212
rect 24535 30209 24547 30243
rect 25682 30240 25688 30252
rect 25643 30212 25688 30240
rect 24489 30203 24547 30209
rect 25682 30200 25688 30212
rect 25740 30200 25746 30252
rect 25848 30249 25876 30348
rect 26050 30336 26056 30348
rect 26108 30376 26114 30388
rect 26326 30376 26332 30388
rect 26108 30348 26234 30376
rect 26287 30348 26332 30376
rect 26108 30336 26114 30348
rect 26206 30308 26234 30348
rect 26326 30336 26332 30348
rect 26384 30336 26390 30388
rect 27706 30336 27712 30388
rect 27764 30376 27770 30388
rect 32122 30376 32128 30388
rect 27764 30348 32128 30376
rect 27764 30336 27770 30348
rect 26694 30308 26700 30320
rect 26206 30280 26700 30308
rect 26694 30268 26700 30280
rect 26752 30268 26758 30320
rect 27062 30308 27068 30320
rect 27023 30280 27068 30308
rect 27062 30268 27068 30280
rect 27120 30268 27126 30320
rect 25833 30243 25891 30249
rect 25833 30209 25845 30243
rect 25879 30209 25891 30243
rect 25958 30240 25964 30252
rect 25919 30212 25964 30240
rect 25833 30203 25891 30209
rect 25958 30200 25964 30212
rect 26016 30200 26022 30252
rect 26050 30200 26056 30252
rect 26108 30240 26114 30252
rect 26191 30243 26249 30249
rect 26108 30212 26153 30240
rect 26108 30200 26114 30212
rect 26191 30209 26203 30243
rect 26237 30209 26249 30243
rect 26970 30240 26976 30252
rect 26931 30212 26976 30240
rect 26191 30203 26249 30209
rect 22005 30175 22063 30181
rect 20272 30144 20484 30172
rect 20456 30116 20484 30144
rect 22005 30141 22017 30175
rect 22051 30141 22063 30175
rect 22005 30135 22063 30141
rect 22281 30175 22339 30181
rect 22281 30141 22293 30175
rect 22327 30172 22339 30175
rect 22830 30172 22836 30184
rect 22327 30144 22836 30172
rect 22327 30141 22339 30144
rect 22281 30135 22339 30141
rect 20346 30104 20352 30116
rect 20180 30076 20352 30104
rect 20346 30064 20352 30076
rect 20404 30064 20410 30116
rect 20438 30064 20444 30116
rect 20496 30064 20502 30116
rect 21177 30039 21235 30045
rect 21177 30036 21189 30039
rect 19352 30008 21189 30036
rect 21177 30005 21189 30008
rect 21223 30005 21235 30039
rect 22020 30036 22048 30135
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 23382 30064 23388 30116
rect 23440 30104 23446 30116
rect 23440 30076 23980 30104
rect 23440 30064 23446 30076
rect 23658 30036 23664 30048
rect 22020 30008 23664 30036
rect 21177 29999 21235 30005
rect 23658 29996 23664 30008
rect 23716 29996 23722 30048
rect 23750 29996 23756 30048
rect 23808 30036 23814 30048
rect 23952 30036 23980 30076
rect 25498 30064 25504 30116
rect 25556 30104 25562 30116
rect 26206 30104 26234 30203
rect 26970 30200 26976 30212
rect 27028 30200 27034 30252
rect 28092 30249 28120 30348
rect 32122 30336 32128 30348
rect 32180 30336 32186 30388
rect 28169 30311 28227 30317
rect 28169 30277 28181 30311
rect 28215 30308 28227 30311
rect 28258 30308 28264 30320
rect 28215 30280 28264 30308
rect 28215 30277 28227 30280
rect 28169 30271 28227 30277
rect 28258 30268 28264 30280
rect 28316 30268 28322 30320
rect 29457 30311 29515 30317
rect 29457 30277 29469 30311
rect 29503 30308 29515 30311
rect 31110 30308 31116 30320
rect 29503 30280 31116 30308
rect 29503 30277 29515 30280
rect 29457 30271 29515 30277
rect 31110 30268 31116 30280
rect 31168 30268 31174 30320
rect 34514 30308 34520 30320
rect 32968 30280 34520 30308
rect 28077 30243 28135 30249
rect 28077 30209 28089 30243
rect 28123 30209 28135 30243
rect 29638 30240 29644 30252
rect 29599 30212 29644 30240
rect 28077 30203 28135 30209
rect 29638 30200 29644 30212
rect 29696 30200 29702 30252
rect 29914 30240 29920 30252
rect 29875 30212 29920 30240
rect 29914 30200 29920 30212
rect 29972 30200 29978 30252
rect 32968 30249 32996 30280
rect 34514 30268 34520 30280
rect 34572 30268 34578 30320
rect 32953 30243 33011 30249
rect 32953 30209 32965 30243
rect 32999 30209 33011 30243
rect 32953 30203 33011 30209
rect 29362 30132 29368 30184
rect 29420 30172 29426 30184
rect 29822 30172 29828 30184
rect 29420 30144 29828 30172
rect 29420 30132 29426 30144
rect 29822 30132 29828 30144
rect 29880 30132 29886 30184
rect 33134 30172 33140 30184
rect 33095 30144 33140 30172
rect 33134 30132 33140 30144
rect 33192 30132 33198 30184
rect 33413 30175 33471 30181
rect 33413 30141 33425 30175
rect 33459 30141 33471 30175
rect 33413 30135 33471 30141
rect 25556 30076 26234 30104
rect 25556 30064 25562 30076
rect 26326 30064 26332 30116
rect 26384 30104 26390 30116
rect 26384 30076 31754 30104
rect 26384 30064 26390 30076
rect 28994 30036 29000 30048
rect 23808 30008 23853 30036
rect 23952 30008 29000 30036
rect 23808 29996 23814 30008
rect 28994 29996 29000 30008
rect 29052 30036 29058 30048
rect 29825 30039 29883 30045
rect 29825 30036 29837 30039
rect 29052 30008 29837 30036
rect 29052 29996 29058 30008
rect 29825 30005 29837 30008
rect 29871 30005 29883 30039
rect 31726 30036 31754 30076
rect 33428 30036 33456 30135
rect 31726 30008 33456 30036
rect 29825 29999 29883 30005
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 16669 29835 16727 29841
rect 16669 29801 16681 29835
rect 16715 29832 16727 29835
rect 16942 29832 16948 29844
rect 16715 29804 16948 29832
rect 16715 29801 16727 29804
rect 16669 29795 16727 29801
rect 16942 29792 16948 29804
rect 17000 29792 17006 29844
rect 20162 29832 20168 29844
rect 19904 29804 20168 29832
rect 14734 29724 14740 29776
rect 14792 29764 14798 29776
rect 19904 29764 19932 29804
rect 20162 29792 20168 29804
rect 20220 29792 20226 29844
rect 20441 29835 20499 29841
rect 20441 29801 20453 29835
rect 20487 29832 20499 29835
rect 21266 29832 21272 29844
rect 20487 29804 21272 29832
rect 20487 29801 20499 29804
rect 20441 29795 20499 29801
rect 21266 29792 21272 29804
rect 21324 29792 21330 29844
rect 21450 29832 21456 29844
rect 21411 29804 21456 29832
rect 21450 29792 21456 29804
rect 21508 29792 21514 29844
rect 21542 29792 21548 29844
rect 21600 29832 21606 29844
rect 22830 29832 22836 29844
rect 21600 29804 22692 29832
rect 22791 29804 22836 29832
rect 21600 29792 21606 29804
rect 22664 29764 22692 29804
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 24581 29835 24639 29841
rect 24581 29801 24593 29835
rect 24627 29832 24639 29835
rect 27338 29832 27344 29844
rect 24627 29804 27344 29832
rect 24627 29801 24639 29804
rect 24581 29795 24639 29801
rect 24394 29764 24400 29776
rect 14792 29736 19932 29764
rect 21284 29736 21680 29764
rect 22664 29736 24400 29764
rect 14792 29724 14798 29736
rect 16574 29696 16580 29708
rect 16040 29668 16580 29696
rect 16040 29637 16068 29668
rect 16574 29656 16580 29668
rect 16632 29656 16638 29708
rect 20714 29696 20720 29708
rect 20272 29668 20720 29696
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29597 16083 29631
rect 16025 29591 16083 29597
rect 16173 29631 16231 29637
rect 16173 29597 16185 29631
rect 16219 29628 16231 29631
rect 16219 29597 16252 29628
rect 16173 29591 16252 29597
rect 16224 29492 16252 29591
rect 16298 29588 16304 29640
rect 16356 29628 16362 29640
rect 16356 29600 16401 29628
rect 16356 29588 16362 29600
rect 16482 29588 16488 29640
rect 16540 29637 16546 29640
rect 16540 29628 16548 29637
rect 17221 29631 17279 29637
rect 16540 29600 16585 29628
rect 16540 29591 16548 29600
rect 17221 29597 17233 29631
rect 17267 29597 17279 29631
rect 17221 29591 17279 29597
rect 17313 29631 17371 29637
rect 17313 29597 17325 29631
rect 17359 29628 17371 29631
rect 17402 29628 17408 29640
rect 17359 29600 17408 29628
rect 17359 29597 17371 29600
rect 17313 29591 17371 29597
rect 16540 29588 16546 29591
rect 16390 29560 16396 29572
rect 16351 29532 16396 29560
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 17236 29560 17264 29591
rect 17402 29588 17408 29600
rect 17460 29588 17466 29640
rect 20272 29637 20300 29668
rect 20714 29656 20720 29668
rect 20772 29656 20778 29708
rect 21284 29696 21312 29736
rect 21652 29708 21680 29736
rect 24394 29724 24400 29736
rect 24452 29724 24458 29776
rect 20916 29668 21312 29696
rect 21361 29699 21419 29705
rect 20257 29631 20315 29637
rect 20257 29597 20269 29631
rect 20303 29597 20315 29631
rect 20257 29591 20315 29597
rect 20441 29631 20499 29637
rect 20441 29597 20453 29631
rect 20487 29628 20499 29631
rect 20916 29628 20944 29668
rect 21361 29665 21373 29699
rect 21407 29696 21419 29699
rect 21542 29696 21548 29708
rect 21407 29668 21548 29696
rect 21407 29665 21419 29668
rect 21361 29659 21419 29665
rect 21542 29656 21548 29668
rect 21600 29656 21606 29708
rect 21634 29656 21640 29708
rect 21692 29696 21698 29708
rect 22373 29699 22431 29705
rect 22373 29696 22385 29699
rect 21692 29668 22385 29696
rect 21692 29656 21698 29668
rect 22373 29665 22385 29668
rect 22419 29696 22431 29699
rect 23750 29696 23756 29708
rect 22419 29668 23756 29696
rect 22419 29665 22431 29668
rect 22373 29659 22431 29665
rect 23750 29656 23756 29668
rect 23808 29656 23814 29708
rect 24596 29696 24624 29795
rect 27338 29792 27344 29804
rect 27396 29792 27402 29844
rect 29641 29835 29699 29841
rect 29641 29801 29653 29835
rect 29687 29801 29699 29835
rect 29641 29795 29699 29801
rect 28813 29767 28871 29773
rect 28813 29764 28825 29767
rect 23860 29668 24624 29696
rect 25148 29736 28825 29764
rect 21082 29628 21088 29640
rect 20487 29600 20944 29628
rect 21043 29600 21088 29628
rect 20487 29597 20499 29600
rect 20441 29591 20499 29597
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 22097 29631 22155 29637
rect 22097 29628 22109 29631
rect 21652 29600 22109 29628
rect 19978 29560 19984 29572
rect 17236 29532 19984 29560
rect 19978 29520 19984 29532
rect 20036 29520 20042 29572
rect 16850 29492 16856 29504
rect 16224 29464 16856 29492
rect 16850 29452 16856 29464
rect 16908 29452 16914 29504
rect 17310 29452 17316 29504
rect 17368 29492 17374 29504
rect 17497 29495 17555 29501
rect 17497 29492 17509 29495
rect 17368 29464 17509 29492
rect 17368 29452 17374 29464
rect 17497 29461 17509 29464
rect 17543 29461 17555 29495
rect 17497 29455 17555 29461
rect 20625 29495 20683 29501
rect 20625 29461 20637 29495
rect 20671 29492 20683 29495
rect 21450 29492 21456 29504
rect 20671 29464 21456 29492
rect 20671 29461 20683 29464
rect 20625 29455 20683 29461
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 21652 29501 21680 29600
rect 22097 29597 22109 29600
rect 22143 29597 22155 29631
rect 22097 29591 22155 29597
rect 22281 29631 22339 29637
rect 22281 29597 22293 29631
rect 22327 29597 22339 29631
rect 22462 29628 22468 29640
rect 22423 29600 22468 29628
rect 22281 29591 22339 29597
rect 21726 29520 21732 29572
rect 21784 29560 21790 29572
rect 22296 29560 22324 29591
rect 22462 29588 22468 29600
rect 22520 29588 22526 29640
rect 22646 29588 22652 29640
rect 22704 29628 22710 29640
rect 23860 29628 23888 29668
rect 22704 29600 23888 29628
rect 22704 29588 22710 29600
rect 24302 29588 24308 29640
rect 24360 29628 24366 29640
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 24360 29600 24409 29628
rect 24360 29588 24366 29600
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 24946 29588 24952 29640
rect 25004 29628 25010 29640
rect 25148 29637 25176 29736
rect 28813 29733 28825 29736
rect 28859 29764 28871 29767
rect 29362 29764 29368 29776
rect 28859 29736 29368 29764
rect 28859 29733 28871 29736
rect 28813 29727 28871 29733
rect 29362 29724 29368 29736
rect 29420 29724 29426 29776
rect 29656 29764 29684 29795
rect 29730 29792 29736 29844
rect 29788 29832 29794 29844
rect 30009 29835 30067 29841
rect 30009 29832 30021 29835
rect 29788 29804 30021 29832
rect 29788 29792 29794 29804
rect 30009 29801 30021 29804
rect 30055 29801 30067 29835
rect 33134 29832 33140 29844
rect 33095 29804 33140 29832
rect 30009 29795 30067 29801
rect 33134 29792 33140 29804
rect 33192 29792 33198 29844
rect 30374 29764 30380 29776
rect 29656 29736 30380 29764
rect 30374 29724 30380 29736
rect 30432 29724 30438 29776
rect 25314 29656 25320 29708
rect 25372 29696 25378 29708
rect 26326 29696 26332 29708
rect 25372 29668 26332 29696
rect 25372 29656 25378 29668
rect 26326 29656 26332 29668
rect 26384 29656 26390 29708
rect 28534 29656 28540 29708
rect 28592 29696 28598 29708
rect 29641 29699 29699 29705
rect 29641 29696 29653 29699
rect 28592 29668 29653 29696
rect 28592 29656 28598 29668
rect 29641 29665 29653 29668
rect 29687 29665 29699 29699
rect 29641 29659 29699 29665
rect 25133 29631 25191 29637
rect 25133 29628 25145 29631
rect 25004 29600 25145 29628
rect 25004 29588 25010 29600
rect 25133 29597 25145 29600
rect 25179 29597 25191 29631
rect 29822 29628 29828 29640
rect 25133 29591 25191 29597
rect 25240 29600 29684 29628
rect 29783 29600 29828 29628
rect 23382 29560 23388 29572
rect 21784 29532 23388 29560
rect 21784 29520 21790 29532
rect 23382 29520 23388 29532
rect 23440 29520 23446 29572
rect 23934 29520 23940 29572
rect 23992 29560 23998 29572
rect 25240 29560 25268 29600
rect 23992 29532 25268 29560
rect 23992 29520 23998 29532
rect 28442 29520 28448 29572
rect 28500 29560 28506 29572
rect 28629 29563 28687 29569
rect 28629 29560 28641 29563
rect 28500 29532 28641 29560
rect 28500 29520 28506 29532
rect 28629 29529 28641 29532
rect 28675 29560 28687 29563
rect 28718 29560 28724 29572
rect 28675 29532 28724 29560
rect 28675 29529 28687 29532
rect 28629 29523 28687 29529
rect 28718 29520 28724 29532
rect 28776 29520 28782 29572
rect 28810 29520 28816 29572
rect 28868 29560 28874 29572
rect 29549 29563 29607 29569
rect 29549 29560 29561 29563
rect 28868 29532 29561 29560
rect 28868 29520 28874 29532
rect 29549 29529 29561 29532
rect 29595 29529 29607 29563
rect 29656 29560 29684 29600
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 29914 29588 29920 29640
rect 29972 29628 29978 29640
rect 30653 29631 30711 29637
rect 30653 29628 30665 29631
rect 29972 29600 30665 29628
rect 29972 29588 29978 29600
rect 30653 29597 30665 29600
rect 30699 29597 30711 29631
rect 30834 29628 30840 29640
rect 30795 29600 30840 29628
rect 30653 29591 30711 29597
rect 30834 29588 30840 29600
rect 30892 29588 30898 29640
rect 30926 29588 30932 29640
rect 30984 29628 30990 29640
rect 30984 29600 31029 29628
rect 30984 29588 30990 29600
rect 32950 29588 32956 29640
rect 33008 29628 33014 29640
rect 33045 29631 33103 29637
rect 33045 29628 33057 29631
rect 33008 29600 33057 29628
rect 33008 29588 33014 29600
rect 33045 29597 33057 29600
rect 33091 29628 33103 29631
rect 46842 29628 46848 29640
rect 33091 29600 46848 29628
rect 33091 29597 33103 29600
rect 33045 29591 33103 29597
rect 46842 29588 46848 29600
rect 46900 29588 46906 29640
rect 48130 29628 48136 29640
rect 48091 29600 48136 29628
rect 48130 29588 48136 29600
rect 48188 29588 48194 29640
rect 32766 29560 32772 29572
rect 29656 29532 32772 29560
rect 29549 29523 29607 29529
rect 32766 29520 32772 29532
rect 32824 29520 32830 29572
rect 21637 29495 21695 29501
rect 21637 29461 21649 29495
rect 21683 29461 21695 29495
rect 21637 29455 21695 29461
rect 23290 29452 23296 29504
rect 23348 29492 23354 29504
rect 25317 29495 25375 29501
rect 25317 29492 25329 29495
rect 23348 29464 25329 29492
rect 23348 29452 23354 29464
rect 25317 29461 25329 29464
rect 25363 29492 25375 29495
rect 26050 29492 26056 29504
rect 25363 29464 26056 29492
rect 25363 29461 25375 29464
rect 25317 29455 25375 29461
rect 26050 29452 26056 29464
rect 26108 29452 26114 29504
rect 30466 29492 30472 29504
rect 30427 29464 30472 29492
rect 30466 29452 30472 29464
rect 30524 29452 30530 29504
rect 47026 29452 47032 29504
rect 47084 29492 47090 29504
rect 47949 29495 48007 29501
rect 47949 29492 47961 29495
rect 47084 29464 47961 29492
rect 47084 29452 47090 29464
rect 47949 29461 47961 29464
rect 47995 29461 48007 29495
rect 47949 29455 48007 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 3326 29248 3332 29300
rect 3384 29288 3390 29300
rect 25314 29288 25320 29300
rect 3384 29260 25320 29288
rect 3384 29248 3390 29260
rect 25314 29248 25320 29260
rect 25372 29248 25378 29300
rect 25961 29291 26019 29297
rect 25961 29257 25973 29291
rect 26007 29288 26019 29291
rect 26050 29288 26056 29300
rect 26007 29260 26056 29288
rect 26007 29257 26019 29260
rect 25961 29251 26019 29257
rect 26050 29248 26056 29260
rect 26108 29248 26114 29300
rect 26878 29248 26884 29300
rect 26936 29288 26942 29300
rect 27341 29291 27399 29297
rect 27341 29288 27353 29291
rect 26936 29260 27353 29288
rect 26936 29248 26942 29260
rect 27341 29257 27353 29260
rect 27387 29257 27399 29291
rect 27341 29251 27399 29257
rect 29825 29291 29883 29297
rect 29825 29257 29837 29291
rect 29871 29288 29883 29291
rect 29914 29288 29920 29300
rect 29871 29260 29920 29288
rect 29871 29257 29883 29260
rect 29825 29251 29883 29257
rect 29914 29248 29920 29260
rect 29972 29248 29978 29300
rect 30006 29248 30012 29300
rect 30064 29248 30070 29300
rect 30282 29288 30288 29300
rect 30243 29260 30288 29288
rect 30282 29248 30288 29260
rect 30340 29248 30346 29300
rect 1670 29180 1676 29232
rect 1728 29220 1734 29232
rect 14458 29220 14464 29232
rect 1728 29192 14464 29220
rect 1728 29180 1734 29192
rect 14458 29180 14464 29192
rect 14516 29180 14522 29232
rect 17589 29223 17647 29229
rect 17589 29189 17601 29223
rect 17635 29220 17647 29223
rect 17635 29192 18092 29220
rect 17635 29189 17647 29192
rect 17589 29183 17647 29189
rect 17310 29152 17316 29164
rect 17271 29124 17316 29152
rect 17310 29112 17316 29124
rect 17368 29112 17374 29164
rect 17402 29112 17408 29164
rect 17460 29152 17466 29164
rect 17678 29155 17736 29161
rect 17460 29124 17505 29152
rect 17460 29112 17466 29124
rect 17678 29121 17690 29155
rect 17724 29121 17736 29155
rect 17678 29115 17736 29121
rect 17817 29155 17875 29161
rect 17817 29121 17829 29155
rect 17863 29152 17875 29155
rect 18064 29152 18092 29192
rect 18138 29180 18144 29232
rect 18196 29220 18202 29232
rect 28810 29220 28816 29232
rect 18196 29192 24072 29220
rect 18196 29180 18202 29192
rect 19978 29152 19984 29164
rect 17863 29124 18000 29152
rect 18064 29124 19840 29152
rect 19939 29124 19984 29152
rect 17863 29121 17875 29124
rect 17817 29115 17875 29121
rect 17218 29044 17224 29096
rect 17276 29084 17282 29096
rect 17696 29084 17724 29115
rect 17276 29056 17724 29084
rect 17276 29044 17282 29056
rect 16298 28976 16304 29028
rect 16356 29016 16362 29028
rect 17972 29016 18000 29124
rect 19812 29084 19840 29124
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 20165 29155 20223 29161
rect 20165 29121 20177 29155
rect 20211 29152 20223 29155
rect 20254 29152 20260 29164
rect 20211 29124 20260 29152
rect 20211 29121 20223 29124
rect 20165 29115 20223 29121
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 20346 29112 20352 29164
rect 20404 29152 20410 29164
rect 20404 29124 20449 29152
rect 20404 29112 20410 29124
rect 21910 29112 21916 29164
rect 21968 29152 21974 29164
rect 23934 29152 23940 29164
rect 21968 29124 23940 29152
rect 21968 29112 21974 29124
rect 23934 29112 23940 29124
rect 23992 29112 23998 29164
rect 20438 29084 20444 29096
rect 19812 29056 20444 29084
rect 20438 29044 20444 29056
rect 20496 29084 20502 29096
rect 24044 29084 24072 29192
rect 28368 29192 28816 29220
rect 25774 29152 25780 29164
rect 25735 29124 25780 29152
rect 25774 29112 25780 29124
rect 25832 29112 25838 29164
rect 28368 29161 28396 29192
rect 28810 29180 28816 29192
rect 28868 29180 28874 29232
rect 30024 29220 30052 29248
rect 29472 29192 30052 29220
rect 29472 29164 29500 29192
rect 26053 29155 26111 29161
rect 26053 29121 26065 29155
rect 26099 29121 26111 29155
rect 28353 29155 28411 29161
rect 28353 29152 28365 29155
rect 26053 29115 26111 29121
rect 27632 29124 28365 29152
rect 26068 29084 26096 29115
rect 27632 29096 27660 29124
rect 28353 29121 28365 29124
rect 28399 29121 28411 29155
rect 28534 29152 28540 29164
rect 28495 29124 28540 29152
rect 28353 29115 28411 29121
rect 28534 29112 28540 29124
rect 28592 29112 28598 29164
rect 29273 29155 29331 29161
rect 29273 29121 29285 29155
rect 29319 29121 29331 29155
rect 29454 29152 29460 29164
rect 29415 29124 29460 29152
rect 29273 29115 29331 29121
rect 27430 29084 27436 29096
rect 20496 29056 23336 29084
rect 24044 29056 26096 29084
rect 27391 29056 27436 29084
rect 20496 29044 20502 29056
rect 20530 29016 20536 29028
rect 16356 28988 20536 29016
rect 16356 28976 16362 28988
rect 20530 28976 20536 28988
rect 20588 28976 20594 29028
rect 23308 29016 23336 29056
rect 27430 29044 27436 29056
rect 27488 29044 27494 29096
rect 27614 29044 27620 29096
rect 27672 29084 27678 29096
rect 27672 29056 27765 29084
rect 27672 29044 27678 29056
rect 24486 29016 24492 29028
rect 23308 28988 24492 29016
rect 24486 28976 24492 28988
rect 24544 28976 24550 29028
rect 26970 29016 26976 29028
rect 26931 28988 26976 29016
rect 26970 28976 26976 28988
rect 27028 28976 27034 29028
rect 17954 28948 17960 28960
rect 17915 28920 17960 28948
rect 17954 28908 17960 28920
rect 18012 28908 18018 28960
rect 25590 28948 25596 28960
rect 25551 28920 25596 28948
rect 25590 28908 25596 28920
rect 25648 28908 25654 28960
rect 27798 28908 27804 28960
rect 27856 28948 27862 28960
rect 27982 28948 27988 28960
rect 27856 28920 27988 28948
rect 27856 28908 27862 28920
rect 27982 28908 27988 28920
rect 28040 28908 28046 28960
rect 28166 28908 28172 28960
rect 28224 28948 28230 28960
rect 28445 28951 28503 28957
rect 28445 28948 28457 28951
rect 28224 28920 28457 28948
rect 28224 28908 28230 28920
rect 28445 28917 28457 28920
rect 28491 28917 28503 28951
rect 29288 28948 29316 29115
rect 29454 29112 29460 29124
rect 29512 29112 29518 29164
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 29641 29155 29699 29161
rect 29641 29121 29653 29155
rect 29687 29152 29699 29155
rect 30006 29152 30012 29164
rect 29687 29124 30012 29152
rect 29687 29121 29699 29124
rect 29641 29115 29699 29121
rect 29362 29044 29368 29096
rect 29420 29084 29426 29096
rect 29564 29084 29592 29115
rect 30006 29112 30012 29124
rect 30064 29112 30070 29164
rect 30469 29155 30527 29161
rect 30469 29121 30481 29155
rect 30515 29152 30527 29155
rect 31754 29152 31760 29164
rect 30515 29124 31760 29152
rect 30515 29121 30527 29124
rect 30469 29115 30527 29121
rect 29420 29056 29592 29084
rect 29420 29044 29426 29056
rect 29822 29044 29828 29096
rect 29880 29084 29886 29096
rect 30484 29084 30512 29115
rect 31754 29112 31760 29124
rect 31812 29112 31818 29164
rect 29880 29056 30512 29084
rect 30745 29087 30803 29093
rect 29880 29044 29886 29056
rect 30745 29053 30757 29087
rect 30791 29084 30803 29087
rect 31294 29084 31300 29096
rect 30791 29056 31300 29084
rect 30791 29053 30803 29056
rect 30745 29047 30803 29053
rect 30282 28976 30288 29028
rect 30340 29016 30346 29028
rect 30653 29019 30711 29025
rect 30653 29016 30665 29019
rect 30340 28988 30665 29016
rect 30340 28976 30346 28988
rect 30653 28985 30665 28988
rect 30699 28985 30711 29019
rect 30653 28979 30711 28985
rect 30374 28948 30380 28960
rect 29288 28920 30380 28948
rect 28445 28911 28503 28917
rect 30374 28908 30380 28920
rect 30432 28948 30438 28960
rect 30760 28948 30788 29047
rect 31294 29044 31300 29056
rect 31352 29044 31358 29096
rect 32306 29084 32312 29096
rect 32267 29056 32312 29084
rect 32306 29044 32312 29056
rect 32364 29044 32370 29096
rect 32490 29084 32496 29096
rect 32451 29056 32496 29084
rect 32490 29044 32496 29056
rect 32548 29044 32554 29096
rect 32766 29084 32772 29096
rect 32727 29056 32772 29084
rect 32766 29044 32772 29056
rect 32824 29044 32830 29096
rect 30432 28920 30788 28948
rect 30432 28908 30438 28920
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 17494 28744 17500 28756
rect 17455 28716 17500 28744
rect 17494 28704 17500 28716
rect 17552 28704 17558 28756
rect 19794 28744 19800 28756
rect 17604 28716 19800 28744
rect 7466 28636 7472 28688
rect 7524 28676 7530 28688
rect 17604 28676 17632 28716
rect 19794 28704 19800 28716
rect 19852 28704 19858 28756
rect 25958 28744 25964 28756
rect 25919 28716 25964 28744
rect 25958 28704 25964 28716
rect 26016 28704 26022 28756
rect 27341 28747 27399 28753
rect 27341 28713 27353 28747
rect 27387 28744 27399 28747
rect 28994 28744 29000 28756
rect 27387 28716 28856 28744
rect 28907 28716 29000 28744
rect 27387 28713 27399 28716
rect 27341 28707 27399 28713
rect 7524 28648 17632 28676
rect 7524 28636 7530 28648
rect 19426 28636 19432 28688
rect 19484 28636 19490 28688
rect 19518 28636 19524 28688
rect 19576 28676 19582 28688
rect 21726 28676 21732 28688
rect 19576 28648 21732 28676
rect 19576 28636 19582 28648
rect 21726 28636 21732 28648
rect 21784 28636 21790 28688
rect 27893 28679 27951 28685
rect 27893 28645 27905 28679
rect 27939 28676 27951 28679
rect 28626 28676 28632 28688
rect 27939 28648 28632 28676
rect 27939 28645 27951 28648
rect 27893 28639 27951 28645
rect 28626 28636 28632 28648
rect 28684 28636 28690 28688
rect 28828 28676 28856 28716
rect 28994 28704 29000 28716
rect 29052 28744 29058 28756
rect 30282 28744 30288 28756
rect 29052 28716 30288 28744
rect 29052 28704 29058 28716
rect 30282 28704 30288 28716
rect 30340 28704 30346 28756
rect 31294 28744 31300 28756
rect 31255 28716 31300 28744
rect 31294 28704 31300 28716
rect 31352 28704 31358 28756
rect 32490 28744 32496 28756
rect 32451 28716 32496 28744
rect 32490 28704 32496 28716
rect 32548 28704 32554 28756
rect 29454 28676 29460 28688
rect 28828 28648 29460 28676
rect 29454 28636 29460 28648
rect 29512 28636 29518 28688
rect 17313 28611 17371 28617
rect 17313 28577 17325 28611
rect 17359 28608 17371 28611
rect 19150 28608 19156 28620
rect 17359 28580 19156 28608
rect 17359 28577 17371 28580
rect 17313 28571 17371 28577
rect 19150 28568 19156 28580
rect 19208 28568 19214 28620
rect 15013 28543 15071 28549
rect 15013 28509 15025 28543
rect 15059 28540 15071 28543
rect 15657 28543 15715 28549
rect 15657 28540 15669 28543
rect 15059 28512 15669 28540
rect 15059 28509 15071 28512
rect 15013 28503 15071 28509
rect 15657 28509 15669 28512
rect 15703 28509 15715 28543
rect 17218 28540 17224 28552
rect 17179 28512 17224 28540
rect 15657 28503 15715 28509
rect 15672 28472 15700 28503
rect 17218 28500 17224 28512
rect 17276 28500 17282 28552
rect 19337 28543 19395 28549
rect 19337 28509 19349 28543
rect 19383 28540 19395 28543
rect 19444 28540 19472 28636
rect 19524 28551 19552 28636
rect 19613 28611 19671 28617
rect 19613 28577 19625 28611
rect 19659 28577 19671 28611
rect 19613 28571 19671 28577
rect 19705 28611 19763 28617
rect 19705 28577 19717 28611
rect 19751 28608 19763 28611
rect 19794 28608 19800 28620
rect 19751 28580 19800 28608
rect 19751 28577 19763 28580
rect 19705 28571 19763 28577
rect 19383 28512 19472 28540
rect 19509 28545 19567 28551
rect 19383 28509 19395 28512
rect 19337 28503 19395 28509
rect 19509 28511 19521 28545
rect 19555 28511 19567 28545
rect 19628 28542 19656 28571
rect 19794 28568 19800 28580
rect 19852 28568 19858 28620
rect 20162 28568 20168 28620
rect 20220 28608 20226 28620
rect 22094 28608 22100 28620
rect 20220 28580 22100 28608
rect 20220 28568 20226 28580
rect 22094 28568 22100 28580
rect 22152 28568 22158 28620
rect 27982 28568 27988 28620
rect 28040 28608 28046 28620
rect 29546 28608 29552 28620
rect 28040 28580 29552 28608
rect 28040 28568 28046 28580
rect 29546 28568 29552 28580
rect 29604 28568 29610 28620
rect 29825 28611 29883 28617
rect 29825 28577 29837 28611
rect 29871 28608 29883 28611
rect 30466 28608 30472 28620
rect 29871 28580 30472 28608
rect 29871 28577 29883 28580
rect 29825 28571 29883 28577
rect 30466 28568 30472 28580
rect 30524 28568 30530 28620
rect 19889 28543 19947 28549
rect 19628 28540 19748 28542
rect 19628 28514 19840 28540
rect 19720 28512 19840 28514
rect 19509 28505 19567 28511
rect 18230 28472 18236 28484
rect 15672 28444 18236 28472
rect 18230 28432 18236 28444
rect 18288 28432 18294 28484
rect 19812 28472 19840 28512
rect 19889 28509 19901 28543
rect 19935 28540 19947 28543
rect 22646 28540 22652 28552
rect 19935 28512 22652 28540
rect 19935 28509 19947 28512
rect 19889 28503 19947 28509
rect 22646 28500 22652 28512
rect 22704 28500 22710 28552
rect 24857 28543 24915 28549
rect 24857 28509 24869 28543
rect 24903 28540 24915 28543
rect 25038 28540 25044 28552
rect 24903 28512 25044 28540
rect 24903 28509 24915 28512
rect 24857 28503 24915 28509
rect 25038 28500 25044 28512
rect 25096 28500 25102 28552
rect 25869 28543 25927 28549
rect 25869 28509 25881 28543
rect 25915 28540 25927 28543
rect 26234 28540 26240 28552
rect 25915 28512 26240 28540
rect 25915 28509 25927 28512
rect 25869 28503 25927 28509
rect 26234 28500 26240 28512
rect 26292 28540 26298 28552
rect 27157 28543 27215 28549
rect 27157 28540 27169 28543
rect 26292 28512 27169 28540
rect 26292 28500 26298 28512
rect 27157 28509 27169 28512
rect 27203 28540 27215 28543
rect 27430 28540 27436 28552
rect 27203 28512 27436 28540
rect 27203 28509 27215 28512
rect 27157 28503 27215 28509
rect 27430 28500 27436 28512
rect 27488 28500 27494 28552
rect 27798 28500 27804 28552
rect 27856 28540 27862 28552
rect 27893 28543 27951 28549
rect 27893 28540 27905 28543
rect 27856 28512 27905 28540
rect 27856 28500 27862 28512
rect 27893 28509 27905 28512
rect 27939 28509 27951 28543
rect 28166 28540 28172 28552
rect 28127 28512 28172 28540
rect 27893 28503 27951 28509
rect 28166 28500 28172 28512
rect 28224 28500 28230 28552
rect 28629 28543 28687 28549
rect 28629 28509 28641 28543
rect 28675 28540 28687 28543
rect 28718 28540 28724 28552
rect 28675 28512 28724 28540
rect 28675 28509 28687 28512
rect 28629 28503 28687 28509
rect 28718 28500 28724 28512
rect 28776 28500 28782 28552
rect 32214 28500 32220 28552
rect 32272 28540 32278 28552
rect 32401 28543 32459 28549
rect 32401 28540 32413 28543
rect 32272 28512 32413 28540
rect 32272 28500 32278 28512
rect 32401 28509 32413 28512
rect 32447 28509 32459 28543
rect 32401 28503 32459 28509
rect 46934 28500 46940 28552
rect 46992 28540 46998 28552
rect 47673 28543 47731 28549
rect 47673 28540 47685 28543
rect 46992 28512 47685 28540
rect 46992 28500 46998 28512
rect 47673 28509 47685 28512
rect 47719 28509 47731 28543
rect 47673 28503 47731 28509
rect 19978 28472 19984 28484
rect 19812 28444 19984 28472
rect 19978 28432 19984 28444
rect 20036 28432 20042 28484
rect 28258 28432 28264 28484
rect 28316 28472 28322 28484
rect 28534 28472 28540 28484
rect 28316 28444 28540 28472
rect 28316 28432 28322 28444
rect 28534 28432 28540 28444
rect 28592 28472 28598 28484
rect 28813 28475 28871 28481
rect 28813 28472 28825 28475
rect 28592 28444 28825 28472
rect 28592 28432 28598 28444
rect 28813 28441 28825 28444
rect 28859 28441 28871 28475
rect 28813 28435 28871 28441
rect 30374 28432 30380 28484
rect 30432 28432 30438 28484
rect 14458 28364 14464 28416
rect 14516 28404 14522 28416
rect 15105 28407 15163 28413
rect 15105 28404 15117 28407
rect 14516 28376 15117 28404
rect 14516 28364 14522 28376
rect 15105 28373 15117 28376
rect 15151 28373 15163 28407
rect 15746 28404 15752 28416
rect 15707 28376 15752 28404
rect 15105 28367 15163 28373
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 19334 28364 19340 28416
rect 19392 28404 19398 28416
rect 20073 28407 20131 28413
rect 20073 28404 20085 28407
rect 19392 28376 20085 28404
rect 19392 28364 19398 28376
rect 20073 28373 20085 28376
rect 20119 28373 20131 28407
rect 20073 28367 20131 28373
rect 24118 28364 24124 28416
rect 24176 28404 24182 28416
rect 24302 28404 24308 28416
rect 24176 28376 24308 28404
rect 24176 28364 24182 28376
rect 24302 28364 24308 28376
rect 24360 28404 24366 28416
rect 24949 28407 25007 28413
rect 24949 28404 24961 28407
rect 24360 28376 24961 28404
rect 24360 28364 24366 28376
rect 24949 28373 24961 28376
rect 24995 28373 25007 28407
rect 24949 28367 25007 28373
rect 28077 28407 28135 28413
rect 28077 28373 28089 28407
rect 28123 28404 28135 28407
rect 28994 28404 29000 28416
rect 28123 28376 29000 28404
rect 28123 28373 28135 28376
rect 28077 28367 28135 28373
rect 28994 28364 29000 28376
rect 29052 28364 29058 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 17218 28160 17224 28212
rect 17276 28200 17282 28212
rect 18785 28203 18843 28209
rect 18785 28200 18797 28203
rect 17276 28172 18797 28200
rect 17276 28160 17282 28172
rect 18785 28169 18797 28172
rect 18831 28169 18843 28203
rect 18785 28163 18843 28169
rect 14458 28132 14464 28144
rect 14419 28104 14464 28132
rect 14458 28092 14464 28104
rect 14516 28092 14522 28144
rect 18598 28132 18604 28144
rect 18538 28104 18604 28132
rect 18598 28092 18604 28104
rect 18656 28092 18662 28144
rect 12710 27956 12716 28008
rect 12768 27996 12774 28008
rect 14277 27999 14335 28005
rect 14277 27996 14289 27999
rect 12768 27968 14289 27996
rect 12768 27956 12774 27968
rect 14277 27965 14289 27968
rect 14323 27965 14335 27999
rect 15838 27996 15844 28008
rect 15799 27968 15844 27996
rect 14277 27959 14335 27965
rect 15838 27956 15844 27968
rect 15896 27956 15902 28008
rect 17034 27996 17040 28008
rect 16995 27968 17040 27996
rect 17034 27956 17040 27968
rect 17092 27956 17098 28008
rect 17313 27999 17371 28005
rect 17313 27965 17325 27999
rect 17359 27996 17371 27999
rect 17954 27996 17960 28008
rect 17359 27968 17960 27996
rect 17359 27965 17371 27968
rect 17313 27959 17371 27965
rect 17954 27956 17960 27968
rect 18012 27956 18018 28008
rect 18800 27996 18828 28163
rect 21174 28160 21180 28212
rect 21232 28200 21238 28212
rect 25869 28203 25927 28209
rect 21232 28172 21956 28200
rect 21232 28160 21238 28172
rect 19978 28132 19984 28144
rect 19444 28104 19984 28132
rect 19444 28073 19472 28104
rect 19978 28092 19984 28104
rect 20036 28132 20042 28144
rect 20533 28135 20591 28141
rect 20036 28104 20392 28132
rect 20036 28092 20042 28104
rect 20364 28073 20392 28104
rect 20533 28101 20545 28135
rect 20579 28132 20591 28135
rect 20579 28104 21036 28132
rect 20579 28101 20591 28104
rect 20533 28095 20591 28101
rect 21008 28076 21036 28104
rect 21450 28092 21456 28144
rect 21508 28132 21514 28144
rect 21821 28135 21879 28141
rect 21821 28132 21833 28135
rect 21508 28104 21833 28132
rect 21508 28092 21514 28104
rect 21821 28101 21833 28104
rect 21867 28101 21879 28135
rect 21928 28132 21956 28172
rect 25869 28169 25881 28203
rect 25915 28200 25927 28203
rect 26234 28200 26240 28212
rect 25915 28172 26240 28200
rect 25915 28169 25927 28172
rect 25869 28163 25927 28169
rect 26234 28160 26240 28172
rect 26292 28160 26298 28212
rect 30561 28203 30619 28209
rect 30561 28169 30573 28203
rect 30607 28200 30619 28203
rect 30926 28200 30932 28212
rect 30607 28172 30932 28200
rect 30607 28169 30619 28172
rect 30561 28163 30619 28169
rect 30926 28160 30932 28172
rect 30984 28160 30990 28212
rect 34514 28160 34520 28212
rect 34572 28200 34578 28212
rect 35621 28203 35679 28209
rect 35621 28200 35633 28203
rect 34572 28172 35633 28200
rect 34572 28160 34578 28172
rect 35621 28169 35633 28172
rect 35667 28169 35679 28203
rect 35621 28163 35679 28169
rect 22005 28135 22063 28141
rect 22005 28132 22017 28135
rect 21928 28104 22017 28132
rect 21821 28095 21879 28101
rect 22005 28101 22017 28104
rect 22051 28101 22063 28135
rect 22005 28095 22063 28101
rect 22186 28092 22192 28144
rect 22244 28132 22250 28144
rect 28626 28132 28632 28144
rect 22244 28104 24256 28132
rect 28587 28104 28632 28132
rect 22244 28092 22250 28104
rect 19429 28067 19487 28073
rect 19429 28033 19441 28067
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 20165 28067 20223 28073
rect 20165 28033 20177 28067
rect 20211 28033 20223 28067
rect 20165 28027 20223 28033
rect 20349 28067 20407 28073
rect 20349 28033 20361 28067
rect 20395 28064 20407 28067
rect 20714 28064 20720 28076
rect 20395 28036 20720 28064
rect 20395 28033 20407 28036
rect 20349 28027 20407 28033
rect 19705 27999 19763 28005
rect 19705 27996 19717 27999
rect 18800 27968 19717 27996
rect 19705 27965 19717 27968
rect 19751 27996 19763 27999
rect 20180 27996 20208 28027
rect 20714 28024 20720 28036
rect 20772 28024 20778 28076
rect 20990 28064 20996 28076
rect 20903 28036 20996 28064
rect 20990 28024 20996 28036
rect 21048 28024 21054 28076
rect 21082 28024 21088 28076
rect 21140 28064 21146 28076
rect 23382 28073 23388 28076
rect 21177 28067 21235 28073
rect 21177 28064 21189 28067
rect 21140 28036 21189 28064
rect 21140 28024 21146 28036
rect 21177 28033 21189 28036
rect 21223 28033 21235 28067
rect 21177 28027 21235 28033
rect 23339 28067 23388 28073
rect 23339 28033 23351 28067
rect 23385 28033 23388 28067
rect 23339 28027 23388 28033
rect 19751 27968 20208 27996
rect 19751 27965 19763 27968
rect 19705 27959 19763 27965
rect 19150 27888 19156 27940
rect 19208 27928 19214 27940
rect 19613 27931 19671 27937
rect 19613 27928 19625 27931
rect 19208 27900 19625 27928
rect 19208 27888 19214 27900
rect 19613 27897 19625 27900
rect 19659 27928 19671 27931
rect 21192 27928 21220 28027
rect 23382 28024 23388 28027
rect 23440 28024 23446 28076
rect 23492 28073 23520 28104
rect 23474 28067 23532 28073
rect 23474 28033 23486 28067
rect 23520 28033 23532 28067
rect 23474 28027 23532 28033
rect 23569 28070 23627 28076
rect 23569 28036 23581 28070
rect 23615 28036 23627 28070
rect 23569 28030 23627 28036
rect 23584 27996 23612 28030
rect 23658 28024 23664 28076
rect 23716 28064 23722 28076
rect 24228 28073 24256 28104
rect 28626 28092 28632 28104
rect 28684 28092 28690 28144
rect 34790 28092 34796 28144
rect 34848 28092 34854 28144
rect 23753 28067 23811 28073
rect 23753 28064 23765 28067
rect 23716 28036 23765 28064
rect 23716 28024 23722 28036
rect 23753 28033 23765 28036
rect 23799 28033 23811 28067
rect 23753 28027 23811 28033
rect 24213 28067 24271 28073
rect 24213 28033 24225 28067
rect 24259 28033 24271 28067
rect 24213 28027 24271 28033
rect 23768 27996 23796 28027
rect 24670 28024 24676 28076
rect 24728 28064 24734 28076
rect 25409 28067 25467 28073
rect 25409 28064 25421 28067
rect 24728 28036 25421 28064
rect 24728 28024 24734 28036
rect 25409 28033 25421 28036
rect 25455 28033 25467 28067
rect 25409 28027 25467 28033
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 27433 28067 27491 28073
rect 27433 28033 27445 28067
rect 27479 28064 27491 28067
rect 27522 28064 27528 28076
rect 27479 28036 27528 28064
rect 27479 28033 27491 28036
rect 27433 28027 27491 28033
rect 24305 27999 24363 28005
rect 24305 27996 24317 27999
rect 23584 27968 23704 27996
rect 23768 27968 24317 27996
rect 22002 27928 22008 27940
rect 19659 27900 22008 27928
rect 19659 27897 19671 27900
rect 19613 27891 19671 27897
rect 22002 27888 22008 27900
rect 22060 27928 22066 27940
rect 22189 27931 22247 27937
rect 22189 27928 22201 27931
rect 22060 27900 22201 27928
rect 22060 27888 22066 27900
rect 22189 27897 22201 27900
rect 22235 27897 22247 27931
rect 23676 27928 23704 27968
rect 24305 27965 24317 27968
rect 24351 27996 24363 27999
rect 24394 27996 24400 28008
rect 24351 27968 24400 27996
rect 24351 27965 24363 27968
rect 24305 27959 24363 27965
rect 24394 27956 24400 27968
rect 24452 27956 24458 28008
rect 25130 27956 25136 28008
rect 25188 27996 25194 28008
rect 25314 27996 25320 28008
rect 25188 27968 25320 27996
rect 25188 27956 25194 27968
rect 25314 27956 25320 27968
rect 25372 27996 25378 28008
rect 25608 27996 25636 28027
rect 27522 28024 27528 28036
rect 27580 28024 27586 28076
rect 28442 28064 28448 28076
rect 28403 28036 28448 28064
rect 28442 28024 28448 28036
rect 28500 28024 28506 28076
rect 30193 28067 30251 28073
rect 30193 28033 30205 28067
rect 30239 28064 30251 28067
rect 31294 28064 31300 28076
rect 30239 28036 31300 28064
rect 30239 28033 30251 28036
rect 30193 28027 30251 28033
rect 31294 28024 31300 28036
rect 31352 28024 31358 28076
rect 45462 28024 45468 28076
rect 45520 28064 45526 28076
rect 47302 28064 47308 28076
rect 45520 28036 47308 28064
rect 45520 28024 45526 28036
rect 47302 28024 47308 28036
rect 47360 28064 47366 28076
rect 47581 28067 47639 28073
rect 47581 28064 47593 28067
rect 47360 28036 47593 28064
rect 47360 28024 47366 28036
rect 47581 28033 47593 28036
rect 47627 28033 47639 28067
rect 47581 28027 47639 28033
rect 25372 27968 25636 27996
rect 25961 27999 26019 28005
rect 25372 27956 25378 27968
rect 25961 27965 25973 27999
rect 26007 27996 26019 27999
rect 27617 27999 27675 28005
rect 27617 27996 27629 27999
rect 26007 27968 27629 27996
rect 26007 27965 26019 27968
rect 25961 27959 26019 27965
rect 27617 27965 27629 27968
rect 27663 27996 27675 27999
rect 28534 27996 28540 28008
rect 27663 27968 28540 27996
rect 27663 27965 27675 27968
rect 27617 27959 27675 27965
rect 28534 27956 28540 27968
rect 28592 27956 28598 28008
rect 30282 27996 30288 28008
rect 30243 27968 30288 27996
rect 30282 27956 30288 27968
rect 30340 27956 30346 28008
rect 33134 27956 33140 28008
rect 33192 27996 33198 28008
rect 33873 27999 33931 28005
rect 33873 27996 33885 27999
rect 33192 27968 33885 27996
rect 33192 27956 33198 27968
rect 33873 27965 33885 27968
rect 33919 27965 33931 27999
rect 34146 27996 34152 28008
rect 34107 27968 34152 27996
rect 33873 27959 33931 27965
rect 34146 27956 34152 27968
rect 34204 27956 34210 28008
rect 24118 27928 24124 27940
rect 23676 27900 24124 27928
rect 22189 27891 22247 27897
rect 24118 27888 24124 27900
rect 24176 27888 24182 27940
rect 24854 27928 24860 27940
rect 24228 27900 24860 27928
rect 19245 27863 19303 27869
rect 19245 27829 19257 27863
rect 19291 27860 19303 27863
rect 19426 27860 19432 27872
rect 19291 27832 19432 27860
rect 19291 27829 19303 27832
rect 19245 27823 19303 27829
rect 19426 27820 19432 27832
rect 19484 27820 19490 27872
rect 20993 27863 21051 27869
rect 20993 27829 21005 27863
rect 21039 27860 21051 27863
rect 21082 27860 21088 27872
rect 21039 27832 21088 27860
rect 21039 27829 21051 27832
rect 20993 27823 21051 27829
rect 21082 27820 21088 27832
rect 21140 27820 21146 27872
rect 23106 27860 23112 27872
rect 23067 27832 23112 27860
rect 23106 27820 23112 27832
rect 23164 27820 23170 27872
rect 23382 27820 23388 27872
rect 23440 27860 23446 27872
rect 24228 27869 24256 27900
rect 24854 27888 24860 27900
rect 24912 27888 24918 27940
rect 24213 27863 24271 27869
rect 24213 27860 24225 27863
rect 23440 27832 24225 27860
rect 23440 27820 23446 27832
rect 24213 27829 24225 27832
rect 24259 27829 24271 27863
rect 24213 27823 24271 27829
rect 24302 27820 24308 27872
rect 24360 27860 24366 27872
rect 24581 27863 24639 27869
rect 24581 27860 24593 27863
rect 24360 27832 24593 27860
rect 24360 27820 24366 27832
rect 24581 27829 24593 27832
rect 24627 27829 24639 27863
rect 24581 27823 24639 27829
rect 28534 27820 28540 27872
rect 28592 27860 28598 27872
rect 28813 27863 28871 27869
rect 28813 27860 28825 27863
rect 28592 27832 28825 27860
rect 28592 27820 28598 27832
rect 28813 27829 28825 27832
rect 28859 27829 28871 27863
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 28813 27823 28871 27829
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 3326 27616 3332 27668
rect 3384 27656 3390 27668
rect 19426 27656 19432 27668
rect 3384 27628 15148 27656
rect 19387 27628 19432 27656
rect 3384 27616 3390 27628
rect 15120 27588 15148 27628
rect 19426 27616 19432 27628
rect 19484 27616 19490 27668
rect 19518 27616 19524 27668
rect 19576 27656 19582 27668
rect 19797 27659 19855 27665
rect 19797 27656 19809 27659
rect 19576 27628 19809 27656
rect 19576 27616 19582 27628
rect 19797 27625 19809 27628
rect 19843 27625 19855 27659
rect 19797 27619 19855 27625
rect 20990 27616 20996 27668
rect 21048 27656 21054 27668
rect 21269 27659 21327 27665
rect 21269 27656 21281 27659
rect 21048 27628 21281 27656
rect 21048 27616 21054 27628
rect 21269 27625 21281 27628
rect 21315 27625 21327 27659
rect 21269 27619 21327 27625
rect 21361 27659 21419 27665
rect 21361 27625 21373 27659
rect 21407 27656 21419 27659
rect 21450 27656 21456 27668
rect 21407 27628 21456 27656
rect 21407 27625 21419 27628
rect 21361 27619 21419 27625
rect 21450 27616 21456 27628
rect 21508 27656 21514 27668
rect 22005 27659 22063 27665
rect 22005 27656 22017 27659
rect 21508 27628 22017 27656
rect 21508 27616 21514 27628
rect 22005 27625 22017 27628
rect 22051 27625 22063 27659
rect 22005 27619 22063 27625
rect 23106 27616 23112 27668
rect 23164 27656 23170 27668
rect 23658 27656 23664 27668
rect 23164 27628 23664 27656
rect 23164 27616 23170 27628
rect 23658 27616 23664 27628
rect 23716 27616 23722 27668
rect 25590 27616 25596 27668
rect 25648 27656 25654 27668
rect 26126 27659 26184 27665
rect 26126 27656 26138 27659
rect 25648 27628 26138 27656
rect 25648 27616 25654 27628
rect 26126 27625 26138 27628
rect 26172 27625 26184 27659
rect 27614 27656 27620 27668
rect 27575 27628 27620 27656
rect 26126 27619 26184 27625
rect 27614 27616 27620 27628
rect 27672 27616 27678 27668
rect 28442 27616 28448 27668
rect 28500 27656 28506 27668
rect 28721 27659 28779 27665
rect 28721 27656 28733 27659
rect 28500 27628 28733 27656
rect 28500 27616 28506 27628
rect 28721 27625 28733 27628
rect 28767 27625 28779 27659
rect 34146 27656 34152 27668
rect 34107 27628 34152 27656
rect 28721 27619 28779 27625
rect 34146 27616 34152 27628
rect 34204 27616 34210 27668
rect 43714 27616 43720 27668
rect 43772 27656 43778 27668
rect 45554 27656 45560 27668
rect 43772 27628 45560 27656
rect 43772 27616 43778 27628
rect 45554 27616 45560 27628
rect 45612 27616 45618 27668
rect 18598 27588 18604 27600
rect 15120 27560 15884 27588
rect 18559 27560 18604 27588
rect 15105 27523 15163 27529
rect 15105 27489 15117 27523
rect 15151 27520 15163 27523
rect 15746 27520 15752 27532
rect 15151 27492 15752 27520
rect 15151 27489 15163 27492
rect 15105 27483 15163 27489
rect 15746 27480 15752 27492
rect 15804 27480 15810 27532
rect 15856 27529 15884 27560
rect 18598 27548 18604 27560
rect 18656 27548 18662 27600
rect 21082 27588 21088 27600
rect 20916 27560 21088 27588
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27489 15899 27523
rect 20162 27520 20168 27532
rect 15841 27483 15899 27489
rect 19444 27492 20168 27520
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 18509 27455 18567 27461
rect 18509 27421 18521 27455
rect 18555 27452 18567 27455
rect 18690 27452 18696 27464
rect 18555 27424 18696 27452
rect 18555 27421 18567 27424
rect 18509 27415 18567 27421
rect 14936 27384 14964 27415
rect 18690 27412 18696 27424
rect 18748 27412 18754 27464
rect 19444 27461 19472 27492
rect 20162 27480 20168 27492
rect 20220 27480 20226 27532
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27452 19671 27455
rect 20916 27452 20944 27560
rect 21082 27548 21088 27560
rect 21140 27548 21146 27600
rect 23382 27548 23388 27600
rect 23440 27588 23446 27600
rect 25314 27588 25320 27600
rect 23440 27560 25320 27588
rect 23440 27548 23446 27560
rect 25314 27548 25320 27560
rect 25372 27548 25378 27600
rect 29825 27591 29883 27597
rect 29825 27557 29837 27591
rect 29871 27588 29883 27591
rect 30374 27588 30380 27600
rect 29871 27560 30380 27588
rect 29871 27557 29883 27560
rect 29825 27551 29883 27557
rect 30374 27548 30380 27560
rect 30432 27548 30438 27600
rect 33045 27591 33103 27597
rect 33045 27557 33057 27591
rect 33091 27588 33103 27591
rect 33134 27588 33140 27600
rect 33091 27560 33140 27588
rect 33091 27557 33103 27560
rect 33045 27551 33103 27557
rect 33134 27548 33140 27560
rect 33192 27548 33198 27600
rect 34790 27548 34796 27600
rect 34848 27588 34854 27600
rect 35069 27591 35127 27597
rect 35069 27588 35081 27591
rect 34848 27560 35081 27588
rect 34848 27548 34854 27560
rect 35069 27557 35081 27560
rect 35115 27557 35127 27591
rect 46934 27588 46940 27600
rect 35069 27551 35127 27557
rect 46308 27560 46940 27588
rect 20990 27480 20996 27532
rect 21048 27520 21054 27532
rect 21818 27520 21824 27532
rect 21048 27492 21824 27520
rect 21048 27480 21054 27492
rect 21818 27480 21824 27492
rect 21876 27520 21882 27532
rect 22097 27523 22155 27529
rect 22097 27520 22109 27523
rect 21876 27492 22109 27520
rect 21876 27480 21882 27492
rect 22097 27489 22109 27492
rect 22143 27489 22155 27523
rect 22097 27483 22155 27489
rect 23477 27523 23535 27529
rect 23477 27489 23489 27523
rect 23523 27520 23535 27523
rect 23750 27520 23756 27532
rect 23523 27492 23756 27520
rect 23523 27489 23535 27492
rect 23477 27483 23535 27489
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 24026 27480 24032 27532
rect 24084 27520 24090 27532
rect 25869 27523 25927 27529
rect 25869 27520 25881 27523
rect 24084 27492 25881 27520
rect 24084 27480 24090 27492
rect 25869 27489 25881 27492
rect 25915 27520 25927 27523
rect 27982 27520 27988 27532
rect 25915 27492 27988 27520
rect 25915 27489 25927 27492
rect 25869 27483 25927 27489
rect 27982 27480 27988 27492
rect 28040 27480 28046 27532
rect 33873 27523 33931 27529
rect 33873 27489 33885 27523
rect 33919 27520 33931 27523
rect 34146 27520 34152 27532
rect 33919 27492 34152 27520
rect 33919 27489 33931 27492
rect 33873 27483 33931 27489
rect 34146 27480 34152 27492
rect 34204 27480 34210 27532
rect 46308 27529 46336 27560
rect 46934 27548 46940 27560
rect 46992 27548 46998 27600
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46293 27483 46351 27489
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 47670 27520 47676 27532
rect 46523 27492 47676 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 47670 27480 47676 27492
rect 47728 27480 47734 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 21082 27452 21088 27464
rect 19659 27424 20944 27452
rect 21043 27424 21088 27452
rect 19659 27421 19671 27424
rect 19613 27415 19671 27421
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 21177 27455 21235 27461
rect 21177 27421 21189 27455
rect 21223 27421 21235 27455
rect 21177 27415 21235 27421
rect 17586 27384 17592 27396
rect 14936 27356 17592 27384
rect 17586 27344 17592 27356
rect 17644 27344 17650 27396
rect 21192 27384 21220 27415
rect 21266 27412 21272 27464
rect 21324 27452 21330 27464
rect 21545 27455 21603 27461
rect 21545 27452 21557 27455
rect 21324 27424 21557 27452
rect 21324 27412 21330 27424
rect 21545 27421 21557 27424
rect 21591 27421 21603 27455
rect 21545 27415 21603 27421
rect 21910 27412 21916 27464
rect 21968 27452 21974 27464
rect 22281 27455 22339 27461
rect 22281 27452 22293 27455
rect 21968 27424 22293 27452
rect 21968 27412 21974 27424
rect 22281 27421 22293 27424
rect 22327 27421 22339 27455
rect 23106 27452 23112 27464
rect 23067 27424 23112 27452
rect 22281 27415 22339 27421
rect 23106 27412 23112 27424
rect 23164 27412 23170 27464
rect 24765 27455 24823 27461
rect 24765 27452 24777 27455
rect 23216 27424 24777 27452
rect 22005 27387 22063 27393
rect 22005 27384 22017 27387
rect 21192 27356 22017 27384
rect 22005 27353 22017 27356
rect 22051 27384 22063 27387
rect 23216 27384 23244 27424
rect 24765 27421 24777 27424
rect 24811 27421 24823 27455
rect 24765 27415 24823 27421
rect 27246 27412 27252 27464
rect 27304 27412 27310 27464
rect 28166 27452 28172 27464
rect 28127 27424 28172 27452
rect 28166 27412 28172 27424
rect 28224 27412 28230 27464
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27452 28595 27455
rect 28810 27452 28816 27464
rect 28583 27424 28816 27452
rect 28583 27421 28595 27424
rect 28537 27415 28595 27421
rect 28810 27412 28816 27424
rect 28868 27412 28874 27464
rect 29546 27412 29552 27464
rect 29604 27452 29610 27464
rect 29733 27455 29791 27461
rect 29733 27452 29745 27455
rect 29604 27424 29745 27452
rect 29604 27412 29610 27424
rect 29733 27421 29745 27424
rect 29779 27421 29791 27455
rect 29733 27415 29791 27421
rect 31202 27412 31208 27464
rect 31260 27452 31266 27464
rect 32953 27455 33011 27461
rect 32953 27452 32965 27455
rect 31260 27424 32965 27452
rect 31260 27412 31266 27424
rect 32953 27421 32965 27424
rect 32999 27421 33011 27455
rect 32953 27415 33011 27421
rect 33781 27455 33839 27461
rect 33781 27421 33793 27455
rect 33827 27452 33839 27455
rect 34514 27452 34520 27464
rect 33827 27424 34520 27452
rect 33827 27421 33839 27424
rect 33781 27415 33839 27421
rect 34514 27412 34520 27424
rect 34572 27412 34578 27464
rect 34977 27455 35035 27461
rect 34977 27421 34989 27455
rect 35023 27452 35035 27455
rect 35526 27452 35532 27464
rect 35023 27424 35532 27452
rect 35023 27421 35035 27424
rect 34977 27415 35035 27421
rect 35526 27412 35532 27424
rect 35584 27412 35590 27464
rect 23382 27384 23388 27396
rect 22051 27356 23244 27384
rect 23343 27356 23388 27384
rect 22051 27353 22063 27356
rect 22005 27347 22063 27353
rect 23382 27344 23388 27356
rect 23440 27344 23446 27396
rect 23594 27387 23652 27393
rect 23594 27353 23606 27387
rect 23640 27384 23652 27387
rect 23934 27384 23940 27396
rect 23640 27356 23940 27384
rect 23640 27353 23652 27356
rect 23594 27347 23652 27353
rect 23934 27344 23940 27356
rect 23992 27344 23998 27396
rect 24394 27384 24400 27396
rect 24355 27356 24400 27384
rect 24394 27344 24400 27356
rect 24452 27344 24458 27396
rect 24578 27384 24584 27396
rect 24539 27356 24584 27384
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 27430 27344 27436 27396
rect 27488 27384 27494 27396
rect 28353 27387 28411 27393
rect 28353 27384 28365 27387
rect 27488 27356 28365 27384
rect 27488 27344 27494 27356
rect 28353 27353 28365 27356
rect 28399 27353 28411 27387
rect 28353 27347 28411 27353
rect 28445 27387 28503 27393
rect 28445 27353 28457 27387
rect 28491 27384 28503 27387
rect 28626 27384 28632 27396
rect 28491 27356 28632 27384
rect 28491 27353 28503 27356
rect 28445 27347 28503 27353
rect 28626 27344 28632 27356
rect 28684 27344 28690 27396
rect 20809 27319 20867 27325
rect 20809 27285 20821 27319
rect 20855 27316 20867 27319
rect 21358 27316 21364 27328
rect 20855 27288 21364 27316
rect 20855 27285 20867 27288
rect 20809 27279 20867 27285
rect 21358 27276 21364 27288
rect 21416 27276 21422 27328
rect 22465 27319 22523 27325
rect 22465 27285 22477 27319
rect 22511 27316 22523 27319
rect 23198 27316 23204 27328
rect 22511 27288 23204 27316
rect 22511 27285 22523 27288
rect 22465 27279 22523 27285
rect 23198 27276 23204 27288
rect 23256 27276 23262 27328
rect 23750 27316 23756 27328
rect 23711 27288 23756 27316
rect 23750 27276 23756 27288
rect 23808 27276 23814 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 20714 27112 20720 27124
rect 20675 27084 20720 27112
rect 20714 27072 20720 27084
rect 20772 27072 20778 27124
rect 22186 27112 22192 27124
rect 22147 27084 22192 27112
rect 22186 27072 22192 27084
rect 22244 27072 22250 27124
rect 23934 27112 23940 27124
rect 23032 27084 23940 27112
rect 17034 27004 17040 27056
rect 17092 27044 17098 27056
rect 19245 27047 19303 27053
rect 17092 27016 19012 27044
rect 17092 27004 17098 27016
rect 12253 26979 12311 26985
rect 12253 26945 12265 26979
rect 12299 26976 12311 26979
rect 12299 26948 13768 26976
rect 12299 26945 12311 26948
rect 12253 26939 12311 26945
rect 13740 26920 13768 26948
rect 18984 26920 19012 27016
rect 19245 27013 19257 27047
rect 19291 27044 19303 27047
rect 19334 27044 19340 27056
rect 19291 27016 19340 27044
rect 19291 27013 19303 27016
rect 19245 27007 19303 27013
rect 19334 27004 19340 27016
rect 19392 27004 19398 27056
rect 19978 27004 19984 27056
rect 20036 27004 20042 27056
rect 21818 27044 21824 27056
rect 21779 27016 21824 27044
rect 21818 27004 21824 27016
rect 21876 27004 21882 27056
rect 22002 27044 22008 27056
rect 21963 27016 22008 27044
rect 22002 27004 22008 27016
rect 22060 27004 22066 27056
rect 23032 26985 23060 27084
rect 23934 27072 23940 27084
rect 23992 27072 23998 27124
rect 24578 27072 24584 27124
rect 24636 27112 24642 27124
rect 25777 27115 25835 27121
rect 25777 27112 25789 27115
rect 24636 27084 25789 27112
rect 24636 27072 24642 27084
rect 25777 27081 25789 27084
rect 25823 27081 25835 27115
rect 25777 27075 25835 27081
rect 27246 27072 27252 27124
rect 27304 27112 27310 27124
rect 27341 27115 27399 27121
rect 27341 27112 27353 27115
rect 27304 27084 27353 27112
rect 27304 27072 27310 27084
rect 27341 27081 27353 27084
rect 27387 27081 27399 27115
rect 27341 27075 27399 27081
rect 28166 27072 28172 27124
rect 28224 27112 28230 27124
rect 29733 27115 29791 27121
rect 29733 27112 29745 27115
rect 28224 27084 29745 27112
rect 28224 27072 28230 27084
rect 29733 27081 29745 27084
rect 29779 27081 29791 27115
rect 29733 27075 29791 27081
rect 32306 27072 32312 27124
rect 32364 27112 32370 27124
rect 33873 27115 33931 27121
rect 33873 27112 33885 27115
rect 32364 27084 33885 27112
rect 32364 27072 32370 27084
rect 33873 27081 33885 27084
rect 33919 27081 33931 27115
rect 33873 27075 33931 27081
rect 23201 27047 23259 27053
rect 23201 27013 23213 27047
rect 23247 27044 23259 27047
rect 24302 27044 24308 27056
rect 23247 27016 24308 27044
rect 23247 27013 23259 27016
rect 23201 27007 23259 27013
rect 24302 27004 24308 27016
rect 24360 27004 24366 27056
rect 25314 27004 25320 27056
rect 25372 27004 25378 27056
rect 29638 27044 29644 27056
rect 29486 27016 29644 27044
rect 29638 27004 29644 27016
rect 29696 27004 29702 27056
rect 33134 27004 33140 27056
rect 33192 27004 33198 27056
rect 34238 27004 34244 27056
rect 34296 27044 34302 27056
rect 34517 27047 34575 27053
rect 34517 27044 34529 27047
rect 34296 27016 34529 27044
rect 34296 27004 34302 27016
rect 34517 27013 34529 27016
rect 34563 27013 34575 27047
rect 34517 27007 34575 27013
rect 23017 26979 23075 26985
rect 23017 26945 23029 26979
rect 23063 26945 23075 26979
rect 23290 26976 23296 26988
rect 23251 26948 23296 26976
rect 23017 26939 23075 26945
rect 23290 26936 23296 26948
rect 23348 26936 23354 26988
rect 23385 26979 23443 26985
rect 23385 26945 23397 26979
rect 23431 26945 23443 26979
rect 24026 26976 24032 26988
rect 23987 26948 24032 26976
rect 23385 26939 23443 26945
rect 12342 26908 12348 26920
rect 12303 26880 12348 26908
rect 12342 26868 12348 26880
rect 12400 26868 12406 26920
rect 13722 26868 13728 26920
rect 13780 26908 13786 26920
rect 16669 26911 16727 26917
rect 16669 26908 16681 26911
rect 13780 26880 16681 26908
rect 13780 26868 13786 26880
rect 16669 26877 16681 26880
rect 16715 26877 16727 26911
rect 16850 26908 16856 26920
rect 16811 26880 16856 26908
rect 16669 26871 16727 26877
rect 16850 26868 16856 26880
rect 16908 26868 16914 26920
rect 17126 26908 17132 26920
rect 17087 26880 17132 26908
rect 17126 26868 17132 26880
rect 17184 26868 17190 26920
rect 18966 26908 18972 26920
rect 18927 26880 18972 26908
rect 18966 26868 18972 26880
rect 19024 26868 19030 26920
rect 22646 26868 22652 26920
rect 22704 26908 22710 26920
rect 23400 26908 23428 26939
rect 24026 26936 24032 26948
rect 24084 26936 24090 26988
rect 27249 26979 27307 26985
rect 27249 26945 27261 26979
rect 27295 26976 27307 26979
rect 27614 26976 27620 26988
rect 27295 26948 27620 26976
rect 27295 26945 27307 26948
rect 27249 26939 27307 26945
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 27982 26976 27988 26988
rect 27943 26948 27988 26976
rect 27982 26936 27988 26948
rect 28040 26936 28046 26988
rect 31202 26936 31208 26988
rect 31260 26976 31266 26988
rect 31297 26979 31355 26985
rect 31297 26976 31309 26979
rect 31260 26948 31309 26976
rect 31260 26936 31266 26948
rect 31297 26945 31309 26948
rect 31343 26945 31355 26979
rect 31297 26939 31355 26945
rect 34054 26936 34060 26988
rect 34112 26976 34118 26988
rect 34333 26979 34391 26985
rect 34333 26976 34345 26979
rect 34112 26948 34345 26976
rect 34112 26936 34118 26948
rect 34333 26945 34345 26948
rect 34379 26945 34391 26979
rect 34333 26939 34391 26945
rect 34609 26979 34667 26985
rect 34609 26945 34621 26979
rect 34655 26945 34667 26979
rect 34609 26939 34667 26945
rect 24305 26911 24363 26917
rect 24305 26908 24317 26911
rect 22704 26880 23428 26908
rect 23584 26880 24317 26908
rect 22704 26868 22710 26880
rect 12618 26840 12624 26852
rect 12579 26812 12624 26840
rect 12618 26800 12624 26812
rect 12676 26800 12682 26852
rect 23584 26849 23612 26880
rect 24305 26877 24317 26880
rect 24351 26877 24363 26911
rect 24305 26871 24363 26877
rect 28261 26911 28319 26917
rect 28261 26877 28273 26911
rect 28307 26908 28319 26911
rect 28350 26908 28356 26920
rect 28307 26880 28356 26908
rect 28307 26877 28319 26880
rect 28261 26871 28319 26877
rect 28350 26868 28356 26880
rect 28408 26868 28414 26920
rect 31573 26911 31631 26917
rect 31573 26877 31585 26911
rect 31619 26908 31631 26911
rect 32125 26911 32183 26917
rect 32125 26908 32137 26911
rect 31619 26880 32137 26908
rect 31619 26877 31631 26880
rect 31573 26871 31631 26877
rect 32125 26877 32137 26880
rect 32171 26877 32183 26911
rect 32398 26908 32404 26920
rect 32359 26880 32404 26908
rect 32125 26871 32183 26877
rect 32398 26868 32404 26880
rect 32456 26868 32462 26920
rect 33962 26868 33968 26920
rect 34020 26908 34026 26920
rect 34624 26908 34652 26939
rect 34020 26880 34652 26908
rect 34020 26868 34026 26880
rect 47118 26868 47124 26920
rect 47176 26908 47182 26920
rect 48038 26908 48044 26920
rect 47176 26880 48044 26908
rect 47176 26868 47182 26880
rect 48038 26868 48044 26880
rect 48096 26868 48102 26920
rect 23569 26843 23627 26849
rect 23569 26809 23581 26843
rect 23615 26809 23627 26843
rect 23569 26803 23627 26809
rect 18782 26732 18788 26784
rect 18840 26772 18846 26784
rect 26142 26772 26148 26784
rect 18840 26744 26148 26772
rect 18840 26732 18846 26744
rect 26142 26732 26148 26744
rect 26200 26732 26206 26784
rect 34333 26775 34391 26781
rect 34333 26741 34345 26775
rect 34379 26772 34391 26775
rect 34790 26772 34796 26784
rect 34379 26744 34796 26772
rect 34379 26741 34391 26744
rect 34333 26735 34391 26741
rect 34790 26732 34796 26744
rect 34848 26732 34854 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 12342 26528 12348 26580
rect 12400 26568 12406 26580
rect 12621 26571 12679 26577
rect 12621 26568 12633 26571
rect 12400 26540 12633 26568
rect 12400 26528 12406 26540
rect 12621 26537 12633 26540
rect 12667 26537 12679 26571
rect 12621 26531 12679 26537
rect 15289 26571 15347 26577
rect 15289 26537 15301 26571
rect 15335 26568 15347 26571
rect 16850 26568 16856 26580
rect 15335 26540 16856 26568
rect 15335 26537 15347 26540
rect 15289 26531 15347 26537
rect 16850 26528 16856 26540
rect 16908 26528 16914 26580
rect 19978 26528 19984 26580
rect 20036 26568 20042 26580
rect 20073 26571 20131 26577
rect 20073 26568 20085 26571
rect 20036 26540 20085 26568
rect 20036 26528 20042 26540
rect 20073 26537 20085 26540
rect 20119 26537 20131 26571
rect 20073 26531 20131 26537
rect 23106 26528 23112 26580
rect 23164 26568 23170 26580
rect 23385 26571 23443 26577
rect 23385 26568 23397 26571
rect 23164 26540 23397 26568
rect 23164 26528 23170 26540
rect 23385 26537 23397 26540
rect 23431 26568 23443 26571
rect 23566 26568 23572 26580
rect 23431 26540 23572 26568
rect 23431 26537 23443 26540
rect 23385 26531 23443 26537
rect 23566 26528 23572 26540
rect 23624 26528 23630 26580
rect 23934 26528 23940 26580
rect 23992 26568 23998 26580
rect 24765 26571 24823 26577
rect 24765 26568 24777 26571
rect 23992 26540 24777 26568
rect 23992 26528 23998 26540
rect 24765 26537 24777 26540
rect 24811 26537 24823 26571
rect 25314 26568 25320 26580
rect 25275 26540 25320 26568
rect 24765 26531 24823 26537
rect 25314 26528 25320 26540
rect 25372 26528 25378 26580
rect 28350 26568 28356 26580
rect 28311 26540 28356 26568
rect 28350 26528 28356 26540
rect 28408 26528 28414 26580
rect 29638 26568 29644 26580
rect 29599 26540 29644 26568
rect 29638 26528 29644 26540
rect 29696 26528 29702 26580
rect 32398 26528 32404 26580
rect 32456 26568 32462 26580
rect 32677 26571 32735 26577
rect 32677 26568 32689 26571
rect 32456 26540 32689 26568
rect 32456 26528 32462 26540
rect 32677 26537 32689 26540
rect 32723 26537 32735 26571
rect 34146 26568 34152 26580
rect 34107 26540 34152 26568
rect 32677 26531 32735 26537
rect 34146 26528 34152 26540
rect 34204 26528 34210 26580
rect 18693 26503 18751 26509
rect 18693 26469 18705 26503
rect 18739 26500 18751 26503
rect 18782 26500 18788 26512
rect 18739 26472 18788 26500
rect 18739 26469 18751 26472
rect 18693 26463 18751 26469
rect 18782 26460 18788 26472
rect 18840 26460 18846 26512
rect 24578 26500 24584 26512
rect 24412 26472 24584 26500
rect 8294 26392 8300 26444
rect 8352 26432 8358 26444
rect 16301 26435 16359 26441
rect 16301 26432 16313 26435
rect 8352 26404 16313 26432
rect 8352 26392 8358 26404
rect 16301 26401 16313 26404
rect 16347 26401 16359 26435
rect 16301 26395 16359 26401
rect 18966 26392 18972 26444
rect 19024 26432 19030 26444
rect 21637 26435 21695 26441
rect 21637 26432 21649 26435
rect 19024 26404 21649 26432
rect 19024 26392 19030 26404
rect 21637 26401 21649 26404
rect 21683 26401 21695 26435
rect 21637 26395 21695 26401
rect 21913 26435 21971 26441
rect 21913 26401 21925 26435
rect 21959 26432 21971 26435
rect 23106 26432 23112 26444
rect 21959 26404 23112 26432
rect 21959 26401 21971 26404
rect 21913 26395 21971 26401
rect 23106 26392 23112 26404
rect 23164 26392 23170 26444
rect 24412 26441 24440 26472
rect 24578 26460 24584 26472
rect 24636 26460 24642 26512
rect 27525 26503 27583 26509
rect 27525 26469 27537 26503
rect 27571 26500 27583 26503
rect 27614 26500 27620 26512
rect 27571 26472 27620 26500
rect 27571 26469 27583 26472
rect 27525 26463 27583 26469
rect 27614 26460 27620 26472
rect 27672 26500 27678 26512
rect 29546 26500 29552 26512
rect 27672 26472 29552 26500
rect 27672 26460 27678 26472
rect 29546 26460 29552 26472
rect 29604 26460 29610 26512
rect 24397 26435 24455 26441
rect 24397 26401 24409 26435
rect 24443 26401 24455 26435
rect 31018 26432 31024 26444
rect 30979 26404 31024 26432
rect 24397 26395 24455 26401
rect 31018 26392 31024 26404
rect 31076 26432 31082 26444
rect 31478 26432 31484 26444
rect 31076 26404 31484 26432
rect 31076 26392 31082 26404
rect 31478 26392 31484 26404
rect 31536 26392 31542 26444
rect 32401 26435 32459 26441
rect 32401 26401 32413 26435
rect 32447 26432 32459 26435
rect 34422 26432 34428 26444
rect 32447 26404 34428 26432
rect 32447 26401 32459 26404
rect 32401 26395 32459 26401
rect 34422 26392 34428 26404
rect 34480 26392 34486 26444
rect 39301 26435 39359 26441
rect 34532 26404 36676 26432
rect 11882 26364 11888 26376
rect 11843 26336 11888 26364
rect 11882 26324 11888 26336
rect 11940 26324 11946 26376
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26333 12587 26367
rect 12710 26364 12716 26376
rect 12671 26336 12716 26364
rect 12529 26327 12587 26333
rect 11977 26299 12035 26305
rect 11977 26265 11989 26299
rect 12023 26296 12035 26299
rect 12434 26296 12440 26308
rect 12023 26268 12440 26296
rect 12023 26265 12035 26268
rect 11977 26259 12035 26265
rect 12434 26256 12440 26268
rect 12492 26256 12498 26308
rect 12544 26296 12572 26327
rect 12710 26324 12716 26336
rect 12768 26364 12774 26376
rect 13078 26364 13084 26376
rect 12768 26336 13084 26364
rect 12768 26324 12774 26336
rect 13078 26324 13084 26336
rect 13136 26324 13142 26376
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26364 13231 26367
rect 14093 26367 14151 26373
rect 14093 26364 14105 26367
rect 13219 26336 14105 26364
rect 13219 26333 13231 26336
rect 13173 26327 13231 26333
rect 14093 26333 14105 26336
rect 14139 26364 14151 26367
rect 14826 26364 14832 26376
rect 14139 26336 14832 26364
rect 14139 26333 14151 26336
rect 14093 26327 14151 26333
rect 14826 26324 14832 26336
rect 14884 26324 14890 26376
rect 15197 26367 15255 26373
rect 15197 26333 15209 26367
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 13354 26296 13360 26308
rect 12544 26268 13360 26296
rect 13354 26256 13360 26268
rect 13412 26256 13418 26308
rect 14182 26296 14188 26308
rect 14143 26268 14188 26296
rect 14182 26256 14188 26268
rect 14240 26256 14246 26308
rect 13262 26228 13268 26240
rect 13223 26200 13268 26228
rect 13262 26188 13268 26200
rect 13320 26188 13326 26240
rect 15212 26228 15240 26327
rect 15286 26324 15292 26376
rect 15344 26364 15350 26376
rect 15841 26367 15899 26373
rect 15841 26364 15853 26367
rect 15344 26336 15853 26364
rect 15344 26324 15350 26336
rect 15841 26333 15853 26336
rect 15887 26333 15899 26367
rect 18506 26364 18512 26376
rect 18419 26336 18512 26364
rect 15841 26327 15899 26333
rect 18506 26324 18512 26336
rect 18564 26364 18570 26376
rect 19242 26364 19248 26376
rect 18564 26336 19248 26364
rect 18564 26324 18570 26336
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 19981 26367 20039 26373
rect 19981 26333 19993 26367
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26364 24639 26367
rect 25038 26364 25044 26376
rect 24627 26336 25044 26364
rect 24627 26333 24639 26336
rect 24581 26327 24639 26333
rect 16025 26299 16083 26305
rect 16025 26265 16037 26299
rect 16071 26296 16083 26299
rect 16942 26296 16948 26308
rect 16071 26268 16948 26296
rect 16071 26265 16083 26268
rect 16025 26259 16083 26265
rect 16942 26256 16948 26268
rect 17000 26256 17006 26308
rect 18690 26256 18696 26308
rect 18748 26296 18754 26308
rect 19996 26296 20024 26327
rect 25038 26324 25044 26336
rect 25096 26324 25102 26376
rect 25225 26367 25283 26373
rect 25225 26333 25237 26367
rect 25271 26333 25283 26367
rect 25225 26327 25283 26333
rect 22186 26296 22192 26308
rect 18748 26268 22192 26296
rect 18748 26256 18754 26268
rect 16298 26228 16304 26240
rect 15212 26200 16304 26228
rect 16298 26188 16304 26200
rect 16356 26188 16362 26240
rect 19444 26237 19472 26268
rect 22186 26256 22192 26268
rect 22244 26256 22250 26308
rect 22554 26256 22560 26308
rect 22612 26256 22618 26308
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 25240 26296 25268 26327
rect 26142 26324 26148 26376
rect 26200 26364 26206 26376
rect 27338 26364 27344 26376
rect 26200 26336 27344 26364
rect 26200 26324 26206 26336
rect 27338 26324 27344 26336
rect 27396 26324 27402 26376
rect 28534 26364 28540 26376
rect 28495 26336 28540 26364
rect 28534 26324 28540 26336
rect 28592 26324 28598 26376
rect 29546 26364 29552 26376
rect 29507 26336 29552 26364
rect 29546 26324 29552 26336
rect 29604 26324 29610 26376
rect 30374 26324 30380 26376
rect 30432 26364 30438 26376
rect 30469 26367 30527 26373
rect 30469 26364 30481 26367
rect 30432 26336 30481 26364
rect 30432 26324 30438 26336
rect 30469 26333 30481 26336
rect 30515 26333 30527 26367
rect 32306 26364 32312 26376
rect 32267 26336 32312 26364
rect 30469 26327 30527 26333
rect 32306 26324 32312 26336
rect 32364 26364 32370 26376
rect 33597 26367 33655 26373
rect 33597 26364 33609 26367
rect 32364 26336 33609 26364
rect 32364 26324 32370 26336
rect 33597 26333 33609 26336
rect 33643 26333 33655 26367
rect 33962 26364 33968 26376
rect 33923 26336 33968 26364
rect 33597 26327 33655 26333
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34238 26324 34244 26376
rect 34296 26364 34302 26376
rect 34532 26364 34560 26404
rect 36648 26376 36676 26404
rect 39301 26401 39313 26435
rect 39347 26432 39359 26435
rect 43714 26432 43720 26444
rect 39347 26404 43720 26432
rect 39347 26401 39359 26404
rect 39301 26395 39359 26401
rect 43714 26392 43720 26404
rect 43772 26392 43778 26444
rect 34698 26364 34704 26376
rect 34296 26336 34560 26364
rect 34659 26336 34704 26364
rect 34296 26324 34302 26336
rect 34698 26324 34704 26336
rect 34756 26324 34762 26376
rect 36630 26324 36636 26376
rect 36688 26364 36694 26376
rect 37461 26367 37519 26373
rect 37461 26364 37473 26367
rect 36688 26336 37473 26364
rect 36688 26324 36694 26336
rect 37461 26333 37473 26336
rect 37507 26333 37519 26367
rect 37461 26327 37519 26333
rect 24544 26268 25268 26296
rect 33781 26299 33839 26305
rect 24544 26256 24550 26268
rect 33781 26265 33793 26299
rect 33827 26296 33839 26299
rect 34974 26296 34980 26308
rect 33827 26268 34100 26296
rect 34935 26268 34980 26296
rect 33827 26265 33839 26268
rect 33781 26259 33839 26265
rect 34072 26240 34100 26268
rect 34974 26256 34980 26268
rect 35032 26256 35038 26308
rect 35986 26256 35992 26308
rect 36044 26256 36050 26308
rect 37642 26296 37648 26308
rect 37603 26268 37648 26296
rect 37642 26256 37648 26268
rect 37700 26256 37706 26308
rect 19429 26231 19487 26237
rect 19429 26197 19441 26231
rect 19475 26197 19487 26231
rect 33870 26228 33876 26240
rect 33831 26200 33876 26228
rect 19429 26191 19487 26197
rect 33870 26188 33876 26200
rect 33928 26188 33934 26240
rect 34054 26188 34060 26240
rect 34112 26228 34118 26240
rect 36449 26231 36507 26237
rect 36449 26228 36461 26231
rect 34112 26200 36461 26228
rect 34112 26188 34118 26200
rect 36449 26197 36461 26200
rect 36495 26228 36507 26231
rect 42150 26228 42156 26240
rect 36495 26200 42156 26228
rect 36495 26197 36507 26200
rect 36449 26191 36507 26197
rect 42150 26188 42156 26200
rect 42208 26188 42214 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 22554 26024 22560 26036
rect 22515 25996 22560 26024
rect 22554 25984 22560 25996
rect 22612 25984 22618 26036
rect 23106 26024 23112 26036
rect 23067 25996 23112 26024
rect 23106 25984 23112 25996
rect 23164 25984 23170 26036
rect 32585 26027 32643 26033
rect 32585 25993 32597 26027
rect 32631 26024 32643 26027
rect 33134 26024 33140 26036
rect 32631 25996 33140 26024
rect 32631 25993 32643 25996
rect 32585 25987 32643 25993
rect 33134 25984 33140 25996
rect 33192 25984 33198 26036
rect 33505 26027 33563 26033
rect 33505 25993 33517 26027
rect 33551 26024 33563 26027
rect 34698 26024 34704 26036
rect 33551 25996 34704 26024
rect 33551 25993 33563 25996
rect 33505 25987 33563 25993
rect 34698 25984 34704 25996
rect 34756 25984 34762 26036
rect 34974 26024 34980 26036
rect 34935 25996 34980 26024
rect 34974 25984 34980 25996
rect 35032 25984 35038 26036
rect 35621 26027 35679 26033
rect 35621 25993 35633 26027
rect 35667 26024 35679 26027
rect 35986 26024 35992 26036
rect 35667 25996 35992 26024
rect 35667 25993 35679 25996
rect 35621 25987 35679 25993
rect 35986 25984 35992 25996
rect 36044 25984 36050 26036
rect 37642 26024 37648 26036
rect 37603 25996 37648 26024
rect 37642 25984 37648 25996
rect 37700 25984 37706 26036
rect 12618 25916 12624 25968
rect 12676 25956 12682 25968
rect 12713 25959 12771 25965
rect 12713 25956 12725 25959
rect 12676 25928 12725 25956
rect 12676 25916 12682 25928
rect 12713 25925 12725 25928
rect 12759 25925 12771 25959
rect 14182 25956 14188 25968
rect 13938 25928 14188 25956
rect 12713 25919 12771 25925
rect 14182 25916 14188 25928
rect 14240 25916 14246 25968
rect 14826 25916 14832 25968
rect 14884 25956 14890 25968
rect 18506 25956 18512 25968
rect 14884 25928 15792 25956
rect 14884 25916 14890 25928
rect 11882 25888 11888 25900
rect 11843 25860 11888 25888
rect 11882 25848 11888 25860
rect 11940 25848 11946 25900
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25888 14979 25891
rect 15102 25888 15108 25900
rect 14967 25860 15108 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 15102 25848 15108 25860
rect 15160 25848 15166 25900
rect 15764 25897 15792 25928
rect 17236 25928 18512 25956
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25888 15807 25891
rect 15838 25888 15844 25900
rect 15795 25860 15844 25888
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 15838 25848 15844 25860
rect 15896 25888 15902 25900
rect 17126 25888 17132 25900
rect 15896 25860 17132 25888
rect 15896 25848 15902 25860
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 17236 25897 17264 25928
rect 18506 25916 18512 25928
rect 18564 25916 18570 25968
rect 23750 25956 23756 25968
rect 23584 25928 23756 25956
rect 17221 25891 17279 25897
rect 17221 25857 17233 25891
rect 17267 25857 17279 25891
rect 18046 25888 18052 25900
rect 18007 25860 18052 25888
rect 17221 25851 17279 25857
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22465 25891 22523 25897
rect 22465 25888 22477 25891
rect 22244 25860 22477 25888
rect 22244 25848 22250 25860
rect 22465 25857 22477 25860
rect 22511 25857 22523 25891
rect 22465 25851 22523 25857
rect 12434 25780 12440 25832
rect 12492 25820 12498 25832
rect 12492 25792 12537 25820
rect 12492 25780 12498 25792
rect 13722 25780 13728 25832
rect 13780 25820 13786 25832
rect 14185 25823 14243 25829
rect 14185 25820 14197 25823
rect 13780 25792 14197 25820
rect 13780 25780 13786 25792
rect 14185 25789 14197 25792
rect 14231 25789 14243 25823
rect 14185 25783 14243 25789
rect 15197 25823 15255 25829
rect 15197 25789 15209 25823
rect 15243 25820 15255 25823
rect 15286 25820 15292 25832
rect 15243 25792 15292 25820
rect 15243 25789 15255 25792
rect 15197 25783 15255 25789
rect 15286 25780 15292 25792
rect 15344 25780 15350 25832
rect 22480 25820 22508 25851
rect 22922 25848 22928 25900
rect 22980 25888 22986 25900
rect 23293 25891 23351 25897
rect 23293 25888 23305 25891
rect 22980 25860 23305 25888
rect 22980 25848 22986 25860
rect 23293 25857 23305 25860
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 23382 25848 23388 25900
rect 23440 25888 23446 25900
rect 23584 25897 23612 25928
rect 23750 25916 23756 25928
rect 23808 25916 23814 25968
rect 31202 25916 31208 25968
rect 31260 25956 31266 25968
rect 34054 25956 34060 25968
rect 31260 25928 33364 25956
rect 34015 25928 34060 25956
rect 31260 25916 31266 25928
rect 23569 25891 23627 25897
rect 23440 25860 23485 25888
rect 23440 25848 23446 25860
rect 23569 25857 23581 25891
rect 23615 25857 23627 25891
rect 23569 25851 23627 25857
rect 23658 25848 23664 25900
rect 23716 25888 23722 25900
rect 25406 25888 25412 25900
rect 23716 25860 23761 25888
rect 25367 25860 25412 25888
rect 23716 25848 23722 25860
rect 25406 25848 25412 25860
rect 25464 25848 25470 25900
rect 32490 25888 32496 25900
rect 32451 25860 32496 25888
rect 32490 25848 32496 25860
rect 32548 25848 32554 25900
rect 33336 25897 33364 25928
rect 34054 25916 34060 25928
rect 34112 25916 34118 25968
rect 34257 25959 34315 25965
rect 34257 25956 34269 25959
rect 34164 25928 34269 25956
rect 34164 25900 34192 25928
rect 34257 25925 34269 25928
rect 34303 25925 34315 25959
rect 34257 25919 34315 25925
rect 34422 25916 34428 25968
rect 34480 25956 34486 25968
rect 34480 25928 35112 25956
rect 34480 25916 34486 25928
rect 33321 25891 33379 25897
rect 33321 25857 33333 25891
rect 33367 25857 33379 25891
rect 33321 25851 33379 25857
rect 33962 25848 33968 25900
rect 34020 25888 34026 25900
rect 34146 25888 34152 25900
rect 34020 25860 34152 25888
rect 34020 25848 34026 25860
rect 34146 25848 34152 25860
rect 34204 25848 34210 25900
rect 34790 25848 34796 25900
rect 34848 25888 34854 25900
rect 35084 25897 35112 25928
rect 35158 25916 35164 25968
rect 35216 25956 35222 25968
rect 41414 25956 41420 25968
rect 35216 25928 41420 25956
rect 35216 25916 35222 25928
rect 41414 25916 41420 25928
rect 41472 25916 41478 25968
rect 34885 25891 34943 25897
rect 34885 25888 34897 25891
rect 34848 25860 34897 25888
rect 34848 25848 34854 25860
rect 34885 25857 34897 25860
rect 34931 25857 34943 25891
rect 34885 25851 34943 25857
rect 35069 25891 35127 25897
rect 35069 25857 35081 25891
rect 35115 25857 35127 25891
rect 35526 25888 35532 25900
rect 35487 25860 35532 25888
rect 35069 25851 35127 25857
rect 35526 25848 35532 25860
rect 35584 25848 35590 25900
rect 37550 25888 37556 25900
rect 37511 25860 37556 25888
rect 37550 25848 37556 25860
rect 37608 25848 37614 25900
rect 41506 25888 41512 25900
rect 41467 25860 41512 25888
rect 41506 25848 41512 25860
rect 41564 25848 41570 25900
rect 46750 25848 46756 25900
rect 46808 25888 46814 25900
rect 48133 25891 48191 25897
rect 48133 25888 48145 25891
rect 46808 25860 48145 25888
rect 46808 25848 46814 25860
rect 48133 25857 48145 25860
rect 48179 25857 48191 25891
rect 48133 25851 48191 25857
rect 24486 25820 24492 25832
rect 22480 25792 24492 25820
rect 24486 25780 24492 25792
rect 24544 25780 24550 25832
rect 25961 25823 26019 25829
rect 25961 25789 25973 25823
rect 26007 25789 26019 25823
rect 25961 25783 26019 25789
rect 13814 25712 13820 25764
rect 13872 25752 13878 25764
rect 15105 25755 15163 25761
rect 15105 25752 15117 25755
rect 13872 25724 15117 25752
rect 13872 25712 13878 25724
rect 15105 25721 15117 25724
rect 15151 25721 15163 25755
rect 18230 25752 18236 25764
rect 18191 25724 18236 25752
rect 15105 25715 15163 25721
rect 18230 25712 18236 25724
rect 18288 25712 18294 25764
rect 25314 25712 25320 25764
rect 25372 25752 25378 25764
rect 25976 25752 26004 25783
rect 28626 25780 28632 25832
rect 28684 25820 28690 25832
rect 29733 25823 29791 25829
rect 29733 25820 29745 25823
rect 28684 25792 29745 25820
rect 28684 25780 28690 25792
rect 29733 25789 29745 25792
rect 29779 25789 29791 25823
rect 29914 25820 29920 25832
rect 29875 25792 29920 25820
rect 29733 25783 29791 25789
rect 29914 25780 29920 25792
rect 29972 25780 29978 25832
rect 31573 25823 31631 25829
rect 31573 25789 31585 25823
rect 31619 25820 31631 25823
rect 36262 25820 36268 25832
rect 31619 25792 36268 25820
rect 31619 25789 31631 25792
rect 31573 25783 31631 25789
rect 36262 25780 36268 25792
rect 36320 25780 36326 25832
rect 36446 25780 36452 25832
rect 36504 25820 36510 25832
rect 45462 25820 45468 25832
rect 36504 25792 45468 25820
rect 36504 25780 36510 25792
rect 45462 25780 45468 25792
rect 45520 25780 45526 25832
rect 35158 25752 35164 25764
rect 25372 25724 35164 25752
rect 25372 25712 25378 25724
rect 35158 25712 35164 25724
rect 35216 25712 35222 25764
rect 11698 25684 11704 25696
rect 11659 25656 11704 25684
rect 11698 25644 11704 25656
rect 11756 25644 11762 25696
rect 14737 25687 14795 25693
rect 14737 25653 14749 25687
rect 14783 25684 14795 25687
rect 14918 25684 14924 25696
rect 14783 25656 14924 25684
rect 14783 25653 14795 25656
rect 14737 25647 14795 25653
rect 14918 25644 14924 25656
rect 14976 25644 14982 25696
rect 15841 25687 15899 25693
rect 15841 25653 15853 25687
rect 15887 25684 15899 25687
rect 15930 25684 15936 25696
rect 15887 25656 15936 25684
rect 15887 25653 15899 25656
rect 15841 25647 15899 25653
rect 15930 25644 15936 25656
rect 15988 25644 15994 25696
rect 17402 25684 17408 25696
rect 17363 25656 17408 25684
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 33870 25644 33876 25696
rect 33928 25684 33934 25696
rect 34238 25684 34244 25696
rect 33928 25656 34244 25684
rect 33928 25644 33934 25656
rect 34238 25644 34244 25656
rect 34296 25644 34302 25696
rect 34422 25684 34428 25696
rect 34383 25656 34428 25684
rect 34422 25644 34428 25656
rect 34480 25644 34486 25696
rect 34514 25644 34520 25696
rect 34572 25684 34578 25696
rect 41506 25684 41512 25696
rect 34572 25656 41512 25684
rect 34572 25644 34578 25656
rect 41506 25644 41512 25656
rect 41564 25644 41570 25696
rect 41601 25687 41659 25693
rect 41601 25653 41613 25687
rect 41647 25684 41659 25687
rect 42334 25684 42340 25696
rect 41647 25656 42340 25684
rect 41647 25653 41659 25656
rect 41601 25647 41659 25653
rect 42334 25644 42340 25656
rect 42392 25644 42398 25696
rect 47578 25644 47584 25696
rect 47636 25684 47642 25696
rect 47949 25687 48007 25693
rect 47949 25684 47961 25687
rect 47636 25656 47961 25684
rect 47636 25644 47642 25656
rect 47949 25653 47961 25656
rect 47995 25653 48007 25687
rect 47949 25647 48007 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 13078 25480 13084 25492
rect 12492 25452 13084 25480
rect 12492 25440 12498 25452
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 15286 25440 15292 25492
rect 15344 25480 15350 25492
rect 16393 25483 16451 25489
rect 16393 25480 16405 25483
rect 15344 25452 16405 25480
rect 15344 25440 15350 25452
rect 16393 25449 16405 25452
rect 16439 25449 16451 25483
rect 16393 25443 16451 25449
rect 17126 25440 17132 25492
rect 17184 25480 17190 25492
rect 17221 25483 17279 25489
rect 17221 25480 17233 25483
rect 17184 25452 17233 25480
rect 17184 25440 17190 25452
rect 17221 25449 17233 25452
rect 17267 25449 17279 25483
rect 17221 25443 17279 25449
rect 17402 25440 17408 25492
rect 17460 25480 17466 25492
rect 17460 25452 22094 25480
rect 17460 25440 17466 25452
rect 16298 25372 16304 25424
rect 16356 25412 16362 25424
rect 17957 25415 18015 25421
rect 17957 25412 17969 25415
rect 16356 25384 17969 25412
rect 16356 25372 16362 25384
rect 17957 25381 17969 25384
rect 18003 25381 18015 25415
rect 22066 25412 22094 25452
rect 25958 25440 25964 25492
rect 26016 25480 26022 25492
rect 26016 25452 31754 25480
rect 26016 25440 26022 25452
rect 30098 25412 30104 25424
rect 22066 25384 30104 25412
rect 17957 25375 18015 25381
rect 30098 25372 30104 25384
rect 30156 25412 30162 25424
rect 31726 25412 31754 25452
rect 32490 25440 32496 25492
rect 32548 25480 32554 25492
rect 32769 25483 32827 25489
rect 32769 25480 32781 25483
rect 32548 25452 32781 25480
rect 32548 25440 32554 25452
rect 32769 25449 32781 25452
rect 32815 25480 32827 25483
rect 35526 25480 35532 25492
rect 32815 25452 35532 25480
rect 32815 25449 32827 25452
rect 32769 25443 32827 25449
rect 35526 25440 35532 25452
rect 35584 25440 35590 25492
rect 39209 25483 39267 25489
rect 39209 25449 39221 25483
rect 39255 25480 39267 25483
rect 40034 25480 40040 25492
rect 39255 25452 40040 25480
rect 39255 25449 39267 25452
rect 39209 25443 39267 25449
rect 40034 25440 40040 25452
rect 40092 25440 40098 25492
rect 46658 25480 46664 25492
rect 41386 25452 46664 25480
rect 37550 25412 37556 25424
rect 30156 25384 30604 25412
rect 31726 25384 37556 25412
rect 30156 25372 30162 25384
rect 11698 25344 11704 25356
rect 11659 25316 11704 25344
rect 11698 25304 11704 25316
rect 11756 25304 11762 25356
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 12526 25344 12532 25356
rect 12023 25316 12532 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 12526 25304 12532 25316
rect 12584 25304 12590 25356
rect 14918 25344 14924 25356
rect 14879 25316 14924 25344
rect 14918 25304 14924 25316
rect 14976 25304 14982 25356
rect 18046 25344 18052 25356
rect 17788 25316 18052 25344
rect 14645 25279 14703 25285
rect 14645 25245 14657 25279
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 17037 25279 17095 25285
rect 17037 25245 17049 25279
rect 17083 25276 17095 25279
rect 17218 25276 17224 25288
rect 17083 25248 17224 25276
rect 17083 25245 17095 25248
rect 17037 25239 17095 25245
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 13262 25208 13268 25220
rect 13202 25180 13268 25208
rect 13262 25168 13268 25180
rect 13320 25168 13326 25220
rect 13354 25168 13360 25220
rect 13412 25208 13418 25220
rect 14660 25208 14688 25239
rect 17218 25236 17224 25248
rect 17276 25276 17282 25288
rect 17402 25276 17408 25288
rect 17276 25248 17408 25276
rect 17276 25236 17282 25248
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 17788 25285 17816 25316
rect 18046 25304 18052 25316
rect 18104 25344 18110 25356
rect 25406 25344 25412 25356
rect 18104 25316 25412 25344
rect 18104 25304 18110 25316
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25245 17831 25279
rect 17773 25239 17831 25245
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25245 19395 25279
rect 19337 25239 19395 25245
rect 19521 25279 19579 25285
rect 19521 25245 19533 25279
rect 19567 25276 19579 25279
rect 20714 25276 20720 25288
rect 19567 25248 20720 25276
rect 19567 25245 19579 25248
rect 19521 25239 19579 25245
rect 15194 25208 15200 25220
rect 13412 25180 13584 25208
rect 14660 25180 15200 25208
rect 13412 25168 13418 25180
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 2038 25140 2044 25152
rect 1995 25112 2044 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 12710 25100 12716 25152
rect 12768 25140 12774 25152
rect 13449 25143 13507 25149
rect 13449 25140 13461 25143
rect 12768 25112 13461 25140
rect 12768 25100 12774 25112
rect 13449 25109 13461 25112
rect 13495 25109 13507 25143
rect 13556 25140 13584 25180
rect 15194 25168 15200 25180
rect 15252 25168 15258 25220
rect 15930 25168 15936 25220
rect 15988 25168 15994 25220
rect 19352 25208 19380 25239
rect 20714 25236 20720 25248
rect 20772 25236 20778 25288
rect 21174 25276 21180 25288
rect 21135 25248 21180 25276
rect 21174 25236 21180 25248
rect 21232 25236 21238 25288
rect 21358 25276 21364 25288
rect 21319 25248 21364 25276
rect 21358 25236 21364 25248
rect 21416 25236 21422 25288
rect 24486 25276 24492 25288
rect 24447 25248 24492 25276
rect 24486 25236 24492 25248
rect 24544 25236 24550 25288
rect 25148 25285 25176 25316
rect 25406 25304 25412 25316
rect 25464 25304 25470 25356
rect 25774 25304 25780 25356
rect 25832 25344 25838 25356
rect 25958 25344 25964 25356
rect 25832 25316 25964 25344
rect 25832 25304 25838 25316
rect 25958 25304 25964 25316
rect 26016 25304 26022 25356
rect 26234 25304 26240 25356
rect 26292 25344 26298 25356
rect 26881 25347 26939 25353
rect 26881 25344 26893 25347
rect 26292 25316 26893 25344
rect 26292 25304 26298 25316
rect 26881 25313 26893 25316
rect 26927 25344 26939 25347
rect 26927 25316 30512 25344
rect 26927 25313 26939 25316
rect 26881 25307 26939 25313
rect 25133 25279 25191 25285
rect 25133 25245 25145 25279
rect 25179 25245 25191 25279
rect 25424 25276 25452 25304
rect 26605 25279 26663 25285
rect 26605 25276 26617 25279
rect 25424 25248 26617 25276
rect 25133 25239 25191 25245
rect 26605 25245 26617 25248
rect 26651 25276 26663 25279
rect 27801 25279 27859 25285
rect 27801 25276 27813 25279
rect 26651 25248 27813 25276
rect 26651 25245 26663 25248
rect 26605 25239 26663 25245
rect 27801 25245 27813 25248
rect 27847 25245 27859 25279
rect 27801 25239 27859 25245
rect 29270 25236 29276 25288
rect 29328 25276 29334 25288
rect 29638 25276 29644 25288
rect 29328 25248 29644 25276
rect 29328 25236 29334 25248
rect 29638 25236 29644 25248
rect 29696 25236 29702 25288
rect 30374 25276 30380 25288
rect 30335 25248 30380 25276
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 19426 25208 19432 25220
rect 19339 25180 19432 25208
rect 19426 25168 19432 25180
rect 19484 25208 19490 25220
rect 24670 25208 24676 25220
rect 19484 25180 24676 25208
rect 19484 25168 19490 25180
rect 24670 25168 24676 25180
rect 24728 25168 24734 25220
rect 27617 25211 27675 25217
rect 27617 25177 27629 25211
rect 27663 25208 27675 25211
rect 29288 25208 29316 25236
rect 27663 25180 29316 25208
rect 30484 25208 30512 25316
rect 30576 25276 30604 25384
rect 37550 25372 37556 25384
rect 37608 25412 37614 25424
rect 39390 25412 39396 25424
rect 37608 25384 39396 25412
rect 37608 25372 37614 25384
rect 39390 25372 39396 25384
rect 39448 25372 39454 25424
rect 31386 25304 31392 25356
rect 31444 25344 31450 25356
rect 32125 25347 32183 25353
rect 32125 25344 32137 25347
rect 31444 25316 32137 25344
rect 31444 25304 31450 25316
rect 32125 25313 32137 25316
rect 32171 25344 32183 25347
rect 41386 25344 41414 25452
rect 46658 25440 46664 25452
rect 46716 25440 46722 25492
rect 46382 25372 46388 25424
rect 46440 25412 46446 25424
rect 47949 25415 48007 25421
rect 47949 25412 47961 25415
rect 46440 25384 47961 25412
rect 46440 25372 46446 25384
rect 47949 25381 47961 25384
rect 47995 25381 48007 25415
rect 47949 25375 48007 25381
rect 41690 25344 41696 25356
rect 32171 25316 41414 25344
rect 41651 25316 41696 25344
rect 32171 25313 32183 25316
rect 32125 25307 32183 25313
rect 41690 25304 41696 25316
rect 41748 25304 41754 25356
rect 42150 25344 42156 25356
rect 42111 25316 42156 25344
rect 42150 25304 42156 25316
rect 42208 25304 42214 25356
rect 42334 25344 42340 25356
rect 42295 25316 42340 25344
rect 42334 25304 42340 25316
rect 42392 25304 42398 25356
rect 46842 25344 46848 25356
rect 46803 25316 46848 25344
rect 46842 25304 46848 25316
rect 46900 25304 46906 25356
rect 32585 25279 32643 25285
rect 32585 25276 32597 25279
rect 30576 25248 32597 25276
rect 32585 25245 32597 25248
rect 32631 25245 32643 25279
rect 39114 25276 39120 25288
rect 39075 25248 39120 25276
rect 32585 25239 32643 25245
rect 39114 25236 39120 25248
rect 39172 25236 39178 25288
rect 39853 25279 39911 25285
rect 39853 25276 39865 25279
rect 39224 25248 39865 25276
rect 30834 25208 30840 25220
rect 30484 25180 30840 25208
rect 27663 25177 27675 25180
rect 27617 25171 27675 25177
rect 30834 25168 30840 25180
rect 30892 25208 30898 25220
rect 34514 25208 34520 25220
rect 30892 25180 34520 25208
rect 30892 25168 30898 25180
rect 34514 25168 34520 25180
rect 34572 25168 34578 25220
rect 15562 25140 15568 25152
rect 13556 25112 15568 25140
rect 13449 25103 13507 25109
rect 15562 25100 15568 25112
rect 15620 25140 15626 25152
rect 19705 25143 19763 25149
rect 19705 25140 19717 25143
rect 15620 25112 19717 25140
rect 15620 25100 15626 25112
rect 19705 25109 19717 25112
rect 19751 25109 19763 25143
rect 19705 25103 19763 25109
rect 21269 25143 21327 25149
rect 21269 25109 21281 25143
rect 21315 25140 21327 25143
rect 21542 25140 21548 25152
rect 21315 25112 21548 25140
rect 21315 25109 21327 25112
rect 21269 25103 21327 25109
rect 21542 25100 21548 25112
rect 21600 25100 21606 25152
rect 24581 25143 24639 25149
rect 24581 25109 24593 25143
rect 24627 25140 24639 25143
rect 24946 25140 24952 25152
rect 24627 25112 24952 25140
rect 24627 25109 24639 25112
rect 24581 25103 24639 25109
rect 24946 25100 24952 25112
rect 25004 25100 25010 25152
rect 29825 25143 29883 25149
rect 29825 25109 29837 25143
rect 29871 25140 29883 25143
rect 30374 25140 30380 25152
rect 29871 25112 30380 25140
rect 29871 25109 29883 25112
rect 29825 25103 29883 25109
rect 30374 25100 30380 25112
rect 30432 25100 30438 25152
rect 33962 25100 33968 25152
rect 34020 25140 34026 25152
rect 39224 25140 39252 25248
rect 39853 25245 39865 25248
rect 39899 25245 39911 25279
rect 39853 25239 39911 25245
rect 45186 25236 45192 25288
rect 45244 25276 45250 25288
rect 45465 25279 45523 25285
rect 45465 25276 45477 25279
rect 45244 25248 45477 25276
rect 45244 25236 45250 25248
rect 45465 25245 45477 25248
rect 45511 25245 45523 25279
rect 45465 25239 45523 25245
rect 40034 25208 40040 25220
rect 39995 25180 40040 25208
rect 40034 25168 40040 25180
rect 40092 25168 40098 25220
rect 43990 25208 43996 25220
rect 43951 25180 43996 25208
rect 43990 25168 43996 25180
rect 44048 25168 44054 25220
rect 45646 25208 45652 25220
rect 45607 25180 45652 25208
rect 45646 25168 45652 25180
rect 45704 25168 45710 25220
rect 34020 25112 39252 25140
rect 34020 25100 34026 25112
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 12434 24936 12440 24948
rect 12406 24896 12440 24936
rect 12492 24896 12498 24948
rect 12618 24896 12624 24948
rect 12676 24936 12682 24948
rect 13081 24939 13139 24945
rect 13081 24936 13093 24939
rect 12676 24908 13093 24936
rect 12676 24896 12682 24908
rect 13081 24905 13093 24908
rect 13127 24936 13139 24939
rect 13722 24936 13728 24948
rect 13127 24908 13728 24936
rect 13127 24905 13139 24908
rect 13081 24899 13139 24905
rect 13722 24896 13728 24908
rect 13780 24936 13786 24948
rect 14737 24939 14795 24945
rect 14737 24936 14749 24939
rect 13780 24908 14749 24936
rect 13780 24896 13786 24908
rect 14737 24905 14749 24908
rect 14783 24905 14795 24939
rect 19426 24936 19432 24948
rect 19387 24908 19432 24936
rect 14737 24899 14795 24905
rect 19426 24896 19432 24908
rect 19484 24896 19490 24948
rect 20530 24896 20536 24948
rect 20588 24936 20594 24948
rect 20809 24939 20867 24945
rect 20809 24936 20821 24939
rect 20588 24908 20821 24936
rect 20588 24896 20594 24908
rect 20809 24905 20821 24908
rect 20855 24905 20867 24939
rect 20809 24899 20867 24905
rect 29825 24939 29883 24945
rect 29825 24905 29837 24939
rect 29871 24936 29883 24939
rect 29914 24936 29920 24948
rect 29871 24908 29920 24936
rect 29871 24905 29883 24908
rect 29825 24899 29883 24905
rect 29914 24896 29920 24908
rect 29972 24896 29978 24948
rect 34238 24896 34244 24948
rect 34296 24896 34302 24948
rect 12161 24871 12219 24877
rect 12161 24837 12173 24871
rect 12207 24868 12219 24871
rect 12406 24868 12434 24896
rect 14645 24871 14703 24877
rect 14645 24868 14657 24871
rect 12207 24840 12434 24868
rect 12728 24840 14657 24868
rect 12207 24837 12219 24840
rect 12161 24831 12219 24837
rect 12066 24800 12072 24812
rect 12027 24772 12072 24800
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24800 12495 24803
rect 12728 24800 12756 24840
rect 14645 24837 14657 24840
rect 14691 24837 14703 24871
rect 14829 24871 14887 24877
rect 14829 24868 14841 24871
rect 14645 24831 14703 24837
rect 14752 24840 14841 24868
rect 12483 24772 12756 24800
rect 12483 24769 12495 24772
rect 12437 24763 12495 24769
rect 12253 24735 12311 24741
rect 12253 24701 12265 24735
rect 12299 24732 12311 24735
rect 12618 24732 12624 24744
rect 12299 24704 12624 24732
rect 12299 24701 12311 24704
rect 12253 24695 12311 24701
rect 12618 24692 12624 24704
rect 12676 24692 12682 24744
rect 12728 24676 12756 24772
rect 13078 24760 13084 24812
rect 13136 24800 13142 24812
rect 13173 24803 13231 24809
rect 13173 24800 13185 24803
rect 13136 24772 13185 24800
rect 13136 24760 13142 24772
rect 13173 24769 13185 24772
rect 13219 24769 13231 24803
rect 13173 24763 13231 24769
rect 13265 24803 13323 24809
rect 13265 24769 13277 24803
rect 13311 24800 13323 24803
rect 13354 24800 13360 24812
rect 13311 24772 13360 24800
rect 13311 24769 13323 24772
rect 13265 24763 13323 24769
rect 13188 24732 13216 24763
rect 13354 24760 13360 24772
rect 13412 24760 13418 24812
rect 13449 24803 13507 24809
rect 13449 24769 13461 24803
rect 13495 24800 13507 24803
rect 13814 24800 13820 24812
rect 13495 24772 13820 24800
rect 13495 24769 13507 24772
rect 13449 24763 13507 24769
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 13538 24732 13544 24744
rect 13188 24704 13544 24732
rect 13538 24692 13544 24704
rect 13596 24732 13602 24744
rect 14752 24732 14780 24840
rect 14829 24837 14841 24840
rect 14875 24837 14887 24871
rect 15562 24868 15568 24880
rect 14829 24831 14887 24837
rect 15488 24840 15568 24868
rect 15488 24809 15516 24840
rect 15562 24828 15568 24840
rect 15620 24828 15626 24880
rect 19613 24871 19671 24877
rect 19613 24837 19625 24871
rect 19659 24868 19671 24871
rect 20714 24868 20720 24880
rect 19659 24840 20720 24868
rect 19659 24837 19671 24840
rect 19613 24831 19671 24837
rect 20714 24828 20720 24840
rect 20772 24828 20778 24880
rect 34256 24868 34284 24896
rect 40221 24871 40279 24877
rect 40221 24868 40233 24871
rect 31956 24840 32444 24868
rect 15473 24803 15531 24809
rect 15473 24769 15485 24803
rect 15519 24769 15531 24803
rect 15473 24763 15531 24769
rect 15657 24803 15715 24809
rect 15657 24769 15669 24803
rect 15703 24769 15715 24803
rect 15657 24763 15715 24769
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 13596 24704 14780 24732
rect 13596 24692 13602 24704
rect 15102 24692 15108 24744
rect 15160 24732 15166 24744
rect 15565 24735 15623 24741
rect 15565 24732 15577 24735
rect 15160 24704 15577 24732
rect 15160 24692 15166 24704
rect 15565 24701 15577 24704
rect 15611 24701 15623 24735
rect 15565 24695 15623 24701
rect 12710 24624 12716 24676
rect 12768 24664 12774 24676
rect 12897 24667 12955 24673
rect 12897 24664 12909 24667
rect 12768 24636 12909 24664
rect 12768 24624 12774 24636
rect 12897 24633 12909 24636
rect 12943 24633 12955 24667
rect 12897 24627 12955 24633
rect 14461 24667 14519 24673
rect 14461 24633 14473 24667
rect 14507 24664 14519 24667
rect 15286 24664 15292 24676
rect 14507 24636 15292 24664
rect 14507 24633 14519 24636
rect 14461 24627 14519 24633
rect 15286 24624 15292 24636
rect 15344 24624 15350 24676
rect 15672 24664 15700 24763
rect 16868 24732 16896 24763
rect 16942 24760 16948 24812
rect 17000 24800 17006 24812
rect 17000 24772 17045 24800
rect 17000 24760 17006 24772
rect 17126 24760 17132 24812
rect 17184 24800 17190 24812
rect 17589 24803 17647 24809
rect 17589 24800 17601 24803
rect 17184 24772 17601 24800
rect 17184 24760 17190 24772
rect 17589 24769 17601 24772
rect 17635 24769 17647 24803
rect 17589 24763 17647 24769
rect 19518 24760 19524 24812
rect 19576 24800 19582 24812
rect 19576 24772 19621 24800
rect 19576 24760 19582 24772
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 20625 24803 20683 24809
rect 20625 24800 20637 24803
rect 20220 24772 20637 24800
rect 20220 24760 20226 24772
rect 20625 24769 20637 24772
rect 20671 24769 20683 24803
rect 20625 24763 20683 24769
rect 20898 24760 20904 24812
rect 20956 24800 20962 24812
rect 21818 24800 21824 24812
rect 20956 24772 21001 24800
rect 21779 24772 21824 24800
rect 20956 24760 20962 24772
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 23201 24803 23259 24809
rect 23201 24769 23213 24803
rect 23247 24769 23259 24803
rect 26142 24800 26148 24812
rect 26103 24772 26148 24800
rect 23201 24763 23259 24769
rect 23216 24732 23244 24763
rect 26142 24760 26148 24772
rect 26200 24760 26206 24812
rect 26510 24760 26516 24812
rect 26568 24800 26574 24812
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26568 24772 26985 24800
rect 26568 24760 26574 24772
rect 26973 24769 26985 24772
rect 27019 24769 27031 24803
rect 26973 24763 27031 24769
rect 27614 24760 27620 24812
rect 27672 24800 27678 24812
rect 27801 24803 27859 24809
rect 27801 24800 27813 24803
rect 27672 24772 27813 24800
rect 27672 24760 27678 24772
rect 27801 24769 27813 24772
rect 27847 24800 27859 24803
rect 28445 24803 28503 24809
rect 28445 24800 28457 24803
rect 27847 24772 28457 24800
rect 27847 24769 27859 24772
rect 27801 24763 27859 24769
rect 28445 24769 28457 24772
rect 28491 24769 28503 24803
rect 28445 24763 28503 24769
rect 29733 24803 29791 24809
rect 29733 24769 29745 24803
rect 29779 24800 29791 24803
rect 30374 24800 30380 24812
rect 29779 24772 30380 24800
rect 29779 24769 29791 24772
rect 29733 24763 29791 24769
rect 30374 24760 30380 24772
rect 30432 24760 30438 24812
rect 31294 24760 31300 24812
rect 31352 24800 31358 24812
rect 31956 24800 31984 24840
rect 32122 24800 32128 24812
rect 31352 24772 31984 24800
rect 32083 24772 32128 24800
rect 31352 24760 31358 24772
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 32416 24800 32444 24840
rect 34072 24840 34284 24868
rect 40052 24840 40233 24868
rect 33870 24800 33876 24812
rect 32416 24772 33876 24800
rect 32309 24763 32367 24769
rect 16868 24704 23244 24732
rect 15672 24636 19196 24664
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 15013 24599 15071 24605
rect 12492 24568 12537 24596
rect 12492 24556 12498 24568
rect 15013 24565 15025 24599
rect 15059 24596 15071 24599
rect 15672 24596 15700 24636
rect 17678 24596 17684 24608
rect 15059 24568 15700 24596
rect 17639 24568 17684 24596
rect 15059 24565 15071 24568
rect 15013 24559 15071 24565
rect 17678 24556 17684 24568
rect 17736 24556 17742 24608
rect 19168 24596 19196 24636
rect 19242 24624 19248 24676
rect 19300 24664 19306 24676
rect 20625 24667 20683 24673
rect 19300 24636 19345 24664
rect 19300 24624 19306 24636
rect 20625 24633 20637 24667
rect 20671 24664 20683 24667
rect 21174 24664 21180 24676
rect 20671 24636 21180 24664
rect 20671 24633 20683 24636
rect 20625 24627 20683 24633
rect 21174 24624 21180 24636
rect 21232 24624 21238 24676
rect 19518 24596 19524 24608
rect 19168 24568 19524 24596
rect 19518 24556 19524 24568
rect 19576 24556 19582 24608
rect 19797 24599 19855 24605
rect 19797 24565 19809 24599
rect 19843 24596 19855 24599
rect 19978 24596 19984 24608
rect 19843 24568 19984 24596
rect 19843 24565 19855 24568
rect 19797 24559 19855 24565
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 21266 24556 21272 24608
rect 21324 24596 21330 24608
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21324 24568 21833 24596
rect 21324 24556 21330 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 23216 24596 23244 24704
rect 23382 24692 23388 24744
rect 23440 24732 23446 24744
rect 23845 24735 23903 24741
rect 23845 24732 23857 24735
rect 23440 24704 23857 24732
rect 23440 24692 23446 24704
rect 23845 24701 23857 24704
rect 23891 24701 23903 24735
rect 23845 24695 23903 24701
rect 24029 24735 24087 24741
rect 24029 24701 24041 24735
rect 24075 24701 24087 24735
rect 24029 24695 24087 24701
rect 25685 24735 25743 24741
rect 25685 24701 25697 24735
rect 25731 24732 25743 24735
rect 28718 24732 28724 24744
rect 25731 24704 28724 24732
rect 25731 24701 25743 24704
rect 25685 24695 25743 24701
rect 23293 24667 23351 24673
rect 23293 24633 23305 24667
rect 23339 24664 23351 24667
rect 24044 24664 24072 24695
rect 28718 24692 28724 24704
rect 28776 24692 28782 24744
rect 31110 24732 31116 24744
rect 31071 24704 31116 24732
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 31662 24692 31668 24744
rect 31720 24732 31726 24744
rect 32324 24732 32352 24763
rect 33870 24760 33876 24772
rect 33928 24760 33934 24812
rect 34072 24809 34100 24840
rect 34057 24803 34115 24809
rect 34057 24769 34069 24803
rect 34103 24769 34115 24803
rect 34057 24763 34115 24769
rect 34238 24760 34244 24812
rect 34296 24800 34302 24812
rect 34885 24803 34943 24809
rect 34885 24800 34897 24803
rect 34296 24772 34897 24800
rect 34296 24760 34302 24772
rect 34885 24769 34897 24772
rect 34931 24769 34943 24803
rect 34885 24763 34943 24769
rect 36262 24760 36268 24812
rect 36320 24760 36326 24812
rect 38746 24800 38752 24812
rect 36372 24772 36768 24800
rect 38707 24772 38752 24800
rect 31720 24704 32352 24732
rect 31720 24692 31726 24704
rect 32398 24692 32404 24744
rect 32456 24732 32462 24744
rect 33962 24732 33968 24744
rect 32456 24704 33968 24732
rect 32456 24692 32462 24704
rect 33962 24692 33968 24704
rect 34020 24692 34026 24744
rect 34146 24732 34152 24744
rect 34107 24704 34152 24732
rect 34146 24692 34152 24704
rect 34204 24692 34210 24744
rect 34425 24735 34483 24741
rect 34425 24701 34437 24735
rect 34471 24732 34483 24735
rect 35161 24735 35219 24741
rect 35161 24732 35173 24735
rect 34471 24704 35173 24732
rect 34471 24701 34483 24704
rect 34425 24695 34483 24701
rect 35161 24701 35173 24704
rect 35207 24701 35219 24735
rect 35161 24695 35219 24701
rect 35250 24692 35256 24744
rect 35308 24732 35314 24744
rect 36372 24732 36400 24772
rect 36630 24732 36636 24744
rect 35308 24704 36400 24732
rect 36591 24704 36636 24732
rect 35308 24692 35314 24704
rect 36630 24692 36636 24704
rect 36688 24692 36694 24744
rect 36740 24732 36768 24772
rect 38746 24760 38752 24772
rect 38804 24760 38810 24812
rect 39390 24800 39396 24812
rect 39351 24772 39396 24800
rect 39390 24760 39396 24772
rect 39448 24760 39454 24812
rect 39485 24803 39543 24809
rect 39485 24769 39497 24803
rect 39531 24800 39543 24803
rect 40052 24800 40080 24840
rect 40221 24837 40233 24840
rect 40267 24837 40279 24871
rect 40221 24831 40279 24837
rect 44910 24800 44916 24812
rect 39531 24772 40080 24800
rect 44871 24772 44916 24800
rect 39531 24769 39543 24772
rect 39485 24763 39543 24769
rect 44910 24760 44916 24772
rect 44968 24760 44974 24812
rect 45005 24803 45063 24809
rect 45005 24769 45017 24803
rect 45051 24800 45063 24803
rect 45646 24800 45652 24812
rect 45051 24772 45652 24800
rect 45051 24769 45063 24772
rect 45005 24763 45063 24769
rect 45646 24760 45652 24772
rect 45704 24760 45710 24812
rect 47210 24760 47216 24812
rect 47268 24800 47274 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47268 24772 47593 24800
rect 47268 24760 47274 24772
rect 47581 24769 47593 24772
rect 47627 24800 47639 24803
rect 47946 24800 47952 24812
rect 47627 24772 47952 24800
rect 47627 24769 47639 24772
rect 47581 24763 47639 24769
rect 47946 24760 47952 24772
rect 48004 24760 48010 24812
rect 40037 24735 40095 24741
rect 40037 24732 40049 24735
rect 36740 24704 40049 24732
rect 40037 24701 40049 24704
rect 40083 24701 40095 24735
rect 41230 24732 41236 24744
rect 41191 24704 41236 24732
rect 40037 24695 40095 24701
rect 41230 24692 41236 24704
rect 41288 24692 41294 24744
rect 23339 24636 24072 24664
rect 23339 24633 23351 24636
rect 23293 24627 23351 24633
rect 24762 24624 24768 24676
rect 24820 24664 24826 24676
rect 45554 24664 45560 24676
rect 24820 24636 35020 24664
rect 24820 24624 24826 24636
rect 26234 24596 26240 24608
rect 23216 24568 26240 24596
rect 21821 24559 21879 24565
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 26329 24599 26387 24605
rect 26329 24565 26341 24599
rect 26375 24596 26387 24599
rect 26418 24596 26424 24608
rect 26375 24568 26424 24596
rect 26375 24565 26387 24568
rect 26329 24559 26387 24565
rect 26418 24556 26424 24568
rect 26476 24556 26482 24608
rect 26970 24596 26976 24608
rect 26931 24568 26976 24596
rect 26970 24556 26976 24568
rect 27028 24556 27034 24608
rect 27890 24596 27896 24608
rect 27851 24568 27896 24596
rect 27890 24556 27896 24568
rect 27948 24556 27954 24608
rect 28534 24596 28540 24608
rect 28495 24568 28540 24596
rect 28534 24556 28540 24568
rect 28592 24556 28598 24608
rect 31938 24556 31944 24608
rect 31996 24596 32002 24608
rect 32125 24599 32183 24605
rect 32125 24596 32137 24599
rect 31996 24568 32137 24596
rect 31996 24556 32002 24568
rect 32125 24565 32137 24568
rect 32171 24565 32183 24599
rect 32125 24559 32183 24565
rect 32766 24556 32772 24608
rect 32824 24596 32830 24608
rect 34790 24596 34796 24608
rect 32824 24568 34796 24596
rect 32824 24556 32830 24568
rect 34790 24556 34796 24568
rect 34848 24556 34854 24608
rect 34992 24596 35020 24636
rect 36188 24636 45560 24664
rect 36188 24596 36216 24636
rect 45554 24624 45560 24636
rect 45612 24624 45618 24676
rect 34992 24568 36216 24596
rect 38841 24599 38899 24605
rect 38841 24565 38853 24599
rect 38887 24596 38899 24599
rect 39022 24596 39028 24608
rect 38887 24568 39028 24596
rect 38887 24565 38899 24568
rect 38841 24559 38899 24565
rect 39022 24556 39028 24568
rect 39080 24556 39086 24608
rect 46290 24556 46296 24608
rect 46348 24596 46354 24608
rect 47029 24599 47087 24605
rect 47029 24596 47041 24599
rect 46348 24568 47041 24596
rect 46348 24556 46354 24568
rect 47029 24565 47041 24568
rect 47075 24565 47087 24599
rect 47670 24596 47676 24608
rect 47631 24568 47676 24596
rect 47029 24559 47087 24565
rect 47670 24556 47676 24568
rect 47728 24556 47734 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 12437 24395 12495 24401
rect 12437 24361 12449 24395
rect 12483 24392 12495 24395
rect 12526 24392 12532 24404
rect 12483 24364 12532 24392
rect 12483 24361 12495 24364
rect 12437 24355 12495 24361
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 15194 24392 15200 24404
rect 15155 24364 15200 24392
rect 15194 24352 15200 24364
rect 15252 24352 15258 24404
rect 20714 24392 20720 24404
rect 20675 24364 20720 24392
rect 20714 24352 20720 24364
rect 20772 24352 20778 24404
rect 32306 24392 32312 24404
rect 28736 24364 32312 24392
rect 12066 24284 12072 24336
rect 12124 24324 12130 24336
rect 13541 24327 13599 24333
rect 13541 24324 13553 24327
rect 12124 24296 13553 24324
rect 12124 24284 12130 24296
rect 13541 24293 13553 24296
rect 13587 24293 13599 24327
rect 28736 24324 28764 24364
rect 32306 24352 32312 24364
rect 32364 24352 32370 24404
rect 32401 24395 32459 24401
rect 32401 24361 32413 24395
rect 32447 24392 32459 24395
rect 32490 24392 32496 24404
rect 32447 24364 32496 24392
rect 32447 24361 32459 24364
rect 32401 24355 32459 24361
rect 32490 24352 32496 24364
rect 32548 24352 32554 24404
rect 34057 24395 34115 24401
rect 34057 24361 34069 24395
rect 34103 24392 34115 24395
rect 34238 24392 34244 24404
rect 34103 24364 34244 24392
rect 34103 24361 34115 24364
rect 34057 24355 34115 24361
rect 34238 24352 34244 24364
rect 34296 24352 34302 24404
rect 35897 24395 35955 24401
rect 35897 24361 35909 24395
rect 35943 24392 35955 24395
rect 36262 24392 36268 24404
rect 35943 24364 36268 24392
rect 35943 24361 35955 24364
rect 35897 24355 35955 24361
rect 36262 24352 36268 24364
rect 36320 24352 36326 24404
rect 38746 24352 38752 24404
rect 38804 24392 38810 24404
rect 44910 24392 44916 24404
rect 38804 24364 44916 24392
rect 38804 24352 38810 24364
rect 44910 24352 44916 24364
rect 44968 24352 44974 24404
rect 13541 24287 13599 24293
rect 28644 24296 28764 24324
rect 13556 24256 13584 24287
rect 20898 24256 20904 24268
rect 13556 24228 20904 24256
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 21266 24256 21272 24268
rect 21227 24228 21272 24256
rect 21266 24216 21272 24228
rect 21324 24216 21330 24268
rect 21542 24256 21548 24268
rect 21503 24228 21548 24256
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 25682 24256 25688 24268
rect 25643 24228 25688 24256
rect 25682 24216 25688 24228
rect 25740 24216 25746 24268
rect 26050 24256 26056 24268
rect 25792 24228 26056 24256
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 12621 24191 12679 24197
rect 12492 24160 12537 24188
rect 12492 24148 12498 24160
rect 12621 24157 12633 24191
rect 12667 24188 12679 24191
rect 13814 24188 13820 24200
rect 12667 24160 13820 24188
rect 12667 24157 12679 24160
rect 12621 24151 12679 24157
rect 13814 24148 13820 24160
rect 13872 24148 13878 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 15930 24188 15936 24200
rect 15151 24160 15936 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 15930 24148 15936 24160
rect 15988 24148 15994 24200
rect 16942 24188 16948 24200
rect 16903 24160 16948 24188
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 19242 24148 19248 24200
rect 19300 24188 19306 24200
rect 19300 24160 19472 24188
rect 19300 24148 19306 24160
rect 13354 24120 13360 24132
rect 13315 24092 13360 24120
rect 13354 24080 13360 24092
rect 13412 24080 13418 24132
rect 14458 24080 14464 24132
rect 14516 24120 14522 24132
rect 16758 24120 16764 24132
rect 14516 24092 16764 24120
rect 14516 24080 14522 24092
rect 16758 24080 16764 24092
rect 16816 24080 16822 24132
rect 17221 24123 17279 24129
rect 17221 24089 17233 24123
rect 17267 24089 17279 24123
rect 17221 24083 17279 24089
rect 15933 24055 15991 24061
rect 15933 24021 15945 24055
rect 15979 24052 15991 24055
rect 16666 24052 16672 24064
rect 15979 24024 16672 24052
rect 15979 24021 15991 24024
rect 15933 24015 15991 24021
rect 16666 24012 16672 24024
rect 16724 24012 16730 24064
rect 17236 24052 17264 24083
rect 17678 24080 17684 24132
rect 17736 24080 17742 24132
rect 19334 24120 19340 24132
rect 19295 24092 19340 24120
rect 19334 24080 19340 24092
rect 19392 24080 19398 24132
rect 19444 24120 19472 24160
rect 19518 24148 19524 24200
rect 19576 24188 19582 24200
rect 19705 24191 19763 24197
rect 19705 24188 19717 24191
rect 19576 24160 19717 24188
rect 19576 24148 19582 24160
rect 19705 24157 19717 24160
rect 19751 24157 19763 24191
rect 20438 24188 20444 24200
rect 20399 24160 20444 24188
rect 19705 24151 19763 24157
rect 20438 24148 20444 24160
rect 20496 24148 20502 24200
rect 25792 24197 25820 24228
rect 26050 24216 26056 24228
rect 26108 24256 26114 24268
rect 28644 24265 28672 24296
rect 30558 24284 30564 24336
rect 30616 24324 30622 24336
rect 31662 24324 31668 24336
rect 30616 24296 31668 24324
rect 30616 24284 30622 24296
rect 31662 24284 31668 24296
rect 31720 24324 31726 24336
rect 33226 24324 33232 24336
rect 31720 24296 33232 24324
rect 31720 24284 31726 24296
rect 33226 24284 33232 24296
rect 33284 24284 33290 24336
rect 33413 24327 33471 24333
rect 33413 24293 33425 24327
rect 33459 24324 33471 24327
rect 34146 24324 34152 24336
rect 33459 24296 34152 24324
rect 33459 24293 33471 24296
rect 33413 24287 33471 24293
rect 34146 24284 34152 24296
rect 34204 24284 34210 24336
rect 35250 24324 35256 24336
rect 35211 24296 35256 24324
rect 35250 24284 35256 24296
rect 35308 24284 35314 24336
rect 40770 24324 40776 24336
rect 36556 24296 40776 24324
rect 28629 24259 28687 24265
rect 28629 24256 28641 24259
rect 26108 24228 28641 24256
rect 26108 24216 26114 24228
rect 28629 24225 28641 24228
rect 28675 24225 28687 24259
rect 28629 24219 28687 24225
rect 28718 24216 28724 24268
rect 28776 24256 28782 24268
rect 36556 24256 36584 24296
rect 40770 24284 40776 24296
rect 40828 24284 40834 24336
rect 47486 24324 47492 24336
rect 41386 24296 47492 24324
rect 38562 24256 38568 24268
rect 28776 24228 36584 24256
rect 38523 24228 38568 24256
rect 28776 24216 28782 24228
rect 38562 24216 38568 24228
rect 38620 24216 38626 24268
rect 39945 24259 40003 24265
rect 39945 24225 39957 24259
rect 39991 24225 40003 24259
rect 39945 24219 40003 24225
rect 20533 24191 20591 24197
rect 20533 24157 20545 24191
rect 20579 24157 20591 24191
rect 20533 24151 20591 24157
rect 24581 24191 24639 24197
rect 24581 24157 24593 24191
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 25777 24191 25835 24197
rect 25777 24157 25789 24191
rect 25823 24157 25835 24191
rect 25777 24151 25835 24157
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 19444 24092 19625 24120
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 19613 24083 19671 24089
rect 20346 24080 20352 24132
rect 20404 24120 20410 24132
rect 20548 24120 20576 24151
rect 22830 24120 22836 24132
rect 20404 24092 20576 24120
rect 22770 24092 22836 24120
rect 20404 24080 20410 24092
rect 22830 24080 22836 24092
rect 22888 24080 22894 24132
rect 24596 24120 24624 24151
rect 26326 24148 26332 24200
rect 26384 24188 26390 24200
rect 26605 24191 26663 24197
rect 26605 24188 26617 24191
rect 26384 24160 26617 24188
rect 26384 24148 26390 24160
rect 26605 24157 26617 24160
rect 26651 24157 26663 24191
rect 26605 24151 26663 24157
rect 29546 24148 29552 24200
rect 29604 24188 29610 24200
rect 29641 24191 29699 24197
rect 29641 24188 29653 24191
rect 29604 24160 29653 24188
rect 29604 24148 29610 24160
rect 29641 24157 29653 24160
rect 29687 24157 29699 24191
rect 30466 24188 30472 24200
rect 30427 24160 30472 24188
rect 29641 24151 29699 24157
rect 30466 24148 30472 24160
rect 30524 24148 30530 24200
rect 31294 24188 31300 24200
rect 31220 24160 31300 24188
rect 26510 24120 26516 24132
rect 24596 24092 26516 24120
rect 26510 24080 26516 24092
rect 26568 24080 26574 24132
rect 26881 24123 26939 24129
rect 26881 24089 26893 24123
rect 26927 24089 26939 24123
rect 26881 24083 26939 24089
rect 18598 24052 18604 24064
rect 17236 24024 18604 24052
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 18693 24055 18751 24061
rect 18693 24021 18705 24055
rect 18739 24052 18751 24055
rect 19426 24052 19432 24064
rect 18739 24024 19432 24052
rect 18739 24021 18751 24024
rect 18693 24015 18751 24021
rect 19426 24012 19432 24024
rect 19484 24052 19490 24064
rect 19521 24055 19579 24061
rect 19521 24052 19533 24055
rect 19484 24024 19533 24052
rect 19484 24012 19490 24024
rect 19521 24021 19533 24024
rect 19567 24021 19579 24055
rect 19521 24015 19579 24021
rect 19889 24055 19947 24061
rect 19889 24021 19901 24055
rect 19935 24052 19947 24055
rect 20530 24052 20536 24064
rect 19935 24024 20536 24052
rect 19935 24021 19947 24024
rect 19889 24015 19947 24021
rect 20530 24012 20536 24024
rect 20588 24012 20594 24064
rect 21910 24012 21916 24064
rect 21968 24052 21974 24064
rect 23017 24055 23075 24061
rect 23017 24052 23029 24055
rect 21968 24024 23029 24052
rect 21968 24012 21974 24024
rect 23017 24021 23029 24024
rect 23063 24021 23075 24055
rect 23017 24015 23075 24021
rect 23934 24012 23940 24064
rect 23992 24052 23998 24064
rect 24673 24055 24731 24061
rect 24673 24052 24685 24055
rect 23992 24024 24685 24052
rect 23992 24012 23998 24024
rect 24673 24021 24685 24024
rect 24719 24021 24731 24055
rect 24673 24015 24731 24021
rect 26145 24055 26203 24061
rect 26145 24021 26157 24055
rect 26191 24052 26203 24055
rect 26896 24052 26924 24083
rect 27890 24080 27896 24132
rect 27948 24080 27954 24132
rect 30374 24080 30380 24132
rect 30432 24120 30438 24132
rect 31220 24129 31248 24160
rect 31294 24148 31300 24160
rect 31352 24148 31358 24200
rect 32766 24188 32772 24200
rect 32232 24160 32772 24188
rect 31205 24123 31263 24129
rect 31205 24120 31217 24123
rect 30432 24092 31217 24120
rect 30432 24080 30438 24092
rect 31205 24089 31217 24092
rect 31251 24089 31263 24123
rect 32030 24120 32036 24132
rect 31205 24083 31263 24089
rect 31312 24092 32036 24120
rect 29730 24052 29736 24064
rect 26191 24024 26924 24052
rect 29691 24024 29736 24052
rect 26191 24021 26203 24024
rect 26145 24015 26203 24021
rect 29730 24012 29736 24024
rect 29788 24012 29794 24064
rect 29822 24012 29828 24064
rect 29880 24052 29886 24064
rect 31312 24052 31340 24092
rect 32030 24080 32036 24092
rect 32088 24080 32094 24132
rect 32232 24129 32260 24160
rect 32766 24148 32772 24160
rect 32824 24148 32830 24200
rect 33134 24188 33140 24200
rect 33095 24160 33140 24188
rect 33134 24148 33140 24160
rect 33192 24148 33198 24200
rect 33229 24191 33287 24197
rect 33229 24157 33241 24191
rect 33275 24157 33287 24191
rect 33229 24151 33287 24157
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 34238 24188 34244 24200
rect 34011 24160 34244 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 32217 24123 32275 24129
rect 32217 24089 32229 24123
rect 32263 24089 32275 24123
rect 32433 24123 32491 24129
rect 32433 24120 32445 24123
rect 32217 24083 32275 24089
rect 32416 24089 32445 24120
rect 32479 24120 32491 24123
rect 33244 24120 33272 24151
rect 34238 24148 34244 24160
rect 34296 24148 34302 24200
rect 35161 24191 35219 24197
rect 35161 24157 35173 24191
rect 35207 24188 35219 24191
rect 35526 24188 35532 24200
rect 35207 24160 35532 24188
rect 35207 24157 35219 24160
rect 35161 24151 35219 24157
rect 35526 24148 35532 24160
rect 35584 24188 35590 24200
rect 35805 24191 35863 24197
rect 35805 24188 35817 24191
rect 35584 24160 35817 24188
rect 35584 24148 35590 24160
rect 35805 24157 35817 24160
rect 35851 24157 35863 24191
rect 35805 24151 35863 24157
rect 36078 24148 36084 24200
rect 36136 24188 36142 24200
rect 37001 24191 37059 24197
rect 37001 24188 37013 24191
rect 36136 24160 37013 24188
rect 36136 24148 36142 24160
rect 37001 24157 37013 24160
rect 37047 24157 37059 24191
rect 37001 24151 37059 24157
rect 32479 24092 33272 24120
rect 32479 24089 32491 24092
rect 32416 24083 32491 24089
rect 29880 24024 31340 24052
rect 29880 24012 29886 24024
rect 31570 24012 31576 24064
rect 31628 24052 31634 24064
rect 32416 24052 32444 24083
rect 33594 24080 33600 24132
rect 33652 24120 33658 24132
rect 36096 24120 36124 24148
rect 33652 24092 36124 24120
rect 37185 24123 37243 24129
rect 33652 24080 33658 24092
rect 37185 24089 37197 24123
rect 37231 24120 37243 24123
rect 37366 24120 37372 24132
rect 37231 24092 37372 24120
rect 37231 24089 37243 24092
rect 37185 24083 37243 24089
rect 37366 24080 37372 24092
rect 37424 24080 37430 24132
rect 38562 24080 38568 24132
rect 38620 24120 38626 24132
rect 39960 24120 39988 24219
rect 40037 24191 40095 24197
rect 40037 24157 40049 24191
rect 40083 24188 40095 24191
rect 41386 24188 41414 24296
rect 47486 24284 47492 24296
rect 47544 24284 47550 24336
rect 46290 24256 46296 24268
rect 46251 24228 46296 24256
rect 46290 24216 46296 24228
rect 46348 24216 46354 24268
rect 46477 24259 46535 24265
rect 46477 24225 46489 24259
rect 46523 24256 46535 24259
rect 47670 24256 47676 24268
rect 46523 24228 47676 24256
rect 46523 24225 46535 24228
rect 46477 24219 46535 24225
rect 47670 24216 47676 24228
rect 47728 24216 47734 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 42978 24188 42984 24200
rect 40083 24160 41414 24188
rect 42939 24160 42984 24188
rect 40083 24157 40095 24160
rect 40037 24151 40095 24157
rect 42978 24148 42984 24160
rect 43036 24148 43042 24200
rect 43162 24188 43168 24200
rect 43123 24160 43168 24188
rect 43162 24148 43168 24160
rect 43220 24148 43226 24200
rect 45002 24120 45008 24132
rect 38620 24092 39988 24120
rect 40052 24092 45008 24120
rect 38620 24080 38626 24092
rect 31628 24024 32444 24052
rect 32585 24055 32643 24061
rect 31628 24012 31634 24024
rect 32585 24021 32597 24055
rect 32631 24052 32643 24055
rect 33226 24052 33232 24064
rect 32631 24024 33232 24052
rect 32631 24021 32643 24024
rect 32585 24015 32643 24021
rect 33226 24012 33232 24024
rect 33284 24012 33290 24064
rect 33870 24012 33876 24064
rect 33928 24052 33934 24064
rect 40052 24052 40080 24092
rect 45002 24080 45008 24092
rect 45060 24080 45066 24132
rect 33928 24024 40080 24052
rect 40405 24055 40463 24061
rect 33928 24012 33934 24024
rect 40405 24021 40417 24055
rect 40451 24052 40463 24055
rect 41230 24052 41236 24064
rect 40451 24024 41236 24052
rect 40451 24021 40463 24024
rect 40405 24015 40463 24021
rect 41230 24012 41236 24024
rect 41288 24012 41294 24064
rect 43073 24055 43131 24061
rect 43073 24021 43085 24055
rect 43119 24052 43131 24055
rect 43530 24052 43536 24064
rect 43119 24024 43536 24052
rect 43119 24021 43131 24024
rect 43073 24015 43131 24021
rect 43530 24012 43536 24024
rect 43588 24012 43594 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 18417 23851 18475 23857
rect 18417 23848 18429 23851
rect 15120 23820 18429 23848
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 11882 23712 11888 23724
rect 11843 23684 11888 23712
rect 11882 23672 11888 23684
rect 11940 23672 11946 23724
rect 14826 23672 14832 23724
rect 14884 23712 14890 23724
rect 15120 23721 15148 23820
rect 18417 23817 18429 23820
rect 18463 23848 18475 23851
rect 19242 23848 19248 23860
rect 18463 23820 19248 23848
rect 18463 23817 18475 23820
rect 18417 23811 18475 23817
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 20349 23851 20407 23857
rect 20349 23817 20361 23851
rect 20395 23848 20407 23851
rect 20438 23848 20444 23860
rect 20395 23820 20444 23848
rect 20395 23817 20407 23820
rect 20349 23811 20407 23817
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 20530 23808 20536 23860
rect 20588 23848 20594 23860
rect 20717 23851 20775 23857
rect 20588 23820 20633 23848
rect 20588 23808 20594 23820
rect 20717 23817 20729 23851
rect 20763 23848 20775 23851
rect 21082 23848 21088 23860
rect 20763 23820 21088 23848
rect 20763 23817 20775 23820
rect 20717 23811 20775 23817
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 22830 23848 22836 23860
rect 22791 23820 22836 23848
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 26326 23848 26332 23860
rect 26287 23820 26332 23848
rect 26326 23808 26332 23820
rect 26384 23808 26390 23860
rect 29822 23848 29828 23860
rect 27632 23820 29828 23848
rect 16025 23783 16083 23789
rect 16025 23749 16037 23783
rect 16071 23780 16083 23783
rect 20162 23780 20168 23792
rect 16071 23752 17434 23780
rect 18984 23752 20168 23780
rect 16071 23749 16083 23752
rect 16025 23743 16083 23749
rect 15105 23715 15163 23721
rect 15105 23712 15117 23715
rect 14884 23684 15117 23712
rect 14884 23672 14890 23684
rect 15105 23681 15117 23684
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 15933 23715 15991 23721
rect 15933 23712 15945 23715
rect 15896 23684 15945 23712
rect 15896 23672 15902 23684
rect 15933 23681 15945 23684
rect 15979 23681 15991 23715
rect 16666 23712 16672 23724
rect 16627 23684 16672 23712
rect 15933 23675 15991 23681
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23613 15255 23647
rect 16945 23647 17003 23653
rect 16945 23644 16957 23647
rect 15197 23607 15255 23613
rect 16316 23616 16957 23644
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 14458 23576 14464 23588
rect 2087 23548 14464 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 14458 23536 14464 23548
rect 14516 23536 14522 23588
rect 15102 23536 15108 23588
rect 15160 23576 15166 23588
rect 15212 23576 15240 23607
rect 15160 23548 15240 23576
rect 15473 23579 15531 23585
rect 15160 23536 15166 23548
rect 15473 23545 15485 23579
rect 15519 23576 15531 23579
rect 16316 23576 16344 23616
rect 16945 23613 16957 23616
rect 16991 23613 17003 23647
rect 16945 23607 17003 23613
rect 17586 23604 17592 23656
rect 17644 23644 17650 23656
rect 18984 23644 19012 23752
rect 20162 23740 20168 23752
rect 20220 23780 20226 23792
rect 21910 23780 21916 23792
rect 20220 23752 21916 23780
rect 20220 23740 20226 23752
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 23934 23780 23940 23792
rect 23895 23752 23940 23780
rect 23934 23740 23940 23752
rect 23992 23740 23998 23792
rect 24946 23740 24952 23792
rect 25004 23740 25010 23792
rect 27632 23780 27660 23820
rect 29822 23808 29828 23820
rect 29880 23808 29886 23860
rect 31395 23851 31453 23857
rect 31395 23817 31407 23851
rect 31441 23848 31453 23851
rect 32122 23848 32128 23860
rect 31441 23820 32128 23848
rect 31441 23817 31453 23820
rect 31395 23811 31453 23817
rect 32122 23808 32128 23820
rect 32180 23808 32186 23860
rect 32769 23851 32827 23857
rect 32769 23817 32781 23851
rect 32815 23848 32827 23851
rect 32858 23848 32864 23860
rect 32815 23820 32864 23848
rect 32815 23817 32827 23820
rect 32769 23811 32827 23817
rect 32858 23808 32864 23820
rect 32916 23808 32922 23860
rect 33134 23848 33140 23860
rect 33095 23820 33140 23848
rect 33134 23808 33140 23820
rect 33192 23808 33198 23860
rect 33226 23808 33232 23860
rect 33284 23848 33290 23860
rect 36078 23848 36084 23860
rect 33284 23820 33916 23848
rect 33284 23808 33290 23820
rect 28534 23780 28540 23792
rect 25608 23752 27660 23780
rect 28474 23752 28540 23780
rect 19061 23715 19119 23721
rect 19061 23681 19073 23715
rect 19107 23712 19119 23715
rect 19426 23712 19432 23724
rect 19107 23684 19432 23712
rect 19107 23681 19119 23684
rect 19061 23675 19119 23681
rect 19426 23672 19432 23684
rect 19484 23672 19490 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23681 20499 23715
rect 21818 23712 21824 23724
rect 21779 23684 21824 23712
rect 20441 23675 20499 23681
rect 17644 23616 19012 23644
rect 19153 23647 19211 23653
rect 17644 23604 17650 23616
rect 19153 23613 19165 23647
rect 19199 23644 19211 23647
rect 19978 23644 19984 23656
rect 19199 23616 19984 23644
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 19978 23604 19984 23616
rect 20036 23604 20042 23656
rect 20162 23604 20168 23656
rect 20220 23644 20226 23656
rect 20346 23644 20352 23656
rect 20220 23616 20352 23644
rect 20220 23604 20226 23616
rect 20346 23604 20352 23616
rect 20404 23644 20410 23656
rect 20456 23644 20484 23675
rect 21818 23672 21824 23684
rect 21876 23672 21882 23724
rect 22738 23712 22744 23724
rect 22699 23684 22744 23712
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 20404 23616 20484 23644
rect 20404 23604 20410 23616
rect 15519 23548 16344 23576
rect 15519 23545 15531 23548
rect 15473 23539 15531 23545
rect 18598 23536 18604 23588
rect 18656 23576 18662 23588
rect 19429 23579 19487 23585
rect 19429 23576 19441 23579
rect 18656 23548 19441 23576
rect 18656 23536 18662 23548
rect 19429 23545 19441 23548
rect 19475 23545 19487 23579
rect 21836 23576 21864 23672
rect 23661 23647 23719 23653
rect 23661 23613 23673 23647
rect 23707 23644 23719 23647
rect 25608 23644 25636 23752
rect 28534 23740 28540 23752
rect 28592 23740 28598 23792
rect 31297 23783 31355 23789
rect 31297 23749 31309 23783
rect 31343 23780 31355 23783
rect 32876 23780 32904 23808
rect 33781 23783 33839 23789
rect 33781 23780 33793 23783
rect 31343 23752 32812 23780
rect 32876 23752 33793 23780
rect 31343 23749 31355 23752
rect 31297 23743 31355 23749
rect 32784 23724 32812 23752
rect 33781 23749 33793 23752
rect 33827 23749 33839 23783
rect 33781 23743 33839 23749
rect 26234 23672 26240 23724
rect 26292 23712 26298 23724
rect 26329 23715 26387 23721
rect 26329 23712 26341 23715
rect 26292 23684 26341 23712
rect 26292 23672 26298 23684
rect 26329 23681 26341 23684
rect 26375 23712 26387 23715
rect 26510 23712 26516 23724
rect 26375 23684 26516 23712
rect 26375 23681 26387 23684
rect 26329 23675 26387 23681
rect 26510 23672 26516 23684
rect 26568 23672 26574 23724
rect 26970 23712 26976 23724
rect 26931 23684 26976 23712
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 29638 23712 29644 23724
rect 29599 23684 29644 23712
rect 29638 23672 29644 23684
rect 29696 23672 29702 23724
rect 30650 23712 30656 23724
rect 30611 23684 30656 23712
rect 30650 23672 30656 23684
rect 30708 23672 30714 23724
rect 30926 23672 30932 23724
rect 30984 23712 30990 23724
rect 31481 23715 31539 23721
rect 31481 23712 31493 23715
rect 30984 23684 31493 23712
rect 30984 23672 30990 23684
rect 31481 23681 31493 23684
rect 31527 23681 31539 23715
rect 31481 23675 31539 23681
rect 23707 23616 25636 23644
rect 25685 23647 25743 23653
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 25685 23613 25697 23647
rect 25731 23613 25743 23647
rect 27246 23644 27252 23656
rect 27207 23616 27252 23644
rect 25685 23607 25743 23613
rect 19429 23539 19487 23545
rect 20272 23548 21864 23576
rect 11790 23508 11796 23520
rect 11751 23480 11796 23508
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 17310 23468 17316 23520
rect 17368 23508 17374 23520
rect 20272 23508 20300 23548
rect 25590 23536 25596 23588
rect 25648 23576 25654 23588
rect 25700 23576 25728 23607
rect 27246 23604 27252 23616
rect 27304 23604 27310 23656
rect 27982 23604 27988 23656
rect 28040 23644 28046 23656
rect 28626 23644 28632 23656
rect 28040 23616 28632 23644
rect 28040 23604 28046 23616
rect 28626 23604 28632 23616
rect 28684 23644 28690 23656
rect 28721 23647 28779 23653
rect 28721 23644 28733 23647
rect 28684 23616 28733 23644
rect 28684 23604 28690 23616
rect 28721 23613 28733 23616
rect 28767 23613 28779 23647
rect 31496 23644 31524 23675
rect 31570 23672 31576 23724
rect 31628 23712 31634 23724
rect 31628 23684 31673 23712
rect 31628 23672 31634 23684
rect 32766 23672 32772 23724
rect 32824 23712 32830 23724
rect 32861 23715 32919 23721
rect 32861 23712 32873 23715
rect 32824 23684 32873 23712
rect 32824 23672 32830 23684
rect 32861 23681 32873 23684
rect 32907 23681 32919 23715
rect 32861 23675 32919 23681
rect 32953 23715 33011 23721
rect 32953 23681 32965 23715
rect 32999 23681 33011 23715
rect 33594 23712 33600 23724
rect 33555 23684 33600 23712
rect 32953 23675 33011 23681
rect 32490 23644 32496 23656
rect 31496 23616 32496 23644
rect 28721 23607 28779 23613
rect 32490 23604 32496 23616
rect 32548 23644 32554 23656
rect 32968 23644 32996 23675
rect 33594 23672 33600 23684
rect 33652 23672 33658 23724
rect 33888 23721 33916 23820
rect 33980 23820 35940 23848
rect 36039 23820 36084 23848
rect 33873 23715 33931 23721
rect 33873 23681 33885 23715
rect 33919 23681 33931 23715
rect 33873 23675 33931 23681
rect 33612 23644 33640 23672
rect 32548 23616 32996 23644
rect 33428 23616 33640 23644
rect 32548 23604 32554 23616
rect 32585 23579 32643 23585
rect 25648 23548 25728 23576
rect 28276 23548 31754 23576
rect 25648 23536 25654 23548
rect 21818 23508 21824 23520
rect 17368 23480 20300 23508
rect 21779 23480 21824 23508
rect 17368 23468 17374 23480
rect 21818 23468 21824 23480
rect 21876 23468 21882 23520
rect 26602 23468 26608 23520
rect 26660 23508 26666 23520
rect 28276 23508 28304 23548
rect 26660 23480 28304 23508
rect 26660 23468 26666 23480
rect 29638 23468 29644 23520
rect 29696 23508 29702 23520
rect 29825 23511 29883 23517
rect 29825 23508 29837 23511
rect 29696 23480 29837 23508
rect 29696 23468 29702 23480
rect 29825 23477 29837 23480
rect 29871 23477 29883 23511
rect 30742 23508 30748 23520
rect 30703 23480 30748 23508
rect 29825 23471 29883 23477
rect 30742 23468 30748 23480
rect 30800 23468 30806 23520
rect 31726 23508 31754 23548
rect 32585 23545 32597 23579
rect 32631 23576 32643 23579
rect 33428 23576 33456 23616
rect 33980 23576 34008 23820
rect 35250 23740 35256 23792
rect 35308 23740 35314 23792
rect 35912 23780 35940 23820
rect 36078 23808 36084 23820
rect 36136 23808 36142 23860
rect 37366 23848 37372 23860
rect 37327 23820 37372 23848
rect 37366 23808 37372 23820
rect 37424 23808 37430 23860
rect 37476 23820 40724 23848
rect 37476 23780 37504 23820
rect 39022 23780 39028 23792
rect 35912 23752 37504 23780
rect 38983 23752 39028 23780
rect 39022 23740 39028 23752
rect 39080 23740 39086 23792
rect 40696 23789 40724 23820
rect 40770 23808 40776 23860
rect 40828 23848 40834 23860
rect 45830 23848 45836 23860
rect 40828 23820 45836 23848
rect 40828 23808 40834 23820
rect 45830 23808 45836 23820
rect 45888 23808 45894 23860
rect 40681 23783 40739 23789
rect 40681 23749 40693 23783
rect 40727 23749 40739 23783
rect 40681 23743 40739 23749
rect 45940 23752 46612 23780
rect 37274 23712 37280 23724
rect 37187 23684 37280 23712
rect 37274 23672 37280 23684
rect 37332 23712 37338 23724
rect 41325 23715 41383 23721
rect 37332 23684 38700 23712
rect 37332 23672 37338 23684
rect 34333 23647 34391 23653
rect 34333 23613 34345 23647
rect 34379 23613 34391 23647
rect 34606 23644 34612 23656
rect 34567 23616 34612 23644
rect 34333 23607 34391 23613
rect 32631 23548 33456 23576
rect 33520 23548 34008 23576
rect 32631 23545 32643 23548
rect 32585 23539 32643 23545
rect 33520 23508 33548 23548
rect 31726 23480 33548 23508
rect 33597 23511 33655 23517
rect 33597 23477 33609 23511
rect 33643 23508 33655 23511
rect 33870 23508 33876 23520
rect 33643 23480 33876 23508
rect 33643 23477 33655 23480
rect 33597 23471 33655 23477
rect 33870 23468 33876 23480
rect 33928 23468 33934 23520
rect 34348 23508 34376 23607
rect 34606 23604 34612 23616
rect 34664 23604 34670 23656
rect 38672 23576 38700 23684
rect 41325 23681 41337 23715
rect 41371 23712 41383 23715
rect 42518 23712 42524 23724
rect 41371 23684 42524 23712
rect 41371 23681 41383 23684
rect 41325 23675 41383 23681
rect 42518 23672 42524 23684
rect 42576 23672 42582 23724
rect 42794 23672 42800 23724
rect 42852 23712 42858 23724
rect 43165 23715 43223 23721
rect 43165 23712 43177 23715
rect 42852 23684 43177 23712
rect 42852 23672 42858 23684
rect 43165 23681 43177 23684
rect 43211 23681 43223 23715
rect 43530 23712 43536 23724
rect 43491 23684 43536 23712
rect 43165 23675 43223 23681
rect 43530 23672 43536 23684
rect 43588 23672 43594 23724
rect 45940 23721 45968 23752
rect 46584 23721 46612 23752
rect 45925 23715 45983 23721
rect 45925 23681 45937 23715
rect 45971 23681 45983 23715
rect 45925 23675 45983 23681
rect 46109 23715 46167 23721
rect 46109 23681 46121 23715
rect 46155 23681 46167 23715
rect 46109 23675 46167 23681
rect 46569 23715 46627 23721
rect 46569 23681 46581 23715
rect 46615 23712 46627 23715
rect 46934 23712 46940 23724
rect 46615 23684 46940 23712
rect 46615 23681 46627 23684
rect 46569 23675 46627 23681
rect 38841 23647 38899 23653
rect 38841 23613 38853 23647
rect 38887 23644 38899 23647
rect 40494 23644 40500 23656
rect 38887 23616 40500 23644
rect 38887 23613 38899 23616
rect 38841 23607 38899 23613
rect 40494 23604 40500 23616
rect 40552 23604 40558 23656
rect 41230 23644 41236 23656
rect 41191 23616 41236 23644
rect 41230 23604 41236 23616
rect 41288 23604 41294 23656
rect 44634 23644 44640 23656
rect 44595 23616 44640 23644
rect 44634 23604 44640 23616
rect 44692 23604 44698 23656
rect 46124 23644 46152 23675
rect 46934 23672 46940 23684
rect 46992 23672 46998 23724
rect 47210 23672 47216 23724
rect 47268 23712 47274 23724
rect 47581 23715 47639 23721
rect 47581 23712 47593 23715
rect 47268 23684 47593 23712
rect 47268 23672 47274 23684
rect 47581 23681 47593 23684
rect 47627 23681 47639 23715
rect 47581 23675 47639 23681
rect 46842 23644 46848 23656
rect 46124 23616 46848 23644
rect 46842 23604 46848 23616
rect 46900 23644 46906 23656
rect 47854 23644 47860 23656
rect 46900 23616 47860 23644
rect 46900 23604 46906 23616
rect 47854 23604 47860 23616
rect 47912 23604 47918 23656
rect 46017 23579 46075 23585
rect 38672 23548 44036 23576
rect 34698 23508 34704 23520
rect 34348 23480 34704 23508
rect 34698 23468 34704 23480
rect 34756 23468 34762 23520
rect 40494 23468 40500 23520
rect 40552 23508 40558 23520
rect 41601 23511 41659 23517
rect 41601 23508 41613 23511
rect 40552 23480 41613 23508
rect 40552 23468 40558 23480
rect 41601 23477 41613 23480
rect 41647 23477 41659 23511
rect 44008 23508 44036 23548
rect 46017 23545 46029 23579
rect 46063 23576 46075 23579
rect 47486 23576 47492 23588
rect 46063 23548 47492 23576
rect 46063 23545 46075 23548
rect 46017 23539 46075 23545
rect 47486 23536 47492 23548
rect 47544 23536 47550 23588
rect 46566 23508 46572 23520
rect 44008 23480 46572 23508
rect 41601 23471 41659 23477
rect 46566 23468 46572 23480
rect 46624 23468 46630 23520
rect 46842 23508 46848 23520
rect 46803 23480 46848 23508
rect 46842 23468 46848 23480
rect 46900 23468 46906 23520
rect 47026 23508 47032 23520
rect 46987 23480 47032 23508
rect 47026 23468 47032 23480
rect 47084 23468 47090 23520
rect 47670 23508 47676 23520
rect 47631 23480 47676 23508
rect 47670 23468 47676 23480
rect 47728 23468 47734 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 16942 23264 16948 23316
rect 17000 23304 17006 23316
rect 17129 23307 17187 23313
rect 17129 23304 17141 23307
rect 17000 23276 17141 23304
rect 17000 23264 17006 23276
rect 17129 23273 17141 23276
rect 17175 23273 17187 23307
rect 17129 23267 17187 23273
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 19518 23304 19524 23316
rect 19392 23276 19524 23304
rect 19392 23264 19398 23276
rect 19518 23264 19524 23276
rect 19576 23304 19582 23316
rect 23201 23307 23259 23313
rect 23201 23304 23213 23307
rect 19576 23276 23213 23304
rect 19576 23264 19582 23276
rect 23201 23273 23213 23276
rect 23247 23304 23259 23307
rect 23382 23304 23388 23316
rect 23247 23276 23388 23304
rect 23247 23273 23259 23276
rect 23201 23267 23259 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 27157 23307 27215 23313
rect 24872 23276 27108 23304
rect 15657 23239 15715 23245
rect 15657 23205 15669 23239
rect 15703 23236 15715 23239
rect 15930 23236 15936 23248
rect 15703 23208 15936 23236
rect 15703 23205 15715 23208
rect 15657 23199 15715 23205
rect 15930 23196 15936 23208
rect 15988 23236 15994 23248
rect 17310 23236 17316 23248
rect 15988 23208 17316 23236
rect 15988 23196 15994 23208
rect 17310 23196 17316 23208
rect 17368 23196 17374 23248
rect 22738 23196 22744 23248
rect 22796 23236 22802 23248
rect 24872 23236 24900 23276
rect 22796 23208 24900 23236
rect 24949 23239 25007 23245
rect 22796 23196 22802 23208
rect 24949 23205 24961 23239
rect 24995 23236 25007 23239
rect 25682 23236 25688 23248
rect 24995 23208 25688 23236
rect 24995 23205 25007 23208
rect 24949 23199 25007 23205
rect 25682 23196 25688 23208
rect 25740 23236 25746 23248
rect 27080 23236 27108 23276
rect 27157 23273 27169 23307
rect 27203 23304 27215 23307
rect 27246 23304 27252 23316
rect 27203 23276 27252 23304
rect 27203 23273 27215 23276
rect 27157 23267 27215 23273
rect 27246 23264 27252 23276
rect 27304 23264 27310 23316
rect 32030 23304 32036 23316
rect 30300 23276 32036 23304
rect 29546 23236 29552 23248
rect 25740 23208 26372 23236
rect 27080 23208 29552 23236
rect 25740 23196 25746 23208
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 11790 23168 11796 23180
rect 11563 23140 11796 23168
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 11790 23128 11796 23140
rect 11848 23128 11854 23180
rect 13538 23168 13544 23180
rect 13499 23140 13544 23168
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 19337 23171 19395 23177
rect 19337 23137 19349 23171
rect 19383 23168 19395 23171
rect 20257 23171 20315 23177
rect 20257 23168 20269 23171
rect 19383 23140 20269 23168
rect 19383 23137 19395 23140
rect 19337 23131 19395 23137
rect 20257 23137 20269 23140
rect 20303 23137 20315 23171
rect 20257 23131 20315 23137
rect 21453 23171 21511 23177
rect 21453 23137 21465 23171
rect 21499 23168 21511 23171
rect 21818 23168 21824 23180
rect 21499 23140 21824 23168
rect 21499 23137 21511 23140
rect 21453 23131 21511 23137
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 26344 23177 26372 23208
rect 29546 23196 29552 23208
rect 29604 23236 29610 23248
rect 30300 23245 30328 23276
rect 32030 23264 32036 23276
rect 32088 23264 32094 23316
rect 32766 23304 32772 23316
rect 32727 23276 32772 23304
rect 32766 23264 32772 23276
rect 32824 23264 32830 23316
rect 34698 23304 34704 23316
rect 34659 23276 34704 23304
rect 34698 23264 34704 23276
rect 34756 23264 34762 23316
rect 43162 23304 43168 23316
rect 43123 23276 43168 23304
rect 43162 23264 43168 23276
rect 43220 23264 43226 23316
rect 47762 23304 47768 23316
rect 43824 23276 47768 23304
rect 30285 23239 30343 23245
rect 30285 23236 30297 23239
rect 29604 23208 30297 23236
rect 29604 23196 29610 23208
rect 30285 23205 30297 23208
rect 30331 23205 30343 23239
rect 30285 23199 30343 23205
rect 26329 23171 26387 23177
rect 26329 23137 26341 23171
rect 26375 23137 26387 23171
rect 28442 23168 28448 23180
rect 28403 23140 28448 23168
rect 26329 23131 26387 23137
rect 28442 23128 28448 23140
rect 28500 23128 28506 23180
rect 28905 23171 28963 23177
rect 28905 23137 28917 23171
rect 28951 23168 28963 23171
rect 28994 23168 29000 23180
rect 28951 23140 29000 23168
rect 28951 23137 28963 23140
rect 28905 23131 28963 23137
rect 28994 23128 29000 23140
rect 29052 23128 29058 23180
rect 30742 23128 30748 23180
rect 30800 23168 30806 23180
rect 31021 23171 31079 23177
rect 31021 23168 31033 23171
rect 30800 23140 31033 23168
rect 30800 23128 30806 23140
rect 31021 23137 31033 23140
rect 31067 23137 31079 23171
rect 31021 23131 31079 23137
rect 31297 23171 31355 23177
rect 31297 23137 31309 23171
rect 31343 23168 31355 23171
rect 31938 23168 31944 23180
rect 31343 23140 31944 23168
rect 31343 23137 31355 23140
rect 31297 23131 31355 23137
rect 31938 23128 31944 23140
rect 31996 23128 32002 23180
rect 33965 23171 34023 23177
rect 33965 23137 33977 23171
rect 34011 23168 34023 23171
rect 34606 23168 34612 23180
rect 34011 23140 34612 23168
rect 34011 23137 34023 23140
rect 33965 23131 34023 23137
rect 34606 23128 34612 23140
rect 34664 23128 34670 23180
rect 40494 23168 40500 23180
rect 40455 23140 40500 23168
rect 40494 23128 40500 23140
rect 40552 23128 40558 23180
rect 43438 23168 43444 23180
rect 42904 23140 43444 23168
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23069 15531 23103
rect 17310 23100 17316 23112
rect 17271 23072 17316 23100
rect 15473 23063 15531 23069
rect 11793 23035 11851 23041
rect 11793 23001 11805 23035
rect 11839 23032 11851 23035
rect 12066 23032 12072 23044
rect 11839 23004 12072 23032
rect 11839 23001 11851 23004
rect 11793 22995 11851 23001
rect 12066 22992 12072 23004
rect 12124 22992 12130 23044
rect 13078 23032 13084 23044
rect 13018 23004 13084 23032
rect 13078 22992 13084 23004
rect 13136 22992 13142 23044
rect 14918 22992 14924 23044
rect 14976 23032 14982 23044
rect 15488 23032 15516 23063
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 19518 23100 19524 23112
rect 19479 23072 19524 23100
rect 19518 23060 19524 23072
rect 19576 23060 19582 23112
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23100 19855 23103
rect 19978 23100 19984 23112
rect 19843 23072 19984 23100
rect 19843 23069 19855 23072
rect 19797 23063 19855 23069
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 20441 23103 20499 23109
rect 20441 23069 20453 23103
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 20456 23032 20484 23063
rect 20530 23060 20536 23112
rect 20588 23100 20594 23112
rect 20625 23103 20683 23109
rect 20625 23100 20637 23103
rect 20588 23072 20637 23100
rect 20588 23060 20594 23072
rect 20625 23069 20637 23072
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23100 20775 23103
rect 20898 23100 20904 23112
rect 20763 23072 20904 23100
rect 20763 23069 20775 23072
rect 20717 23063 20775 23069
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 22830 23060 22836 23112
rect 22888 23060 22894 23112
rect 24857 23103 24915 23109
rect 24857 23069 24869 23103
rect 24903 23069 24915 23103
rect 24857 23063 24915 23069
rect 21729 23035 21787 23041
rect 21729 23032 21741 23035
rect 14976 23004 19840 23032
rect 20456 23004 21741 23032
rect 14976 22992 14982 23004
rect 19426 22924 19432 22976
rect 19484 22964 19490 22976
rect 19705 22967 19763 22973
rect 19705 22964 19717 22967
rect 19484 22936 19717 22964
rect 19484 22924 19490 22936
rect 19705 22933 19717 22936
rect 19751 22933 19763 22967
rect 19812 22964 19840 23004
rect 21729 23001 21741 23004
rect 21775 23001 21787 23035
rect 24872 23032 24900 23063
rect 24946 23060 24952 23112
rect 25004 23100 25010 23112
rect 25041 23103 25099 23109
rect 25041 23100 25053 23103
rect 25004 23072 25053 23100
rect 25004 23060 25010 23072
rect 25041 23069 25053 23072
rect 25087 23100 25099 23103
rect 25685 23103 25743 23109
rect 25685 23100 25697 23103
rect 25087 23072 25697 23100
rect 25087 23069 25099 23072
rect 25041 23063 25099 23069
rect 25685 23069 25697 23072
rect 25731 23069 25743 23103
rect 25685 23063 25743 23069
rect 26513 23103 26571 23109
rect 26513 23069 26525 23103
rect 26559 23069 26571 23103
rect 26513 23063 26571 23069
rect 26697 23103 26755 23109
rect 26697 23069 26709 23103
rect 26743 23100 26755 23103
rect 27341 23103 27399 23109
rect 27341 23100 27353 23103
rect 26743 23072 27353 23100
rect 26743 23069 26755 23072
rect 26697 23063 26755 23069
rect 27341 23069 27353 23072
rect 27387 23069 27399 23103
rect 27341 23063 27399 23069
rect 25222 23032 25228 23044
rect 24872 23004 25228 23032
rect 21729 22995 21787 23001
rect 25222 22992 25228 23004
rect 25280 23032 25286 23044
rect 25501 23035 25559 23041
rect 25501 23032 25513 23035
rect 25280 23004 25513 23032
rect 25280 22992 25286 23004
rect 25501 23001 25513 23004
rect 25547 23001 25559 23035
rect 25501 22995 25559 23001
rect 25869 23035 25927 23041
rect 25869 23001 25881 23035
rect 25915 23032 25927 23035
rect 26528 23032 26556 23063
rect 28258 23060 28264 23112
rect 28316 23100 28322 23112
rect 28537 23103 28595 23109
rect 28537 23100 28549 23103
rect 28316 23072 28549 23100
rect 28316 23060 28322 23072
rect 28537 23069 28549 23072
rect 28583 23069 28595 23103
rect 30098 23100 30104 23112
rect 30059 23072 30104 23100
rect 28537 23063 28595 23069
rect 30098 23060 30104 23072
rect 30156 23060 30162 23112
rect 33870 23100 33876 23112
rect 33831 23072 33876 23100
rect 33870 23060 33876 23072
rect 33928 23060 33934 23112
rect 34057 23103 34115 23109
rect 34057 23069 34069 23103
rect 34103 23100 34115 23103
rect 34146 23100 34152 23112
rect 34103 23072 34152 23100
rect 34103 23069 34115 23072
rect 34057 23063 34115 23069
rect 34146 23060 34152 23072
rect 34204 23060 34210 23112
rect 34238 23060 34244 23112
rect 34296 23100 34302 23112
rect 34698 23100 34704 23112
rect 34296 23072 34704 23100
rect 34296 23060 34302 23072
rect 34698 23060 34704 23072
rect 34756 23060 34762 23112
rect 40034 23100 40040 23112
rect 39995 23072 40040 23100
rect 40034 23060 40040 23072
rect 40092 23060 40098 23112
rect 42904 23109 42932 23140
rect 43438 23128 43444 23140
rect 43496 23168 43502 23180
rect 43824 23168 43852 23276
rect 47762 23264 47768 23276
rect 47820 23264 47826 23316
rect 47026 23236 47032 23248
rect 43496 23140 43852 23168
rect 43496 23128 43502 23140
rect 42889 23103 42947 23109
rect 42889 23069 42901 23103
rect 42935 23069 42947 23103
rect 42889 23063 42947 23069
rect 42981 23103 43039 23109
rect 42981 23069 42993 23103
rect 43027 23100 43039 23103
rect 43530 23100 43536 23112
rect 43027 23072 43536 23100
rect 43027 23069 43039 23072
rect 42981 23063 43039 23069
rect 43530 23060 43536 23072
rect 43588 23100 43594 23112
rect 43824 23109 43852 23140
rect 45848 23208 47032 23236
rect 45848 23109 45876 23208
rect 47026 23196 47032 23208
rect 47084 23196 47090 23248
rect 46290 23168 46296 23180
rect 46251 23140 46296 23168
rect 46290 23128 46296 23140
rect 46348 23128 46354 23180
rect 46477 23171 46535 23177
rect 46477 23137 46489 23171
rect 46523 23168 46535 23171
rect 47670 23168 47676 23180
rect 46523 23140 47676 23168
rect 46523 23137 46535 23140
rect 46477 23131 46535 23137
rect 47670 23128 47676 23140
rect 47728 23128 47734 23180
rect 48133 23171 48191 23177
rect 48133 23137 48145 23171
rect 48179 23168 48191 23171
rect 48222 23168 48228 23180
rect 48179 23140 48228 23168
rect 48179 23137 48191 23140
rect 48133 23131 48191 23137
rect 48222 23128 48228 23140
rect 48280 23128 48286 23180
rect 43625 23103 43683 23109
rect 43625 23100 43637 23103
rect 43588 23072 43637 23100
rect 43588 23060 43594 23072
rect 43625 23069 43637 23072
rect 43671 23069 43683 23103
rect 43625 23063 43683 23069
rect 43809 23103 43867 23109
rect 43809 23069 43821 23103
rect 43855 23069 43867 23103
rect 43809 23063 43867 23069
rect 45833 23103 45891 23109
rect 45833 23069 45845 23103
rect 45879 23069 45891 23103
rect 45833 23063 45891 23069
rect 25915 23004 26556 23032
rect 25915 23001 25927 23004
rect 25869 22995 25927 23001
rect 28442 22992 28448 23044
rect 28500 23032 28506 23044
rect 31570 23032 31576 23044
rect 28500 23004 31576 23032
rect 28500 22992 28506 23004
rect 31570 22992 31576 23004
rect 31628 22992 31634 23044
rect 32306 22992 32312 23044
rect 32364 22992 32370 23044
rect 40681 23035 40739 23041
rect 40681 23001 40693 23035
rect 40727 23001 40739 23035
rect 40681 22995 40739 23001
rect 42337 23035 42395 23041
rect 42337 23001 42349 23035
rect 42383 23032 42395 23035
rect 45738 23032 45744 23044
rect 42383 23004 45744 23032
rect 42383 23001 42395 23004
rect 42337 22995 42395 23001
rect 25590 22964 25596 22976
rect 19812 22936 25596 22964
rect 19705 22927 19763 22933
rect 25590 22924 25596 22936
rect 25648 22964 25654 22976
rect 27338 22964 27344 22976
rect 25648 22936 27344 22964
rect 25648 22924 25654 22936
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 31938 22924 31944 22976
rect 31996 22964 32002 22976
rect 32214 22964 32220 22976
rect 31996 22936 32220 22964
rect 31996 22924 32002 22936
rect 32214 22924 32220 22936
rect 32272 22924 32278 22976
rect 39853 22967 39911 22973
rect 39853 22933 39865 22967
rect 39899 22964 39911 22967
rect 40696 22964 40724 22995
rect 45738 22992 45744 23004
rect 45796 22992 45802 23044
rect 43714 22964 43720 22976
rect 39899 22936 40724 22964
rect 43675 22936 43720 22964
rect 39899 22933 39911 22936
rect 39853 22927 39911 22933
rect 43714 22924 43720 22936
rect 43772 22924 43778 22976
rect 45370 22924 45376 22976
rect 45428 22964 45434 22976
rect 45649 22967 45707 22973
rect 45649 22964 45661 22967
rect 45428 22936 45661 22964
rect 45428 22924 45434 22936
rect 45649 22933 45661 22936
rect 45695 22933 45707 22967
rect 45649 22927 45707 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 13078 22760 13084 22772
rect 13039 22732 13084 22760
rect 13078 22720 13084 22732
rect 13136 22720 13142 22772
rect 22830 22760 22836 22772
rect 22791 22732 22836 22760
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 28258 22720 28264 22772
rect 28316 22760 28322 22772
rect 30469 22763 30527 22769
rect 30469 22760 30481 22763
rect 28316 22732 30481 22760
rect 28316 22720 28322 22732
rect 30469 22729 30481 22732
rect 30515 22760 30527 22763
rect 30926 22760 30932 22772
rect 30515 22732 30932 22760
rect 30515 22729 30527 22732
rect 30469 22723 30527 22729
rect 30926 22720 30932 22732
rect 30984 22720 30990 22772
rect 32217 22763 32275 22769
rect 32217 22729 32229 22763
rect 32263 22760 32275 22763
rect 32306 22760 32312 22772
rect 32263 22732 32312 22760
rect 32263 22729 32275 22732
rect 32217 22723 32275 22729
rect 32306 22720 32312 22732
rect 32364 22720 32370 22772
rect 40034 22720 40040 22772
rect 40092 22760 40098 22772
rect 40681 22763 40739 22769
rect 40681 22760 40693 22763
rect 40092 22732 40693 22760
rect 40092 22720 40098 22732
rect 40681 22729 40693 22732
rect 40727 22729 40739 22763
rect 42978 22760 42984 22772
rect 40681 22723 40739 22729
rect 42536 22732 42984 22760
rect 13538 22692 13544 22704
rect 11716 22664 13544 22692
rect 11716 22633 11744 22664
rect 13538 22652 13544 22664
rect 13596 22652 13602 22704
rect 21358 22652 21364 22704
rect 21416 22692 21422 22704
rect 28442 22692 28448 22704
rect 21416 22664 28448 22692
rect 21416 22652 21422 22664
rect 28442 22652 28448 22664
rect 28500 22652 28506 22704
rect 28994 22692 29000 22704
rect 28955 22664 29000 22692
rect 28994 22652 29000 22664
rect 29052 22652 29058 22704
rect 29730 22652 29736 22704
rect 29788 22652 29794 22704
rect 34698 22692 34704 22704
rect 31726 22664 34704 22692
rect 11701 22627 11759 22633
rect 11701 22593 11713 22627
rect 11747 22593 11759 22627
rect 11974 22624 11980 22636
rect 11701 22587 11759 22593
rect 11808 22596 11980 22624
rect 11808 22565 11836 22596
rect 11974 22584 11980 22596
rect 12032 22624 12038 22636
rect 12342 22624 12348 22636
rect 12032 22596 12348 22624
rect 12032 22584 12038 22596
rect 12342 22584 12348 22596
rect 12400 22584 12406 22636
rect 12986 22624 12992 22636
rect 12947 22596 12992 22624
rect 12986 22584 12992 22596
rect 13044 22584 13050 22636
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22624 15163 22627
rect 18230 22624 18236 22636
rect 15151 22596 18236 22624
rect 15151 22593 15163 22596
rect 15105 22587 15163 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 22738 22624 22744 22636
rect 22699 22596 22744 22624
rect 22738 22584 22744 22596
rect 22796 22584 22802 22636
rect 25590 22624 25596 22636
rect 25551 22596 25596 22624
rect 25590 22584 25596 22596
rect 25648 22584 25654 22636
rect 27338 22584 27344 22636
rect 27396 22624 27402 22636
rect 27893 22627 27951 22633
rect 27893 22624 27905 22627
rect 27396 22596 27905 22624
rect 27396 22584 27402 22596
rect 27893 22593 27905 22596
rect 27939 22593 27951 22627
rect 30650 22624 30656 22636
rect 27893 22587 27951 22593
rect 30392 22596 30656 22624
rect 11793 22559 11851 22565
rect 11793 22525 11805 22559
rect 11839 22525 11851 22559
rect 12066 22556 12072 22568
rect 12027 22528 12072 22556
rect 11793 22519 11851 22525
rect 12066 22516 12072 22528
rect 12124 22516 12130 22568
rect 28721 22559 28779 22565
rect 28721 22525 28733 22559
rect 28767 22556 28779 22559
rect 29546 22556 29552 22568
rect 28767 22528 29552 22556
rect 28767 22525 28779 22528
rect 28721 22519 28779 22525
rect 29546 22516 29552 22528
rect 29604 22516 29610 22568
rect 15194 22420 15200 22432
rect 15155 22392 15200 22420
rect 15194 22380 15200 22392
rect 15252 22380 15258 22432
rect 25409 22423 25467 22429
rect 25409 22389 25421 22423
rect 25455 22420 25467 22423
rect 25682 22420 25688 22432
rect 25455 22392 25688 22420
rect 25455 22389 25467 22392
rect 25409 22383 25467 22389
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 28077 22423 28135 22429
rect 28077 22389 28089 22423
rect 28123 22420 28135 22423
rect 30190 22420 30196 22432
rect 28123 22392 30196 22420
rect 28123 22389 28135 22392
rect 28077 22383 28135 22389
rect 30190 22380 30196 22392
rect 30248 22420 30254 22432
rect 30392 22420 30420 22596
rect 30650 22584 30656 22596
rect 30708 22624 30714 22636
rect 31113 22627 31171 22633
rect 31113 22624 31125 22627
rect 30708 22596 31125 22624
rect 30708 22584 30714 22596
rect 31113 22593 31125 22596
rect 31159 22624 31171 22627
rect 31726 22624 31754 22664
rect 34698 22652 34704 22664
rect 34756 22652 34762 22704
rect 42536 22701 42564 22732
rect 42978 22720 42984 22732
rect 43036 22760 43042 22772
rect 43714 22760 43720 22772
rect 43036 22732 43720 22760
rect 43036 22720 43042 22732
rect 43714 22720 43720 22732
rect 43772 22720 43778 22772
rect 42521 22695 42579 22701
rect 42521 22661 42533 22695
rect 42567 22661 42579 22695
rect 42521 22655 42579 22661
rect 42705 22695 42763 22701
rect 42705 22661 42717 22695
rect 42751 22692 42763 22695
rect 43349 22695 43407 22701
rect 43349 22692 43361 22695
rect 42751 22664 43361 22692
rect 42751 22661 42763 22664
rect 42705 22655 42763 22661
rect 43349 22661 43361 22664
rect 43395 22661 43407 22695
rect 45370 22692 45376 22704
rect 45331 22664 45376 22692
rect 43349 22655 43407 22661
rect 45370 22652 45376 22664
rect 45428 22652 45434 22704
rect 31159 22596 31754 22624
rect 31159 22593 31171 22596
rect 31113 22587 31171 22593
rect 32030 22584 32036 22636
rect 32088 22624 32094 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 32088 22596 32137 22624
rect 32088 22584 32094 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 40221 22627 40279 22633
rect 40221 22593 40233 22627
rect 40267 22624 40279 22627
rect 40310 22624 40316 22636
rect 40267 22596 40316 22624
rect 40267 22593 40279 22596
rect 40221 22587 40279 22593
rect 40310 22584 40316 22596
rect 40368 22584 40374 22636
rect 42794 22624 42800 22636
rect 42755 22596 42800 22624
rect 42794 22584 42800 22596
rect 42852 22584 42858 22636
rect 43257 22627 43315 22633
rect 43257 22593 43269 22627
rect 43303 22593 43315 22627
rect 43438 22624 43444 22636
rect 43399 22596 43444 22624
rect 43257 22587 43315 22593
rect 43272 22556 43300 22587
rect 43438 22584 43444 22596
rect 43496 22584 43502 22636
rect 44729 22627 44787 22633
rect 44729 22593 44741 22627
rect 44775 22593 44787 22627
rect 45186 22624 45192 22636
rect 45147 22596 45192 22624
rect 44729 22587 44787 22593
rect 43530 22556 43536 22568
rect 43272 22528 43536 22556
rect 43530 22516 43536 22528
rect 43588 22516 43594 22568
rect 42518 22488 42524 22500
rect 42479 22460 42524 22488
rect 42518 22448 42524 22460
rect 42576 22448 42582 22500
rect 44744 22488 44772 22587
rect 45186 22584 45192 22596
rect 45244 22584 45250 22636
rect 47578 22624 47584 22636
rect 47539 22596 47584 22624
rect 47578 22584 47584 22596
rect 47636 22624 47642 22636
rect 47946 22624 47952 22636
rect 47636 22596 47952 22624
rect 47636 22584 47642 22596
rect 47946 22584 47952 22596
rect 48004 22584 48010 22636
rect 45738 22556 45744 22568
rect 45699 22528 45744 22556
rect 45738 22516 45744 22528
rect 45796 22516 45802 22568
rect 47670 22516 47676 22568
rect 47728 22556 47734 22568
rect 47857 22559 47915 22565
rect 47857 22556 47869 22559
rect 47728 22528 47869 22556
rect 47728 22516 47734 22528
rect 47857 22525 47869 22528
rect 47903 22525 47915 22559
rect 47857 22519 47915 22525
rect 48133 22491 48191 22497
rect 48133 22488 48145 22491
rect 44744 22460 48145 22488
rect 48133 22457 48145 22460
rect 48179 22457 48191 22491
rect 48133 22451 48191 22457
rect 31294 22420 31300 22432
rect 30248 22392 30420 22420
rect 31255 22392 31300 22420
rect 30248 22380 30254 22392
rect 31294 22380 31300 22392
rect 31352 22380 31358 22432
rect 40126 22380 40132 22432
rect 40184 22420 40190 22432
rect 40313 22423 40371 22429
rect 40313 22420 40325 22423
rect 40184 22392 40325 22420
rect 40184 22380 40190 22392
rect 40313 22389 40325 22392
rect 40359 22389 40371 22423
rect 40313 22383 40371 22389
rect 44545 22423 44603 22429
rect 44545 22389 44557 22423
rect 44591 22420 44603 22423
rect 45370 22420 45376 22432
rect 44591 22392 45376 22420
rect 44591 22389 44603 22392
rect 44545 22383 44603 22389
rect 45370 22380 45376 22392
rect 45428 22380 45434 22432
rect 47486 22380 47492 22432
rect 47544 22420 47550 22432
rect 47673 22423 47731 22429
rect 47673 22420 47685 22423
rect 47544 22392 47685 22420
rect 47544 22380 47550 22392
rect 47673 22389 47685 22392
rect 47719 22389 47731 22423
rect 47673 22383 47731 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 25590 22176 25596 22228
rect 25648 22216 25654 22228
rect 26145 22219 26203 22225
rect 26145 22216 26157 22219
rect 25648 22188 26157 22216
rect 25648 22176 25654 22188
rect 26145 22185 26157 22188
rect 26191 22185 26203 22219
rect 29546 22216 29552 22228
rect 29507 22188 29552 22216
rect 26145 22179 26203 22185
rect 29546 22176 29552 22188
rect 29604 22176 29610 22228
rect 35069 22219 35127 22225
rect 35069 22185 35081 22219
rect 35115 22216 35127 22219
rect 35434 22216 35440 22228
rect 35115 22188 35440 22216
rect 35115 22185 35127 22188
rect 35069 22179 35127 22185
rect 35434 22176 35440 22188
rect 35492 22216 35498 22228
rect 35529 22219 35587 22225
rect 35529 22216 35541 22219
rect 35492 22188 35541 22216
rect 35492 22176 35498 22188
rect 35529 22185 35541 22188
rect 35575 22185 35587 22219
rect 35529 22179 35587 22185
rect 13173 22151 13231 22157
rect 13173 22117 13185 22151
rect 13219 22148 13231 22151
rect 25958 22148 25964 22160
rect 13219 22120 13253 22148
rect 25919 22120 25964 22148
rect 13219 22117 13231 22120
rect 13173 22111 13231 22117
rect 14 22040 20 22092
rect 72 22080 78 22092
rect 13188 22080 13216 22111
rect 25958 22108 25964 22120
rect 26016 22108 26022 22160
rect 26694 22148 26700 22160
rect 26655 22120 26700 22148
rect 26694 22108 26700 22120
rect 26752 22108 26758 22160
rect 30837 22151 30895 22157
rect 30837 22117 30849 22151
rect 30883 22148 30895 22151
rect 30883 22120 31432 22148
rect 30883 22117 30895 22120
rect 30837 22111 30895 22117
rect 14826 22080 14832 22092
rect 72 22052 6914 22080
rect 72 22040 78 22052
rect 6886 21944 6914 22052
rect 11900 22052 13216 22080
rect 14787 22052 14832 22080
rect 11900 22024 11928 22052
rect 14826 22040 14832 22052
rect 14884 22040 14890 22092
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22080 15071 22083
rect 15194 22080 15200 22092
rect 15059 22052 15200 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 19978 22080 19984 22092
rect 15344 22052 15389 22080
rect 18524 22052 19984 22080
rect 15344 22040 15350 22052
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 11882 22012 11888 22024
rect 11839 21984 11888 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 12342 22012 12348 22024
rect 12303 21984 12348 22012
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12492 21984 12541 22012
rect 12492 21972 12498 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 12989 22015 13047 22021
rect 12989 21981 13001 22015
rect 13035 22012 13047 22015
rect 14734 22012 14740 22024
rect 13035 21984 14740 22012
rect 13035 21981 13047 21984
rect 12989 21975 13047 21981
rect 14734 21972 14740 21984
rect 14792 21972 14798 22024
rect 16298 21972 16304 22024
rect 16356 22012 16362 22024
rect 18524 22021 18552 22052
rect 19978 22040 19984 22052
rect 20036 22040 20042 22092
rect 23382 22040 23388 22092
rect 23440 22080 23446 22092
rect 24397 22083 24455 22089
rect 24397 22080 24409 22083
rect 23440 22052 24409 22080
rect 23440 22040 23446 22052
rect 24397 22049 24409 22052
rect 24443 22080 24455 22083
rect 27982 22080 27988 22092
rect 24443 22052 27988 22080
rect 24443 22049 24455 22052
rect 24397 22043 24455 22049
rect 27982 22040 27988 22052
rect 28040 22040 28046 22092
rect 30558 22080 30564 22092
rect 30519 22052 30564 22080
rect 30558 22040 30564 22052
rect 30616 22040 30622 22092
rect 31294 22080 31300 22092
rect 31255 22052 31300 22080
rect 31294 22040 31300 22052
rect 31352 22040 31358 22092
rect 31404 22080 31432 22120
rect 31573 22083 31631 22089
rect 31573 22080 31585 22083
rect 31404 22052 31585 22080
rect 31573 22049 31585 22052
rect 31619 22049 31631 22083
rect 31573 22043 31631 22049
rect 31662 22040 31668 22092
rect 31720 22080 31726 22092
rect 31938 22080 31944 22092
rect 31720 22052 31944 22080
rect 31720 22040 31726 22052
rect 31938 22040 31944 22052
rect 31996 22080 32002 22092
rect 37274 22080 37280 22092
rect 31996 22052 37280 22080
rect 31996 22040 32002 22052
rect 37274 22040 37280 22052
rect 37332 22040 37338 22092
rect 40126 22040 40132 22092
rect 40184 22080 40190 22092
rect 40184 22052 40448 22080
rect 40184 22040 40190 22052
rect 17129 22015 17187 22021
rect 17129 22012 17141 22015
rect 16356 21984 17141 22012
rect 16356 21972 16362 21984
rect 17129 21981 17141 21984
rect 17175 21981 17187 22015
rect 18509 22015 18567 22021
rect 18509 22012 18521 22015
rect 17129 21975 17187 21981
rect 18156 21984 18521 22012
rect 16574 21944 16580 21956
rect 6886 21916 16580 21944
rect 16574 21904 16580 21916
rect 16632 21904 16638 21956
rect 18156 21944 18184 21984
rect 18509 21981 18521 21984
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 19245 22015 19303 22021
rect 19245 21981 19257 22015
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 20349 22015 20407 22021
rect 20349 21981 20361 22015
rect 20395 22012 20407 22015
rect 22186 22012 22192 22024
rect 20395 21984 22192 22012
rect 20395 21981 20407 21984
rect 20349 21975 20407 21981
rect 16776 21916 18184 21944
rect 11514 21836 11520 21888
rect 11572 21876 11578 21888
rect 11793 21879 11851 21885
rect 11793 21876 11805 21879
rect 11572 21848 11805 21876
rect 11572 21836 11578 21848
rect 11793 21845 11805 21848
rect 11839 21845 11851 21879
rect 11793 21839 11851 21845
rect 11882 21836 11888 21888
rect 11940 21876 11946 21888
rect 12437 21879 12495 21885
rect 12437 21876 12449 21879
rect 11940 21848 12449 21876
rect 11940 21836 11946 21848
rect 12437 21845 12449 21848
rect 12483 21845 12495 21879
rect 12437 21839 12495 21845
rect 16390 21836 16396 21888
rect 16448 21876 16454 21888
rect 16776 21876 16804 21916
rect 18230 21904 18236 21956
rect 18288 21944 18294 21956
rect 19260 21944 19288 21975
rect 22186 21972 22192 21984
rect 22244 22012 22250 22024
rect 22465 22015 22523 22021
rect 22465 22012 22477 22015
rect 22244 21984 22477 22012
rect 22244 21972 22250 21984
rect 22465 21981 22477 21984
rect 22511 22012 22523 22015
rect 24673 22015 24731 22021
rect 22511 21984 24624 22012
rect 22511 21981 22523 21984
rect 22465 21975 22523 21981
rect 18288 21916 19288 21944
rect 18288 21904 18294 21916
rect 20622 21904 20628 21956
rect 20680 21944 20686 21956
rect 20898 21944 20904 21956
rect 20680 21916 20904 21944
rect 20680 21904 20686 21916
rect 20898 21904 20904 21916
rect 20956 21904 20962 21956
rect 22738 21904 22744 21956
rect 22796 21944 22802 21956
rect 22833 21947 22891 21953
rect 22833 21944 22845 21947
rect 22796 21916 22845 21944
rect 22796 21904 22802 21916
rect 22833 21913 22845 21916
rect 22879 21913 22891 21947
rect 22833 21907 22891 21913
rect 16448 21848 16804 21876
rect 16448 21836 16454 21848
rect 16850 21836 16856 21888
rect 16908 21876 16914 21888
rect 17221 21879 17279 21885
rect 17221 21876 17233 21879
rect 16908 21848 17233 21876
rect 16908 21836 16914 21848
rect 17221 21845 17233 21848
rect 17267 21845 17279 21879
rect 18598 21876 18604 21888
rect 18559 21848 18604 21876
rect 17221 21839 17279 21845
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 19334 21876 19340 21888
rect 19295 21848 19340 21876
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 24596 21876 24624 21984
rect 24673 21981 24685 22015
rect 24719 22012 24731 22015
rect 24946 22012 24952 22024
rect 24719 21984 24952 22012
rect 24719 21981 24731 21984
rect 24673 21975 24731 21981
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 26418 21972 26424 22024
rect 26476 22012 26482 22024
rect 26605 22015 26663 22021
rect 26605 22012 26617 22015
rect 26476 21984 26617 22012
rect 26476 21972 26482 21984
rect 26605 21981 26617 21984
rect 26651 21981 26663 22015
rect 26605 21975 26663 21981
rect 28353 22015 28411 22021
rect 28353 21981 28365 22015
rect 28399 22012 28411 22015
rect 29638 22012 29644 22024
rect 28399 21984 29644 22012
rect 28399 21981 28411 21984
rect 28353 21975 28411 21981
rect 25130 21904 25136 21956
rect 25188 21944 25194 21956
rect 25685 21947 25743 21953
rect 25685 21944 25697 21947
rect 25188 21916 25697 21944
rect 25188 21904 25194 21916
rect 25685 21913 25697 21916
rect 25731 21913 25743 21947
rect 25685 21907 25743 21913
rect 28368 21876 28396 21975
rect 29638 21972 29644 21984
rect 29696 21972 29702 22024
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 22012 29791 22015
rect 30190 22012 30196 22024
rect 29779 21984 30196 22012
rect 29779 21981 29791 21984
rect 29733 21975 29791 21981
rect 30190 21972 30196 21984
rect 30248 21972 30254 22024
rect 30466 22012 30472 22024
rect 30427 21984 30472 22012
rect 30466 21972 30472 21984
rect 30524 21972 30530 22024
rect 34793 22015 34851 22021
rect 34793 21981 34805 22015
rect 34839 22012 34851 22015
rect 35894 22012 35900 22024
rect 34839 21984 35900 22012
rect 34839 21981 34851 21984
rect 34793 21975 34851 21981
rect 35894 21972 35900 21984
rect 35952 21972 35958 22024
rect 40310 22012 40316 22024
rect 40271 21984 40316 22012
rect 40310 21972 40316 21984
rect 40368 21972 40374 22024
rect 40420 22021 40448 22052
rect 44634 22040 44640 22092
rect 44692 22080 44698 22092
rect 45189 22083 45247 22089
rect 45189 22080 45201 22083
rect 44692 22052 45201 22080
rect 44692 22040 44698 22052
rect 45189 22049 45201 22052
rect 45235 22049 45247 22083
rect 45370 22080 45376 22092
rect 45331 22052 45376 22080
rect 45189 22043 45247 22049
rect 45370 22040 45376 22052
rect 45428 22040 45434 22092
rect 45738 22080 45744 22092
rect 45699 22052 45744 22080
rect 45738 22040 45744 22052
rect 45796 22040 45802 22092
rect 47489 22083 47547 22089
rect 47489 22049 47501 22083
rect 47535 22080 47547 22083
rect 47854 22080 47860 22092
rect 47535 22052 47860 22080
rect 47535 22049 47547 22052
rect 47489 22043 47547 22049
rect 47854 22040 47860 22052
rect 47912 22040 47918 22092
rect 40405 22015 40463 22021
rect 40405 21981 40417 22015
rect 40451 21981 40463 22015
rect 40405 21975 40463 21981
rect 40494 21972 40500 22024
rect 40552 22012 40558 22024
rect 40552 21984 41414 22012
rect 40552 21972 40558 21984
rect 28534 21904 28540 21956
rect 28592 21944 28598 21956
rect 28629 21947 28687 21953
rect 28629 21944 28641 21947
rect 28592 21916 28641 21944
rect 28592 21904 28598 21916
rect 28629 21913 28641 21916
rect 28675 21944 28687 21947
rect 31662 21944 31668 21956
rect 28675 21916 31668 21944
rect 28675 21913 28687 21916
rect 28629 21907 28687 21913
rect 31662 21904 31668 21916
rect 31720 21904 31726 21956
rect 32214 21904 32220 21956
rect 32272 21904 32278 21956
rect 40589 21947 40647 21953
rect 40589 21944 40601 21947
rect 40420 21916 40601 21944
rect 40420 21888 40448 21916
rect 40589 21913 40601 21916
rect 40635 21913 40647 21947
rect 41386 21944 41414 21984
rect 43254 21972 43260 22024
rect 43312 22012 43318 22024
rect 43349 22015 43407 22021
rect 43349 22012 43361 22015
rect 43312 21984 43361 22012
rect 43312 21972 43318 21984
rect 43349 21981 43361 21984
rect 43395 21981 43407 22015
rect 43349 21975 43407 21981
rect 43438 21972 43444 22024
rect 43496 22012 43502 22024
rect 43533 22015 43591 22021
rect 43533 22012 43545 22015
rect 43496 21984 43545 22012
rect 43496 21972 43502 21984
rect 43533 21981 43545 21984
rect 43579 22012 43591 22015
rect 44177 22015 44235 22021
rect 44177 22012 44189 22015
rect 43579 21984 44189 22012
rect 43579 21981 43591 21984
rect 43533 21975 43591 21981
rect 44177 21981 44189 21984
rect 44223 21981 44235 22015
rect 44177 21975 44235 21981
rect 44361 22015 44419 22021
rect 44361 21981 44373 22015
rect 44407 22012 44419 22015
rect 45094 22012 45100 22024
rect 44407 21984 45100 22012
rect 44407 21981 44419 21984
rect 44361 21975 44419 21981
rect 45094 21972 45100 21984
rect 45152 21972 45158 22024
rect 47673 22015 47731 22021
rect 47673 21981 47685 22015
rect 47719 22012 47731 22015
rect 47762 22012 47768 22024
rect 47719 21984 47768 22012
rect 47719 21981 47731 21984
rect 47673 21975 47731 21981
rect 47762 21972 47768 21984
rect 47820 22012 47826 22024
rect 47946 22012 47952 22024
rect 47820 21984 47952 22012
rect 47820 21972 47826 21984
rect 47946 21972 47952 21984
rect 48004 21972 48010 22024
rect 48041 21947 48099 21953
rect 48041 21944 48053 21947
rect 41386 21916 44496 21944
rect 40589 21907 40647 21913
rect 24596 21848 28396 21876
rect 30466 21836 30472 21888
rect 30524 21876 30530 21888
rect 32858 21876 32864 21888
rect 30524 21848 32864 21876
rect 30524 21836 30530 21848
rect 32858 21836 32864 21848
rect 32916 21876 32922 21888
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32916 21848 33057 21876
rect 32916 21836 32922 21848
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 34606 21836 34612 21888
rect 34664 21876 34670 21888
rect 35253 21879 35311 21885
rect 35253 21876 35265 21879
rect 34664 21848 35265 21876
rect 34664 21836 34670 21848
rect 35253 21845 35265 21848
rect 35299 21845 35311 21879
rect 35253 21839 35311 21845
rect 40402 21836 40408 21888
rect 40460 21836 40466 21888
rect 43438 21876 43444 21888
rect 43399 21848 43444 21876
rect 43438 21836 43444 21848
rect 43496 21836 43502 21888
rect 44358 21876 44364 21888
rect 44319 21848 44364 21876
rect 44358 21836 44364 21848
rect 44416 21836 44422 21888
rect 44468 21876 44496 21916
rect 47136 21916 48053 21944
rect 47136 21876 47164 21916
rect 48041 21913 48053 21916
rect 48087 21913 48099 21947
rect 48041 21907 48099 21913
rect 44468 21848 47164 21876
rect 47670 21836 47676 21888
rect 47728 21876 47734 21888
rect 47765 21879 47823 21885
rect 47765 21876 47777 21879
rect 47728 21848 47777 21876
rect 47728 21836 47734 21848
rect 47765 21845 47777 21848
rect 47811 21845 47823 21879
rect 47765 21839 47823 21845
rect 47854 21836 47860 21888
rect 47912 21876 47918 21888
rect 47912 21848 47957 21876
rect 47912 21836 47918 21848
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 3694 21632 3700 21684
rect 3752 21672 3758 21684
rect 18046 21672 18052 21684
rect 3752 21644 10180 21672
rect 3752 21632 3758 21644
rect 3510 21564 3516 21616
rect 3568 21604 3574 21616
rect 3568 21576 6914 21604
rect 3568 21564 3574 21576
rect 6886 21332 6914 21576
rect 10152 21400 10180 21644
rect 10796 21644 11836 21672
rect 10796 21545 10824 21644
rect 11808 21616 11836 21644
rect 16684 21644 18052 21672
rect 10873 21607 10931 21613
rect 10873 21573 10885 21607
rect 10919 21604 10931 21607
rect 11701 21607 11759 21613
rect 11701 21604 11713 21607
rect 10919 21576 11713 21604
rect 10919 21573 10931 21576
rect 10873 21567 10931 21573
rect 11701 21573 11713 21576
rect 11747 21573 11759 21607
rect 11701 21567 11759 21573
rect 11790 21564 11796 21616
rect 11848 21604 11854 21616
rect 16390 21604 16396 21616
rect 11848 21576 16396 21604
rect 11848 21564 11854 21576
rect 16390 21564 16396 21576
rect 16448 21564 16454 21616
rect 16684 21545 16712 21644
rect 18046 21632 18052 21644
rect 18104 21632 18110 21684
rect 19978 21632 19984 21684
rect 20036 21672 20042 21684
rect 20530 21672 20536 21684
rect 20036 21644 20536 21672
rect 20036 21632 20042 21644
rect 20530 21632 20536 21644
rect 20588 21672 20594 21684
rect 22373 21675 22431 21681
rect 22373 21672 22385 21675
rect 20588 21644 22385 21672
rect 20588 21632 20594 21644
rect 22373 21641 22385 21644
rect 22419 21641 22431 21675
rect 22373 21635 22431 21641
rect 25041 21675 25099 21681
rect 25041 21641 25053 21675
rect 25087 21672 25099 21675
rect 25222 21672 25228 21684
rect 25087 21644 25228 21672
rect 25087 21641 25099 21644
rect 25041 21635 25099 21641
rect 25222 21632 25228 21644
rect 25280 21672 25286 21684
rect 25590 21672 25596 21684
rect 25280 21644 25596 21672
rect 25280 21632 25286 21644
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 25685 21675 25743 21681
rect 25685 21641 25697 21675
rect 25731 21672 25743 21675
rect 25958 21672 25964 21684
rect 25731 21644 25964 21672
rect 25731 21641 25743 21644
rect 25685 21635 25743 21641
rect 25958 21632 25964 21644
rect 26016 21632 26022 21684
rect 26970 21632 26976 21684
rect 27028 21672 27034 21684
rect 27525 21675 27583 21681
rect 27525 21672 27537 21675
rect 27028 21644 27537 21672
rect 27028 21632 27034 21644
rect 27525 21641 27537 21644
rect 27571 21672 27583 21675
rect 31202 21672 31208 21684
rect 27571 21644 31208 21672
rect 27571 21641 27583 21644
rect 27525 21635 27583 21641
rect 31202 21632 31208 21644
rect 31260 21632 31266 21684
rect 32214 21672 32220 21684
rect 32175 21644 32220 21672
rect 32214 21632 32220 21644
rect 32272 21632 32278 21684
rect 46106 21672 46112 21684
rect 35176 21644 46112 21672
rect 16850 21604 16856 21616
rect 16811 21576 16856 21604
rect 16850 21564 16856 21576
rect 16908 21564 16914 21616
rect 19334 21564 19340 21616
rect 19392 21604 19398 21616
rect 19613 21607 19671 21613
rect 19613 21604 19625 21607
rect 19392 21576 19625 21604
rect 19392 21564 19398 21576
rect 19613 21573 19625 21576
rect 19659 21573 19671 21607
rect 19613 21567 19671 21573
rect 21269 21607 21327 21613
rect 21269 21573 21281 21607
rect 21315 21604 21327 21607
rect 35176 21604 35204 21644
rect 46106 21632 46112 21644
rect 46164 21632 46170 21684
rect 46934 21632 46940 21684
rect 46992 21672 46998 21684
rect 47854 21672 47860 21684
rect 46992 21644 47860 21672
rect 46992 21632 46998 21644
rect 47854 21632 47860 21644
rect 47912 21632 47918 21684
rect 21315 21576 35204 21604
rect 21315 21573 21327 21576
rect 21269 21567 21327 21573
rect 35250 21564 35256 21616
rect 35308 21604 35314 21616
rect 42797 21607 42855 21613
rect 35308 21576 35353 21604
rect 35308 21564 35314 21576
rect 42797 21573 42809 21607
rect 42843 21604 42855 21607
rect 43070 21604 43076 21616
rect 42843 21576 43076 21604
rect 42843 21573 42855 21576
rect 42797 21567 42855 21573
rect 43070 21564 43076 21576
rect 43128 21564 43134 21616
rect 45186 21604 45192 21616
rect 45147 21576 45192 21604
rect 45186 21564 45192 21576
rect 45244 21564 45250 21616
rect 47578 21604 47584 21616
rect 47539 21576 47584 21604
rect 47578 21564 47584 21576
rect 47636 21564 47642 21616
rect 47762 21604 47768 21616
rect 47723 21576 47768 21604
rect 47762 21564 47768 21576
rect 47820 21564 47826 21616
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22281 21539 22339 21545
rect 22281 21536 22293 21539
rect 22244 21508 22293 21536
rect 22244 21496 22250 21508
rect 22281 21505 22293 21508
rect 22327 21505 22339 21539
rect 23198 21536 23204 21548
rect 23159 21508 23204 21536
rect 22281 21499 22339 21505
rect 23198 21496 23204 21508
rect 23256 21496 23262 21548
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21536 23443 21539
rect 24670 21536 24676 21548
rect 23431 21508 24676 21536
rect 23431 21505 23443 21508
rect 23385 21499 23443 21505
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21468 11575 21471
rect 11698 21468 11704 21480
rect 11563 21440 11704 21468
rect 11563 21437 11575 21440
rect 11517 21431 11575 21437
rect 11698 21428 11704 21440
rect 11756 21428 11762 21480
rect 11977 21471 12035 21477
rect 11977 21437 11989 21471
rect 12023 21437 12035 21471
rect 14274 21468 14280 21480
rect 14235 21440 14280 21468
rect 11977 21431 12035 21437
rect 11992 21400 12020 21431
rect 14274 21428 14280 21440
rect 14332 21428 14338 21480
rect 14458 21468 14464 21480
rect 14419 21440 14464 21468
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 14737 21471 14795 21477
rect 14737 21437 14749 21471
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21437 17187 21471
rect 17129 21431 17187 21437
rect 19429 21471 19487 21477
rect 19429 21437 19441 21471
rect 19475 21468 19487 21471
rect 19978 21468 19984 21480
rect 19475 21440 19984 21468
rect 19475 21437 19487 21440
rect 19429 21431 19487 21437
rect 10152 21372 12020 21400
rect 14752 21332 14780 21431
rect 16574 21360 16580 21412
rect 16632 21400 16638 21412
rect 17144 21400 17172 21431
rect 19978 21428 19984 21440
rect 20036 21428 20042 21480
rect 21634 21428 21640 21480
rect 21692 21468 21698 21480
rect 23400 21468 23428 21499
rect 24670 21496 24676 21508
rect 24728 21496 24734 21548
rect 24854 21536 24860 21548
rect 24815 21508 24860 21536
rect 24854 21496 24860 21508
rect 24912 21496 24918 21548
rect 24946 21496 24952 21548
rect 25004 21536 25010 21548
rect 25004 21508 25049 21536
rect 25004 21496 25010 21508
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 25225 21539 25283 21545
rect 25225 21536 25237 21539
rect 25188 21508 25237 21536
rect 25188 21496 25194 21508
rect 25225 21505 25237 21508
rect 25271 21505 25283 21539
rect 25225 21499 25283 21505
rect 25590 21496 25596 21548
rect 25648 21536 25654 21548
rect 25869 21539 25927 21545
rect 25869 21536 25881 21539
rect 25648 21508 25881 21536
rect 25648 21496 25654 21508
rect 25869 21505 25881 21508
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 26145 21539 26203 21545
rect 26145 21505 26157 21539
rect 26191 21536 26203 21539
rect 27338 21536 27344 21548
rect 26191 21508 26280 21536
rect 27299 21508 27344 21536
rect 26191 21505 26203 21508
rect 26145 21499 26203 21505
rect 21692 21440 23428 21468
rect 24964 21468 24992 21496
rect 25961 21471 26019 21477
rect 25961 21468 25973 21471
rect 24964 21440 25973 21468
rect 21692 21428 21698 21440
rect 25961 21437 25973 21440
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 26050 21428 26056 21480
rect 26108 21468 26114 21480
rect 26108 21440 26201 21468
rect 26108 21428 26114 21440
rect 16632 21372 17172 21400
rect 16632 21360 16638 21372
rect 22738 21360 22744 21412
rect 22796 21400 22802 21412
rect 22796 21372 24348 21400
rect 22796 21360 22802 21372
rect 6886 21304 14780 21332
rect 24320 21332 24348 21372
rect 24394 21360 24400 21412
rect 24452 21400 24458 21412
rect 24673 21403 24731 21409
rect 24673 21400 24685 21403
rect 24452 21372 24685 21400
rect 24452 21360 24458 21372
rect 24673 21369 24685 21372
rect 24719 21369 24731 21403
rect 24673 21363 24731 21369
rect 24578 21332 24584 21344
rect 24320 21304 24584 21332
rect 24578 21292 24584 21304
rect 24636 21292 24642 21344
rect 24688 21332 24716 21363
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 26068 21400 26096 21428
rect 24912 21372 26096 21400
rect 24912 21360 24918 21372
rect 26252 21332 26280 21508
rect 27338 21496 27344 21508
rect 27396 21496 27402 21548
rect 28258 21536 28264 21548
rect 28219 21508 28264 21536
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 29638 21496 29644 21548
rect 29696 21536 29702 21548
rect 30653 21539 30711 21545
rect 30653 21536 30665 21539
rect 29696 21508 30665 21536
rect 29696 21496 29702 21508
rect 30653 21505 30665 21508
rect 30699 21505 30711 21539
rect 30653 21499 30711 21505
rect 32030 21496 32036 21548
rect 32088 21536 32094 21548
rect 32125 21539 32183 21545
rect 32125 21536 32137 21539
rect 32088 21508 32137 21536
rect 32088 21496 32094 21508
rect 32125 21505 32137 21508
rect 32171 21505 32183 21539
rect 34606 21536 34612 21548
rect 34567 21508 34612 21536
rect 32125 21499 32183 21505
rect 34606 21496 34612 21508
rect 34664 21496 34670 21548
rect 42886 21496 42892 21548
rect 42944 21536 42950 21548
rect 42981 21539 43039 21545
rect 42981 21536 42993 21539
rect 42944 21508 42993 21536
rect 42944 21496 42950 21508
rect 42981 21505 42993 21508
rect 43027 21505 43039 21539
rect 42981 21499 43039 21505
rect 43901 21539 43959 21545
rect 43901 21505 43913 21539
rect 43947 21505 43959 21539
rect 43901 21499 43959 21505
rect 28445 21471 28503 21477
rect 28445 21437 28457 21471
rect 28491 21468 28503 21471
rect 28626 21468 28632 21480
rect 28491 21440 28632 21468
rect 28491 21437 28503 21440
rect 28445 21431 28503 21437
rect 28626 21428 28632 21440
rect 28684 21428 28690 21480
rect 28994 21468 29000 21480
rect 28955 21440 29000 21468
rect 28994 21428 29000 21440
rect 29052 21428 29058 21480
rect 31481 21471 31539 21477
rect 31481 21437 31493 21471
rect 31527 21468 31539 21471
rect 32950 21468 32956 21480
rect 31527 21440 32956 21468
rect 31527 21437 31539 21440
rect 31481 21431 31539 21437
rect 32950 21428 32956 21440
rect 33008 21428 33014 21480
rect 35161 21471 35219 21477
rect 35161 21468 35173 21471
rect 33428 21440 35173 21468
rect 27154 21332 27160 21344
rect 24688 21304 27160 21332
rect 27154 21292 27160 21304
rect 27212 21292 27218 21344
rect 27706 21292 27712 21344
rect 27764 21332 27770 21344
rect 33428 21332 33456 21440
rect 35161 21437 35173 21440
rect 35207 21437 35219 21471
rect 36170 21468 36176 21480
rect 36131 21440 36176 21468
rect 35161 21431 35219 21437
rect 36170 21428 36176 21440
rect 36228 21428 36234 21480
rect 34425 21403 34483 21409
rect 34425 21369 34437 21403
rect 34471 21400 34483 21403
rect 35250 21400 35256 21412
rect 34471 21372 35256 21400
rect 34471 21369 34483 21372
rect 34425 21363 34483 21369
rect 35250 21360 35256 21372
rect 35308 21360 35314 21412
rect 43916 21400 43944 21499
rect 44358 21496 44364 21548
rect 44416 21536 44422 21548
rect 46198 21536 46204 21548
rect 44416 21508 44574 21536
rect 46159 21508 46204 21536
rect 44416 21496 44422 21508
rect 46198 21496 46204 21508
rect 46256 21496 46262 21548
rect 44634 21468 44640 21480
rect 44595 21440 44640 21468
rect 44634 21428 44640 21440
rect 44692 21428 44698 21480
rect 45646 21428 45652 21480
rect 45704 21468 45710 21480
rect 46477 21471 46535 21477
rect 46477 21468 46489 21471
rect 45704 21440 46489 21468
rect 45704 21428 45710 21440
rect 46477 21437 46489 21440
rect 46523 21437 46535 21471
rect 46477 21431 46535 21437
rect 47949 21403 48007 21409
rect 47949 21400 47961 21403
rect 43916 21372 47961 21400
rect 47949 21369 47961 21372
rect 47995 21369 48007 21403
rect 47949 21363 48007 21369
rect 43162 21332 43168 21344
rect 27764 21304 33456 21332
rect 43123 21304 43168 21332
rect 27764 21292 27770 21304
rect 43162 21292 43168 21304
rect 43220 21292 43226 21344
rect 43717 21335 43775 21341
rect 43717 21301 43729 21335
rect 43763 21332 43775 21335
rect 44266 21332 44272 21344
rect 43763 21304 44272 21332
rect 43763 21301 43775 21304
rect 43717 21295 43775 21301
rect 44266 21292 44272 21304
rect 44324 21292 44330 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 12342 21088 12348 21140
rect 12400 21128 12406 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 12400 21100 14105 21128
rect 12400 21088 12406 21100
rect 14093 21097 14105 21100
rect 14139 21097 14151 21131
rect 14093 21091 14151 21097
rect 14458 21088 14464 21140
rect 14516 21128 14522 21140
rect 15657 21131 15715 21137
rect 15657 21128 15669 21131
rect 14516 21100 15669 21128
rect 14516 21088 14522 21100
rect 15657 21097 15669 21100
rect 15703 21097 15715 21131
rect 15657 21091 15715 21097
rect 20162 21088 20168 21140
rect 20220 21128 20226 21140
rect 20220 21100 21772 21128
rect 20220 21088 20226 21100
rect 16574 21020 16580 21072
rect 16632 21060 16638 21072
rect 17310 21060 17316 21072
rect 16632 21032 17316 21060
rect 16632 21020 16638 21032
rect 17310 21020 17316 21032
rect 17368 21020 17374 21072
rect 18322 21020 18328 21072
rect 18380 21060 18386 21072
rect 21744 21060 21772 21100
rect 23106 21088 23112 21140
rect 23164 21128 23170 21140
rect 27154 21128 27160 21140
rect 23164 21100 26740 21128
rect 27115 21100 27160 21128
rect 23164 21088 23170 21100
rect 23753 21063 23811 21069
rect 23753 21060 23765 21063
rect 18380 21032 21128 21060
rect 18380 21020 18386 21032
rect 3418 20952 3424 21004
rect 3476 20992 3482 21004
rect 3476 20964 20668 20992
rect 3476 20952 3482 20964
rect 11514 20924 11520 20936
rect 11475 20896 11520 20924
rect 11514 20884 11520 20896
rect 11572 20884 11578 20936
rect 12894 20884 12900 20936
rect 12952 20884 12958 20936
rect 14366 20924 14372 20936
rect 14327 20896 14372 20924
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14826 20924 14832 20936
rect 14787 20896 14832 20924
rect 14826 20884 14832 20896
rect 14884 20884 14890 20936
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 15930 20924 15936 20936
rect 15611 20896 15936 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 15930 20884 15936 20896
rect 15988 20924 15994 20936
rect 16298 20924 16304 20936
rect 15988 20896 16304 20924
rect 15988 20884 15994 20896
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20924 16635 20927
rect 17126 20924 17132 20936
rect 16623 20896 17132 20924
rect 16623 20893 16635 20896
rect 16577 20887 16635 20893
rect 17126 20884 17132 20896
rect 17184 20924 17190 20936
rect 17184 20896 17264 20924
rect 17184 20884 17190 20896
rect 11793 20859 11851 20865
rect 11793 20825 11805 20859
rect 11839 20856 11851 20859
rect 11882 20856 11888 20868
rect 11839 20828 11888 20856
rect 11839 20825 11851 20828
rect 11793 20819 11851 20825
rect 11882 20816 11888 20828
rect 11940 20816 11946 20868
rect 14093 20859 14151 20865
rect 14093 20856 14105 20859
rect 13280 20828 14105 20856
rect 11698 20748 11704 20800
rect 11756 20788 11762 20800
rect 13280 20797 13308 20828
rect 14093 20825 14105 20828
rect 14139 20856 14151 20859
rect 17034 20856 17040 20868
rect 14139 20828 17040 20856
rect 14139 20825 14151 20828
rect 14093 20819 14151 20825
rect 17034 20816 17040 20828
rect 17092 20816 17098 20868
rect 17236 20856 17264 20896
rect 17310 20884 17316 20936
rect 17368 20924 17374 20936
rect 18049 20927 18107 20933
rect 17368 20896 17413 20924
rect 17368 20884 17374 20896
rect 18049 20893 18061 20927
rect 18095 20924 18107 20927
rect 18230 20924 18236 20936
rect 18095 20896 18236 20924
rect 18095 20893 18107 20896
rect 18049 20887 18107 20893
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 19242 20924 19248 20936
rect 19203 20896 19248 20924
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 17586 20856 17592 20868
rect 17236 20828 17592 20856
rect 17586 20816 17592 20828
rect 17644 20816 17650 20868
rect 18598 20816 18604 20868
rect 18656 20856 18662 20868
rect 19429 20859 19487 20865
rect 19429 20856 19441 20859
rect 18656 20828 19441 20856
rect 18656 20816 18662 20828
rect 19429 20825 19441 20828
rect 19475 20825 19487 20859
rect 20640 20856 20668 20964
rect 21100 20933 21128 21032
rect 21744 21032 23765 21060
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20893 21143 20927
rect 21634 20924 21640 20936
rect 21595 20896 21640 20924
rect 21085 20887 21143 20893
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 21744 20933 21772 21032
rect 23753 21029 23765 21032
rect 23799 21029 23811 21063
rect 23753 21023 23811 21029
rect 23842 21020 23848 21072
rect 23900 21060 23906 21072
rect 24949 21063 25007 21069
rect 24949 21060 24961 21063
rect 23900 21032 24961 21060
rect 23900 21020 23906 21032
rect 24949 21029 24961 21032
rect 24995 21029 25007 21063
rect 24949 21023 25007 21029
rect 24394 20992 24400 21004
rect 23216 20964 24400 20992
rect 21729 20927 21787 20933
rect 21729 20893 21741 20927
rect 21775 20893 21787 20927
rect 21729 20887 21787 20893
rect 23106 20856 23112 20868
rect 20640 20828 23112 20856
rect 19429 20819 19487 20825
rect 23106 20816 23112 20828
rect 23164 20816 23170 20868
rect 23216 20865 23244 20964
rect 24394 20952 24400 20964
rect 24452 20952 24458 21004
rect 24578 20952 24584 21004
rect 24636 20992 24642 21004
rect 25682 20992 25688 21004
rect 24636 20964 25268 20992
rect 25643 20964 25688 20992
rect 24636 20952 24642 20964
rect 24670 20924 24676 20936
rect 24631 20896 24676 20924
rect 24670 20884 24676 20896
rect 24728 20884 24734 20936
rect 24946 20884 24952 20936
rect 25004 20884 25010 20936
rect 23201 20859 23259 20865
rect 23201 20825 23213 20859
rect 23247 20825 23259 20859
rect 23566 20856 23572 20868
rect 23527 20828 23572 20856
rect 23201 20819 23259 20825
rect 13265 20791 13323 20797
rect 13265 20788 13277 20791
rect 11756 20760 13277 20788
rect 11756 20748 11762 20760
rect 13265 20757 13277 20760
rect 13311 20757 13323 20791
rect 13265 20751 13323 20757
rect 14277 20791 14335 20797
rect 14277 20757 14289 20791
rect 14323 20788 14335 20791
rect 14458 20788 14464 20800
rect 14323 20760 14464 20788
rect 14323 20757 14335 20760
rect 14277 20751 14335 20757
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 15013 20791 15071 20797
rect 15013 20757 15025 20791
rect 15059 20788 15071 20791
rect 16574 20788 16580 20800
rect 15059 20760 16580 20788
rect 15059 20757 15071 20760
rect 15013 20751 15071 20757
rect 16574 20748 16580 20760
rect 16632 20748 16638 20800
rect 16758 20788 16764 20800
rect 16719 20760 16764 20788
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 16942 20748 16948 20800
rect 17000 20788 17006 20800
rect 17497 20791 17555 20797
rect 17497 20788 17509 20791
rect 17000 20760 17509 20788
rect 17000 20748 17006 20760
rect 17497 20757 17509 20760
rect 17543 20757 17555 20791
rect 18138 20788 18144 20800
rect 18099 20760 18144 20788
rect 17497 20751 17555 20757
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 21913 20791 21971 20797
rect 21913 20788 21925 20791
rect 20772 20760 21925 20788
rect 20772 20748 20778 20760
rect 21913 20757 21925 20760
rect 21959 20757 21971 20791
rect 21913 20751 21971 20757
rect 22830 20748 22836 20800
rect 22888 20788 22894 20800
rect 23216 20788 23244 20819
rect 23566 20816 23572 20828
rect 23624 20816 23630 20868
rect 24581 20859 24639 20865
rect 24581 20825 24593 20859
rect 24627 20856 24639 20859
rect 24964 20856 24992 20884
rect 24627 20828 24992 20856
rect 25240 20856 25268 20964
rect 25682 20952 25688 20964
rect 25740 20952 25746 21004
rect 26712 20992 26740 21100
rect 27154 21088 27160 21100
rect 27212 21088 27218 21140
rect 28626 21128 28632 21140
rect 28587 21100 28632 21128
rect 28626 21088 28632 21100
rect 28684 21088 28690 21140
rect 41386 21100 43208 21128
rect 41386 21060 41414 21100
rect 31726 21032 41414 21060
rect 30009 20995 30067 21001
rect 30009 20992 30021 20995
rect 26712 20964 30021 20992
rect 30009 20961 30021 20964
rect 30055 20961 30067 20995
rect 30009 20955 30067 20961
rect 25406 20924 25412 20936
rect 25367 20896 25412 20924
rect 25406 20884 25412 20896
rect 25464 20884 25470 20936
rect 27985 20927 28043 20933
rect 27985 20893 27997 20927
rect 28031 20924 28043 20927
rect 28534 20924 28540 20936
rect 28031 20896 28540 20924
rect 28031 20893 28043 20896
rect 27985 20887 28043 20893
rect 28534 20884 28540 20896
rect 28592 20884 28598 20936
rect 29546 20924 29552 20936
rect 29507 20896 29552 20924
rect 29546 20884 29552 20896
rect 29604 20884 29610 20936
rect 25240 20828 26096 20856
rect 24627 20825 24639 20828
rect 24581 20819 24639 20825
rect 23382 20788 23388 20800
rect 22888 20760 23244 20788
rect 23343 20760 23388 20788
rect 22888 20748 22894 20760
rect 23382 20748 23388 20760
rect 23440 20748 23446 20800
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 23532 20760 23577 20788
rect 23532 20748 23538 20760
rect 24762 20748 24768 20800
rect 24820 20788 24826 20800
rect 24820 20760 24865 20788
rect 24820 20748 24826 20760
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25682 20788 25688 20800
rect 25372 20760 25688 20788
rect 25372 20748 25378 20760
rect 25682 20748 25688 20760
rect 25740 20748 25746 20800
rect 26068 20788 26096 20828
rect 26694 20816 26700 20868
rect 26752 20816 26758 20868
rect 29730 20856 29736 20868
rect 27540 20828 29592 20856
rect 29691 20828 29736 20856
rect 27540 20788 27568 20828
rect 26068 20760 27568 20788
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 27985 20791 28043 20797
rect 27985 20788 27997 20791
rect 27672 20760 27997 20788
rect 27672 20748 27678 20760
rect 27985 20757 27997 20760
rect 28031 20757 28043 20791
rect 29564 20788 29592 20828
rect 29730 20816 29736 20828
rect 29788 20816 29794 20868
rect 31726 20788 31754 21032
rect 43070 21020 43076 21072
rect 43128 21020 43134 21072
rect 43180 21060 43208 21100
rect 45094 21088 45100 21140
rect 45152 21128 45158 21140
rect 45373 21131 45431 21137
rect 45373 21128 45385 21131
rect 45152 21100 45385 21128
rect 45152 21088 45158 21100
rect 45373 21097 45385 21100
rect 45419 21097 45431 21131
rect 45373 21091 45431 21097
rect 47210 21060 47216 21072
rect 43180 21032 47216 21060
rect 47210 21020 47216 21032
rect 47268 21020 47274 21072
rect 36170 20952 36176 21004
rect 36228 20992 36234 21004
rect 36541 20995 36599 21001
rect 36541 20992 36553 20995
rect 36228 20964 36553 20992
rect 36228 20952 36234 20964
rect 36541 20961 36553 20964
rect 36587 20992 36599 20995
rect 43088 20992 43116 21020
rect 48130 20992 48136 21004
rect 36587 20964 41414 20992
rect 36587 20961 36599 20964
rect 36541 20955 36599 20961
rect 35526 20856 35532 20868
rect 35487 20828 35532 20856
rect 35526 20816 35532 20828
rect 35584 20816 35590 20868
rect 35621 20859 35679 20865
rect 35621 20825 35633 20859
rect 35667 20856 35679 20859
rect 35894 20856 35900 20868
rect 35667 20828 35900 20856
rect 35667 20825 35679 20828
rect 35621 20819 35679 20825
rect 35894 20816 35900 20828
rect 35952 20856 35958 20868
rect 36354 20856 36360 20868
rect 35952 20828 36360 20856
rect 35952 20816 35958 20828
rect 36354 20816 36360 20828
rect 36412 20816 36418 20868
rect 41386 20856 41414 20964
rect 42352 20964 43116 20992
rect 48091 20964 48136 20992
rect 42352 20933 42380 20964
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 42337 20927 42395 20933
rect 42337 20893 42349 20927
rect 42383 20893 42395 20927
rect 42337 20887 42395 20893
rect 42521 20927 42579 20933
rect 42521 20893 42533 20927
rect 42567 20924 42579 20927
rect 42886 20924 42892 20936
rect 42567 20896 42892 20924
rect 42567 20893 42579 20896
rect 42521 20887 42579 20893
rect 42886 20884 42892 20896
rect 42944 20884 42950 20936
rect 43070 20924 43076 20936
rect 43031 20896 43076 20924
rect 43070 20884 43076 20896
rect 43128 20884 43134 20936
rect 43438 20924 43444 20936
rect 43399 20896 43444 20924
rect 43438 20884 43444 20896
rect 43496 20884 43502 20936
rect 44726 20884 44732 20936
rect 44784 20924 44790 20936
rect 45189 20927 45247 20933
rect 45189 20924 45201 20927
rect 44784 20896 45201 20924
rect 44784 20884 44790 20896
rect 45189 20893 45201 20896
rect 45235 20893 45247 20927
rect 46290 20924 46296 20936
rect 46251 20896 46296 20924
rect 45189 20887 45247 20893
rect 46290 20884 46296 20896
rect 46348 20884 46354 20936
rect 44358 20856 44364 20868
rect 41386 20828 44364 20856
rect 44358 20816 44364 20828
rect 44416 20856 44422 20868
rect 45005 20859 45063 20865
rect 45005 20856 45017 20859
rect 44416 20828 45017 20856
rect 44416 20816 44422 20828
rect 45005 20825 45017 20828
rect 45051 20825 45063 20859
rect 45005 20819 45063 20825
rect 46477 20859 46535 20865
rect 46477 20825 46489 20859
rect 46523 20856 46535 20859
rect 47670 20856 47676 20868
rect 46523 20828 47676 20856
rect 46523 20825 46535 20828
rect 46477 20819 46535 20825
rect 47670 20816 47676 20828
rect 47728 20816 47734 20868
rect 29564 20760 31754 20788
rect 42521 20791 42579 20797
rect 27985 20751 28043 20757
rect 42521 20757 42533 20791
rect 42567 20788 42579 20791
rect 42610 20788 42616 20800
rect 42567 20760 42616 20788
rect 42567 20757 42579 20760
rect 42521 20751 42579 20757
rect 42610 20748 42616 20760
rect 42668 20748 42674 20800
rect 44082 20788 44088 20800
rect 44043 20760 44088 20788
rect 44082 20748 44088 20760
rect 44140 20748 44146 20800
rect 47210 20748 47216 20800
rect 47268 20788 47274 20800
rect 47762 20788 47768 20800
rect 47268 20760 47768 20788
rect 47268 20748 47274 20760
rect 47762 20748 47768 20760
rect 47820 20748 47826 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3050 20544 3056 20596
rect 3108 20584 3114 20596
rect 3108 20556 22094 20584
rect 3108 20544 3114 20556
rect 13630 20476 13636 20528
rect 13688 20476 13694 20528
rect 14921 20519 14979 20525
rect 14921 20516 14933 20519
rect 14384 20488 14933 20516
rect 11974 20448 11980 20460
rect 11935 20420 11980 20448
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 12161 20383 12219 20389
rect 12161 20349 12173 20383
rect 12207 20380 12219 20383
rect 12621 20383 12679 20389
rect 12621 20380 12633 20383
rect 12207 20352 12633 20380
rect 12207 20349 12219 20352
rect 12161 20343 12219 20349
rect 12621 20349 12633 20352
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 12897 20383 12955 20389
rect 12897 20349 12909 20383
rect 12943 20380 12955 20383
rect 14090 20380 14096 20392
rect 12943 20352 14096 20380
rect 12943 20349 12955 20352
rect 12897 20343 12955 20349
rect 14090 20340 14096 20352
rect 14148 20340 14154 20392
rect 14274 20340 14280 20392
rect 14332 20380 14338 20392
rect 14384 20389 14412 20488
rect 14921 20485 14933 20488
rect 14967 20485 14979 20519
rect 15121 20519 15179 20525
rect 15121 20516 15133 20519
rect 14921 20479 14979 20485
rect 15028 20488 15133 20516
rect 15028 20448 15056 20488
rect 15121 20485 15133 20488
rect 15167 20485 15179 20519
rect 15121 20479 15179 20485
rect 17034 20476 17040 20528
rect 17092 20516 17098 20528
rect 18969 20519 19027 20525
rect 18969 20516 18981 20519
rect 17092 20488 18981 20516
rect 17092 20476 17098 20488
rect 18969 20485 18981 20488
rect 19015 20485 19027 20519
rect 18969 20479 19027 20485
rect 19185 20519 19243 20525
rect 19185 20485 19197 20519
rect 19231 20516 19243 20519
rect 19794 20516 19800 20528
rect 19231 20488 19800 20516
rect 19231 20485 19243 20488
rect 19185 20479 19243 20485
rect 19794 20476 19800 20488
rect 19852 20476 19858 20528
rect 19886 20476 19892 20528
rect 19944 20516 19950 20528
rect 19981 20519 20039 20525
rect 19981 20516 19993 20519
rect 19944 20488 19993 20516
rect 19944 20476 19950 20488
rect 19981 20485 19993 20488
rect 20027 20485 20039 20519
rect 19981 20479 20039 20485
rect 20162 20476 20168 20528
rect 20220 20525 20226 20528
rect 20220 20519 20239 20525
rect 20227 20485 20239 20519
rect 20220 20479 20239 20485
rect 20220 20476 20226 20479
rect 16761 20451 16819 20457
rect 16761 20448 16773 20451
rect 14936 20420 15056 20448
rect 16684 20420 16773 20448
rect 14936 20392 14964 20420
rect 14369 20383 14427 20389
rect 14369 20380 14381 20383
rect 14332 20352 14381 20380
rect 14332 20340 14338 20352
rect 14369 20349 14381 20352
rect 14415 20349 14427 20383
rect 14369 20343 14427 20349
rect 14918 20340 14924 20392
rect 14976 20340 14982 20392
rect 16298 20340 16304 20392
rect 16356 20380 16362 20392
rect 16684 20380 16712 20420
rect 16761 20417 16773 20420
rect 16807 20417 16819 20451
rect 16761 20411 16819 20417
rect 16850 20408 16856 20460
rect 16908 20448 16914 20460
rect 17589 20451 17647 20457
rect 17589 20448 17601 20451
rect 16908 20420 17601 20448
rect 16908 20408 16914 20420
rect 17589 20417 17601 20420
rect 17635 20417 17647 20451
rect 17862 20448 17868 20460
rect 17823 20420 17868 20448
rect 17589 20411 17647 20417
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 18046 20448 18052 20460
rect 18007 20420 18052 20448
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 21818 20448 21824 20460
rect 21779 20420 21824 20448
rect 21818 20408 21824 20420
rect 21876 20408 21882 20460
rect 22066 20448 22094 20556
rect 23474 20544 23480 20596
rect 23532 20584 23538 20596
rect 24305 20587 24363 20593
rect 24305 20584 24317 20587
rect 23532 20556 24317 20584
rect 23532 20544 23538 20556
rect 24305 20553 24317 20556
rect 24351 20584 24363 20587
rect 24762 20584 24768 20596
rect 24351 20556 24768 20584
rect 24351 20553 24363 20556
rect 24305 20547 24363 20553
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 25406 20544 25412 20596
rect 25464 20584 25470 20596
rect 25501 20587 25559 20593
rect 25501 20584 25513 20587
rect 25464 20556 25513 20584
rect 25464 20544 25470 20556
rect 25501 20553 25513 20556
rect 25547 20553 25559 20587
rect 25501 20547 25559 20553
rect 26234 20544 26240 20596
rect 26292 20584 26298 20596
rect 27157 20587 27215 20593
rect 27157 20584 27169 20587
rect 26292 20556 27169 20584
rect 26292 20544 26298 20556
rect 27157 20553 27169 20556
rect 27203 20553 27215 20587
rect 27157 20547 27215 20553
rect 29181 20587 29239 20593
rect 29181 20553 29193 20587
rect 29227 20584 29239 20587
rect 29730 20584 29736 20596
rect 29227 20556 29736 20584
rect 29227 20553 29239 20556
rect 29181 20547 29239 20553
rect 29730 20544 29736 20556
rect 29788 20544 29794 20596
rect 42613 20587 42671 20593
rect 42613 20553 42625 20587
rect 42659 20584 42671 20587
rect 43070 20584 43076 20596
rect 42659 20556 43076 20584
rect 42659 20553 42671 20556
rect 42613 20547 42671 20553
rect 43070 20544 43076 20556
rect 43128 20544 43134 20596
rect 43346 20584 43352 20596
rect 43307 20556 43352 20584
rect 43346 20544 43352 20556
rect 43404 20544 43410 20596
rect 43441 20587 43499 20593
rect 43441 20553 43453 20587
rect 43487 20553 43499 20587
rect 48041 20587 48099 20593
rect 48041 20584 48053 20587
rect 43441 20547 43499 20553
rect 44192 20556 48053 20584
rect 23566 20476 23572 20528
rect 23624 20516 23630 20528
rect 23937 20519 23995 20525
rect 23937 20516 23949 20519
rect 23624 20488 23949 20516
rect 23624 20476 23630 20488
rect 23937 20485 23949 20488
rect 23983 20485 23995 20519
rect 23937 20479 23995 20485
rect 24153 20519 24211 20525
rect 24153 20485 24165 20519
rect 24199 20516 24211 20519
rect 24854 20516 24860 20528
rect 24199 20488 24860 20516
rect 24199 20485 24211 20488
rect 24153 20479 24211 20485
rect 24854 20476 24860 20488
rect 24912 20476 24918 20528
rect 28994 20516 29000 20528
rect 24964 20488 29000 20516
rect 24964 20448 24992 20488
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 43456 20516 43484 20547
rect 42628 20488 43484 20516
rect 42628 20460 42656 20488
rect 22066 20420 24992 20448
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20448 25559 20451
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 25547 20420 26065 20448
rect 25547 20417 25559 20420
rect 25501 20411 25559 20417
rect 26053 20417 26065 20420
rect 26099 20448 26111 20451
rect 26234 20448 26240 20460
rect 26099 20420 26240 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 26970 20448 26976 20460
rect 26931 20420 26976 20448
rect 26970 20408 26976 20420
rect 27028 20408 27034 20460
rect 29089 20451 29147 20457
rect 29089 20417 29101 20451
rect 29135 20448 29147 20451
rect 29730 20448 29736 20460
rect 29135 20420 29736 20448
rect 29135 20417 29147 20420
rect 29089 20411 29147 20417
rect 29730 20408 29736 20420
rect 29788 20448 29794 20460
rect 30374 20448 30380 20460
rect 29788 20420 30380 20448
rect 29788 20408 29794 20420
rect 30374 20408 30380 20420
rect 30432 20408 30438 20460
rect 30469 20451 30527 20457
rect 30469 20417 30481 20451
rect 30515 20448 30527 20451
rect 30834 20448 30840 20460
rect 30515 20420 30840 20448
rect 30515 20417 30527 20420
rect 30469 20411 30527 20417
rect 30834 20408 30840 20420
rect 30892 20408 30898 20460
rect 33410 20448 33416 20460
rect 33371 20420 33416 20448
rect 33410 20408 33416 20420
rect 33468 20408 33474 20460
rect 42429 20451 42487 20457
rect 42429 20417 42441 20451
rect 42475 20417 42487 20451
rect 42610 20448 42616 20460
rect 42571 20420 42616 20448
rect 42429 20411 42487 20417
rect 42444 20380 42472 20411
rect 42610 20408 42616 20420
rect 42668 20408 42674 20460
rect 42794 20408 42800 20460
rect 42852 20448 42858 20460
rect 43073 20451 43131 20457
rect 43073 20448 43085 20451
rect 42852 20420 43085 20448
rect 42852 20408 42858 20420
rect 43073 20417 43085 20420
rect 43119 20417 43131 20451
rect 43254 20448 43260 20460
rect 43215 20420 43260 20448
rect 43073 20411 43131 20417
rect 43254 20408 43260 20420
rect 43312 20408 43318 20460
rect 43622 20448 43628 20460
rect 43583 20420 43628 20448
rect 43622 20408 43628 20420
rect 43680 20408 43686 20460
rect 43162 20380 43168 20392
rect 16356 20352 20576 20380
rect 42444 20352 43168 20380
rect 16356 20340 16362 20352
rect 14458 20272 14464 20324
rect 14516 20312 14522 20324
rect 15289 20315 15347 20321
rect 15289 20312 15301 20315
rect 14516 20284 15301 20312
rect 14516 20272 14522 20284
rect 15289 20281 15301 20284
rect 15335 20312 15347 20315
rect 19337 20315 19395 20321
rect 15335 20284 19196 20312
rect 15335 20281 15347 20284
rect 15289 20275 15347 20281
rect 15102 20244 15108 20256
rect 15063 20216 15108 20244
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 16850 20244 16856 20256
rect 16811 20216 16856 20244
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 19168 20253 19196 20284
rect 19337 20281 19349 20315
rect 19383 20312 19395 20315
rect 20438 20312 20444 20324
rect 19383 20284 20444 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 20438 20272 20444 20284
rect 20496 20272 20502 20324
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 17276 20216 17417 20244
rect 17276 20204 17282 20216
rect 17405 20213 17417 20216
rect 17451 20213 17463 20247
rect 17405 20207 17463 20213
rect 19153 20247 19211 20253
rect 19153 20213 19165 20247
rect 19199 20213 19211 20247
rect 19153 20207 19211 20213
rect 19794 20204 19800 20256
rect 19852 20244 19858 20256
rect 20165 20247 20223 20253
rect 20165 20244 20177 20247
rect 19852 20216 20177 20244
rect 19852 20204 19858 20216
rect 20165 20213 20177 20216
rect 20211 20213 20223 20247
rect 20165 20207 20223 20213
rect 20349 20247 20407 20253
rect 20349 20213 20361 20247
rect 20395 20244 20407 20247
rect 20548 20244 20576 20352
rect 43162 20340 43168 20352
rect 43220 20340 43226 20392
rect 43806 20340 43812 20392
rect 43864 20380 43870 20392
rect 44085 20383 44143 20389
rect 44085 20380 44097 20383
rect 43864 20352 44097 20380
rect 43864 20340 43870 20352
rect 44085 20349 44097 20352
rect 44131 20349 44143 20383
rect 44085 20343 44143 20349
rect 28810 20272 28816 20324
rect 28868 20312 28874 20324
rect 44192 20312 44220 20556
rect 48041 20553 48053 20556
rect 48087 20553 48099 20587
rect 48041 20547 48099 20553
rect 44266 20476 44272 20528
rect 44324 20516 44330 20528
rect 45373 20519 45431 20525
rect 45373 20516 45385 20519
rect 44324 20488 45385 20516
rect 44324 20476 44330 20488
rect 45373 20485 45385 20488
rect 45419 20485 45431 20519
rect 47946 20516 47952 20528
rect 47907 20488 47952 20516
rect 45373 20479 45431 20485
rect 47946 20476 47952 20488
rect 48004 20476 48010 20528
rect 44358 20448 44364 20460
rect 44319 20420 44364 20448
rect 44358 20408 44364 20420
rect 44416 20408 44422 20460
rect 44545 20451 44603 20457
rect 44545 20417 44557 20451
rect 44591 20448 44603 20451
rect 44726 20448 44732 20460
rect 44591 20420 44732 20448
rect 44591 20417 44603 20420
rect 44545 20411 44603 20417
rect 44726 20408 44732 20420
rect 44784 20408 44790 20460
rect 44450 20340 44456 20392
rect 44508 20380 44514 20392
rect 45189 20383 45247 20389
rect 45189 20380 45201 20383
rect 44508 20352 45201 20380
rect 44508 20340 44514 20352
rect 45189 20349 45201 20352
rect 45235 20349 45247 20383
rect 45738 20380 45744 20392
rect 45699 20352 45744 20380
rect 45189 20343 45247 20349
rect 45738 20340 45744 20352
rect 45796 20340 45802 20392
rect 28868 20284 44220 20312
rect 28868 20272 28874 20284
rect 20395 20216 20576 20244
rect 20395 20213 20407 20216
rect 20349 20207 20407 20213
rect 21726 20204 21732 20256
rect 21784 20244 21790 20256
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 21784 20216 22017 20244
rect 21784 20204 21790 20216
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 24118 20244 24124 20256
rect 24079 20216 24124 20244
rect 22005 20207 22063 20213
rect 24118 20204 24124 20216
rect 24176 20204 24182 20256
rect 25314 20204 25320 20256
rect 25372 20244 25378 20256
rect 26145 20247 26203 20253
rect 26145 20244 26157 20247
rect 25372 20216 26157 20244
rect 25372 20204 25378 20216
rect 26145 20213 26157 20216
rect 26191 20213 26203 20247
rect 26145 20207 26203 20213
rect 30561 20247 30619 20253
rect 30561 20213 30573 20247
rect 30607 20244 30619 20247
rect 30650 20244 30656 20256
rect 30607 20216 30656 20244
rect 30607 20213 30619 20216
rect 30561 20207 30619 20213
rect 30650 20204 30656 20216
rect 30708 20204 30714 20256
rect 33226 20244 33232 20256
rect 33187 20216 33232 20244
rect 33226 20204 33232 20216
rect 33284 20204 33290 20256
rect 43254 20204 43260 20256
rect 43312 20244 43318 20256
rect 44361 20247 44419 20253
rect 44361 20244 44373 20247
rect 43312 20216 44373 20244
rect 43312 20204 43318 20216
rect 44361 20213 44373 20216
rect 44407 20213 44419 20247
rect 44361 20207 44419 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 12894 20040 12900 20052
rect 12855 20012 12900 20040
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 14090 20040 14096 20052
rect 14051 20012 14096 20040
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14645 20043 14703 20049
rect 14645 20040 14657 20043
rect 14332 20012 14657 20040
rect 14332 20000 14338 20012
rect 14645 20009 14657 20012
rect 14691 20009 14703 20043
rect 14645 20003 14703 20009
rect 14918 20000 14924 20052
rect 14976 20040 14982 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 14976 20012 16313 20040
rect 14976 20000 14982 20012
rect 16301 20009 16313 20012
rect 16347 20009 16359 20043
rect 16301 20003 16359 20009
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 19794 20040 19800 20052
rect 17920 20012 19380 20040
rect 19755 20012 19800 20040
rect 17920 20000 17926 20012
rect 15194 19932 15200 19984
rect 15252 19972 15258 19984
rect 15473 19975 15531 19981
rect 15473 19972 15485 19975
rect 15252 19944 15485 19972
rect 15252 19932 15258 19944
rect 15473 19941 15485 19944
rect 15519 19941 15531 19975
rect 15473 19935 15531 19941
rect 16485 19975 16543 19981
rect 16485 19941 16497 19975
rect 16531 19941 16543 19975
rect 19352 19972 19380 20012
rect 19794 20000 19800 20012
rect 19852 20000 19858 20052
rect 20162 20000 20168 20052
rect 20220 20040 20226 20052
rect 43073 20043 43131 20049
rect 20220 20012 22094 20040
rect 20220 20000 20226 20012
rect 20809 19975 20867 19981
rect 20809 19972 20821 19975
rect 19352 19944 20821 19972
rect 16485 19935 16543 19941
rect 20809 19941 20821 19944
rect 20855 19941 20867 19975
rect 20809 19935 20867 19941
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19836 12863 19839
rect 12986 19836 12992 19848
rect 12851 19808 12992 19836
rect 12851 19805 12863 19808
rect 12805 19799 12863 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 14274 19839 14332 19845
rect 14274 19805 14286 19839
rect 14320 19836 14332 19839
rect 14458 19836 14464 19848
rect 14320 19808 14464 19836
rect 14320 19805 14332 19808
rect 14274 19799 14332 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19836 14795 19839
rect 15197 19839 15255 19845
rect 15197 19836 15209 19839
rect 14783 19808 15209 19836
rect 14783 19805 14795 19808
rect 14737 19799 14795 19805
rect 15197 19805 15209 19808
rect 15243 19836 15255 19839
rect 16500 19836 16528 19935
rect 16942 19904 16948 19916
rect 16903 19876 16948 19904
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17218 19904 17224 19916
rect 17179 19876 17224 19904
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 17586 19864 17592 19916
rect 17644 19904 17650 19916
rect 21818 19904 21824 19916
rect 17644 19876 21824 19904
rect 17644 19864 17650 19876
rect 21818 19864 21824 19876
rect 21876 19864 21882 19916
rect 19426 19836 19432 19848
rect 15243 19808 16528 19836
rect 19339 19808 19432 19836
rect 15243 19805 15255 19808
rect 15197 19799 15255 19805
rect 19426 19796 19432 19808
rect 19484 19836 19490 19848
rect 19978 19836 19984 19848
rect 19484 19808 19984 19836
rect 19484 19796 19490 19808
rect 19978 19796 19984 19808
rect 20036 19836 20042 19848
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 20036 19808 20269 19836
rect 20036 19796 20042 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 20714 19836 20720 19848
rect 20671 19808 20720 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 21726 19836 21732 19848
rect 21687 19808 21732 19836
rect 21726 19796 21732 19808
rect 21784 19796 21790 19848
rect 15102 19728 15108 19780
rect 15160 19768 15166 19780
rect 16117 19771 16175 19777
rect 16117 19768 16129 19771
rect 15160 19740 16129 19768
rect 15160 19728 15166 19740
rect 16117 19737 16129 19740
rect 16163 19737 16175 19771
rect 16117 19731 16175 19737
rect 16298 19728 16304 19780
rect 16356 19777 16362 19780
rect 16356 19771 16375 19777
rect 16363 19737 16375 19771
rect 19150 19768 19156 19780
rect 18446 19740 19156 19768
rect 16356 19731 16375 19737
rect 16356 19728 16362 19731
rect 19150 19728 19156 19740
rect 19208 19728 19214 19780
rect 19245 19771 19303 19777
rect 19245 19737 19257 19771
rect 19291 19737 19303 19771
rect 19245 19731 19303 19737
rect 19521 19771 19579 19777
rect 19521 19737 19533 19771
rect 19567 19768 19579 19771
rect 20346 19768 20352 19780
rect 19567 19740 20352 19768
rect 19567 19737 19579 19740
rect 19521 19731 19579 19737
rect 14274 19700 14280 19712
rect 14235 19672 14280 19700
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 15528 19672 15669 19700
rect 15528 19660 15534 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 15657 19663 15715 19669
rect 18046 19660 18052 19712
rect 18104 19700 18110 19712
rect 18693 19703 18751 19709
rect 18693 19700 18705 19703
rect 18104 19672 18705 19700
rect 18104 19660 18110 19672
rect 18693 19669 18705 19672
rect 18739 19700 18751 19703
rect 19260 19700 19288 19731
rect 20346 19728 20352 19740
rect 20404 19768 20410 19780
rect 20441 19771 20499 19777
rect 20441 19768 20453 19771
rect 20404 19740 20453 19768
rect 20404 19728 20410 19740
rect 20441 19737 20453 19740
rect 20487 19737 20499 19771
rect 21744 19768 21772 19796
rect 20441 19731 20499 19737
rect 20640 19740 21772 19768
rect 22066 19768 22094 20012
rect 43073 20009 43085 20043
rect 43119 20040 43131 20043
rect 43622 20040 43628 20052
rect 43119 20012 43628 20040
rect 43119 20009 43131 20012
rect 43073 20003 43131 20009
rect 43622 20000 43628 20012
rect 43680 20000 43686 20052
rect 43806 20000 43812 20052
rect 43864 20040 43870 20052
rect 44174 20040 44180 20052
rect 43864 20012 44180 20040
rect 43864 20000 43870 20012
rect 44174 20000 44180 20012
rect 44232 20040 44238 20052
rect 44634 20040 44640 20052
rect 44232 20012 44640 20040
rect 44232 20000 44238 20012
rect 44634 20000 44640 20012
rect 44692 20000 44698 20052
rect 45833 20043 45891 20049
rect 45833 20009 45845 20043
rect 45879 20040 45891 20043
rect 46290 20040 46296 20052
rect 45879 20012 46296 20040
rect 45879 20009 45891 20012
rect 45833 20003 45891 20009
rect 46290 20000 46296 20012
rect 46348 20000 46354 20052
rect 23474 19932 23480 19984
rect 23532 19972 23538 19984
rect 23569 19975 23627 19981
rect 23569 19972 23581 19975
rect 23532 19944 23581 19972
rect 23532 19932 23538 19944
rect 23569 19941 23581 19944
rect 23615 19941 23627 19975
rect 23569 19935 23627 19941
rect 29178 19932 29184 19984
rect 29236 19972 29242 19984
rect 32214 19972 32220 19984
rect 29236 19944 32220 19972
rect 29236 19932 29242 19944
rect 32214 19932 32220 19944
rect 32272 19932 32278 19984
rect 43346 19932 43352 19984
rect 43404 19972 43410 19984
rect 43901 19975 43959 19981
rect 43901 19972 43913 19975
rect 43404 19944 43913 19972
rect 43404 19932 43410 19944
rect 43901 19941 43913 19944
rect 43947 19941 43959 19975
rect 43901 19935 43959 19941
rect 45002 19932 45008 19984
rect 45060 19972 45066 19984
rect 47394 19972 47400 19984
rect 45060 19944 47400 19972
rect 45060 19932 45066 19944
rect 47394 19932 47400 19944
rect 47452 19932 47458 19984
rect 24949 19907 25007 19913
rect 24949 19873 24961 19907
rect 24995 19904 25007 19907
rect 25130 19904 25136 19916
rect 24995 19876 25136 19904
rect 24995 19873 25007 19876
rect 24949 19867 25007 19873
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19836 23903 19839
rect 24964 19836 24992 19867
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 25406 19904 25412 19916
rect 25367 19876 25412 19904
rect 25406 19864 25412 19876
rect 25464 19864 25470 19916
rect 30466 19904 30472 19916
rect 30427 19876 30472 19904
rect 30466 19864 30472 19876
rect 30524 19864 30530 19916
rect 30650 19904 30656 19916
rect 30611 19876 30656 19904
rect 30650 19864 30656 19876
rect 30708 19864 30714 19916
rect 33137 19907 33195 19913
rect 33137 19873 33149 19907
rect 33183 19904 33195 19907
rect 33183 19876 41414 19904
rect 33183 19873 33195 19876
rect 33137 19867 33195 19873
rect 23891 19808 24992 19836
rect 25041 19839 25099 19845
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 25041 19805 25053 19839
rect 25087 19805 25099 19839
rect 25041 19799 25099 19805
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19836 26019 19839
rect 26970 19836 26976 19848
rect 26007 19808 26976 19836
rect 26007 19805 26019 19808
rect 25961 19799 26019 19805
rect 23566 19768 23572 19780
rect 22066 19740 23572 19768
rect 20640 19712 20668 19740
rect 23566 19728 23572 19740
rect 23624 19728 23630 19780
rect 23753 19771 23811 19777
rect 23753 19737 23765 19771
rect 23799 19768 23811 19771
rect 24118 19768 24124 19780
rect 23799 19740 24124 19768
rect 23799 19737 23811 19740
rect 23753 19731 23811 19737
rect 24118 19728 24124 19740
rect 24176 19768 24182 19780
rect 24762 19768 24768 19780
rect 24176 19740 24768 19768
rect 24176 19728 24182 19740
rect 24762 19728 24768 19740
rect 24820 19768 24826 19780
rect 25056 19768 25084 19799
rect 26970 19796 26976 19808
rect 27028 19796 27034 19848
rect 29638 19796 29644 19848
rect 29696 19836 29702 19848
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 29696 19808 29745 19836
rect 29696 19796 29702 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 32306 19768 32312 19780
rect 24820 19740 25084 19768
rect 32267 19740 32312 19768
rect 24820 19728 24826 19740
rect 32306 19728 32312 19740
rect 32364 19728 32370 19780
rect 33226 19728 33232 19780
rect 33284 19768 33290 19780
rect 34146 19768 34152 19780
rect 33284 19740 33329 19768
rect 34107 19740 34152 19768
rect 33284 19728 33290 19740
rect 34146 19728 34152 19740
rect 34204 19728 34210 19780
rect 41386 19768 41414 19876
rect 42886 19864 42892 19916
rect 42944 19904 42950 19916
rect 44542 19904 44548 19916
rect 42944 19876 43300 19904
rect 42944 19864 42950 19876
rect 43272 19848 43300 19876
rect 43824 19876 44548 19904
rect 42978 19796 42984 19848
rect 43036 19836 43042 19848
rect 43073 19839 43131 19845
rect 43073 19836 43085 19839
rect 43036 19808 43085 19836
rect 43036 19796 43042 19808
rect 43073 19805 43085 19808
rect 43119 19805 43131 19839
rect 43254 19836 43260 19848
rect 43215 19808 43260 19836
rect 43073 19799 43131 19805
rect 43254 19796 43260 19808
rect 43312 19796 43318 19848
rect 43824 19845 43852 19876
rect 44542 19864 44548 19876
rect 44600 19864 44606 19916
rect 45189 19907 45247 19913
rect 45189 19873 45201 19907
rect 45235 19904 45247 19907
rect 46293 19907 46351 19913
rect 46293 19904 46305 19907
rect 45235 19876 46305 19904
rect 45235 19873 45247 19876
rect 45189 19867 45247 19873
rect 46293 19873 46305 19876
rect 46339 19873 46351 19907
rect 46293 19867 46351 19873
rect 43809 19839 43867 19845
rect 43809 19805 43821 19839
rect 43855 19805 43867 19839
rect 43809 19799 43867 19805
rect 43993 19839 44051 19845
rect 43993 19805 44005 19839
rect 44039 19836 44051 19839
rect 44634 19836 44640 19848
rect 44039 19808 44640 19836
rect 44039 19805 44051 19808
rect 43993 19799 44051 19805
rect 44634 19796 44640 19808
rect 44692 19796 44698 19848
rect 45646 19768 45652 19780
rect 41386 19740 45652 19768
rect 45646 19728 45652 19740
rect 45704 19728 45710 19780
rect 46477 19771 46535 19777
rect 46477 19737 46489 19771
rect 46523 19768 46535 19771
rect 47210 19768 47216 19780
rect 46523 19740 47216 19768
rect 46523 19737 46535 19740
rect 46477 19731 46535 19737
rect 47210 19728 47216 19740
rect 47268 19728 47274 19780
rect 48130 19768 48136 19780
rect 48091 19740 48136 19768
rect 48130 19728 48136 19740
rect 48188 19728 48194 19780
rect 18739 19672 19288 19700
rect 19613 19703 19671 19709
rect 18739 19669 18751 19672
rect 18693 19663 18751 19669
rect 19613 19669 19625 19703
rect 19659 19700 19671 19703
rect 20530 19700 20536 19712
rect 19659 19672 20536 19700
rect 19659 19669 19671 19672
rect 19613 19663 19671 19669
rect 20530 19660 20536 19672
rect 20588 19660 20594 19712
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 21818 19700 21824 19712
rect 21779 19672 21824 19700
rect 21818 19660 21824 19672
rect 21876 19660 21882 19712
rect 24670 19660 24676 19712
rect 24728 19700 24734 19712
rect 26053 19703 26111 19709
rect 26053 19700 26065 19703
rect 24728 19672 26065 19700
rect 24728 19660 24734 19672
rect 26053 19669 26065 19672
rect 26099 19669 26111 19703
rect 29546 19700 29552 19712
rect 29459 19672 29552 19700
rect 26053 19663 26111 19669
rect 29546 19660 29552 19672
rect 29604 19700 29610 19712
rect 29914 19700 29920 19712
rect 29604 19672 29920 19700
rect 29604 19660 29610 19672
rect 29914 19660 29920 19672
rect 29972 19660 29978 19712
rect 31110 19660 31116 19712
rect 31168 19700 31174 19712
rect 36538 19700 36544 19712
rect 31168 19672 36544 19700
rect 31168 19660 31174 19672
rect 36538 19660 36544 19672
rect 36596 19660 36602 19712
rect 45922 19660 45928 19712
rect 45980 19700 45986 19712
rect 47394 19700 47400 19712
rect 45980 19672 47400 19700
rect 45980 19660 45986 19672
rect 47394 19660 47400 19672
rect 47452 19660 47458 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 13630 19456 13636 19508
rect 13688 19496 13694 19508
rect 13725 19499 13783 19505
rect 13725 19496 13737 19499
rect 13688 19468 13737 19496
rect 13688 19456 13694 19468
rect 13725 19465 13737 19468
rect 13771 19465 13783 19499
rect 13725 19459 13783 19465
rect 14918 19456 14924 19508
rect 14976 19496 14982 19508
rect 15473 19499 15531 19505
rect 15473 19496 15485 19499
rect 14976 19468 15485 19496
rect 14976 19456 14982 19468
rect 15473 19465 15485 19468
rect 15519 19465 15531 19499
rect 15473 19459 15531 19465
rect 19150 19456 19156 19508
rect 19208 19496 19214 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19208 19468 19625 19496
rect 19208 19456 19214 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 20732 19468 23520 19496
rect 15102 19388 15108 19440
rect 15160 19428 15166 19440
rect 16942 19428 16948 19440
rect 15160 19400 16948 19428
rect 15160 19388 15166 19400
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 12802 19360 12808 19372
rect 12763 19332 12808 19360
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 13633 19363 13691 19369
rect 13633 19360 13645 19363
rect 13044 19332 13645 19360
rect 13044 19320 13050 19332
rect 13633 19329 13645 19332
rect 13679 19360 13691 19363
rect 13722 19360 13728 19372
rect 13679 19332 13728 19360
rect 13679 19329 13691 19332
rect 13633 19323 13691 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 15304 19369 15332 19400
rect 16942 19388 16948 19400
rect 17000 19428 17006 19440
rect 17405 19431 17463 19437
rect 17000 19400 17264 19428
rect 17000 19388 17006 19400
rect 15289 19363 15347 19369
rect 15289 19329 15301 19363
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 15565 19363 15623 19369
rect 15565 19329 15577 19363
rect 15611 19360 15623 19363
rect 16850 19360 16856 19372
rect 15611 19332 16856 19360
rect 15611 19329 15623 19332
rect 15565 19323 15623 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 14274 19292 14280 19304
rect 12943 19264 14280 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19292 15163 19295
rect 15194 19292 15200 19304
rect 15151 19264 15200 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15580 19292 15608 19323
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 17236 19369 17264 19400
rect 17405 19397 17417 19431
rect 17451 19428 17463 19431
rect 18138 19428 18144 19440
rect 17451 19400 18144 19428
rect 17451 19397 17463 19400
rect 17405 19391 17463 19397
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 20622 19428 20628 19440
rect 19536 19400 20628 19428
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 19058 19360 19064 19372
rect 19019 19332 19064 19360
rect 17221 19323 17279 19329
rect 19058 19320 19064 19332
rect 19116 19320 19122 19372
rect 19150 19320 19156 19372
rect 19208 19360 19214 19372
rect 19536 19369 19564 19400
rect 20622 19388 20628 19400
rect 20680 19388 20686 19440
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19208 19332 19533 19360
rect 19208 19320 19214 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 20732 19369 20760 19468
rect 21818 19388 21824 19440
rect 21876 19428 21882 19440
rect 23492 19428 23520 19468
rect 23566 19456 23572 19508
rect 23624 19496 23630 19508
rect 26053 19499 26111 19505
rect 26053 19496 26065 19499
rect 23624 19468 26065 19496
rect 23624 19456 23630 19468
rect 26053 19465 26065 19468
rect 26099 19465 26111 19499
rect 28074 19496 28080 19508
rect 28035 19468 28080 19496
rect 26053 19459 26111 19465
rect 28074 19456 28080 19468
rect 28132 19496 28138 19508
rect 29638 19496 29644 19508
rect 28132 19468 28672 19496
rect 29599 19468 29644 19496
rect 28132 19456 28138 19468
rect 28644 19440 28672 19468
rect 29638 19456 29644 19468
rect 29696 19456 29702 19508
rect 33594 19496 33600 19508
rect 32048 19468 33600 19496
rect 21876 19400 22586 19428
rect 23492 19400 23888 19428
rect 21876 19388 21882 19400
rect 23860 19369 23888 19400
rect 24854 19388 24860 19440
rect 24912 19428 24918 19440
rect 28626 19428 28632 19440
rect 24912 19400 25070 19428
rect 28539 19400 28632 19428
rect 24912 19388 24918 19400
rect 28626 19388 28632 19400
rect 28684 19428 28690 19440
rect 29089 19431 29147 19437
rect 29089 19428 29101 19431
rect 28684 19400 29101 19428
rect 28684 19388 28690 19400
rect 29089 19397 29101 19400
rect 29135 19397 29147 19431
rect 29089 19391 29147 19397
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20588 19332 20729 19360
rect 20588 19320 20594 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19360 23903 19363
rect 24026 19360 24032 19372
rect 23891 19332 24032 19360
rect 23891 19329 23903 19332
rect 23845 19323 23903 19329
rect 24026 19320 24032 19332
rect 24084 19320 24090 19372
rect 26418 19320 26424 19372
rect 26476 19360 26482 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26476 19332 26985 19360
rect 26476 19320 26482 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 28445 19363 28503 19369
rect 28445 19329 28457 19363
rect 28491 19329 28503 19363
rect 29457 19363 29515 19369
rect 29457 19360 29469 19363
rect 28445 19323 28503 19329
rect 29196 19332 29469 19360
rect 20806 19292 20812 19304
rect 15488 19264 15608 19292
rect 20767 19264 20812 19292
rect 14292 19224 14320 19252
rect 15488 19224 15516 19264
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 21818 19292 21824 19304
rect 21779 19264 21824 19292
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 22097 19295 22155 19301
rect 22097 19292 22109 19295
rect 21928 19264 22109 19292
rect 14292 19196 15516 19224
rect 21085 19227 21143 19233
rect 21085 19193 21097 19227
rect 21131 19224 21143 19227
rect 21928 19224 21956 19264
rect 22097 19261 22109 19264
rect 22143 19261 22155 19295
rect 24302 19292 24308 19304
rect 24263 19264 24308 19292
rect 22097 19255 22155 19261
rect 24302 19252 24308 19264
rect 24360 19252 24366 19304
rect 24578 19292 24584 19304
rect 24539 19264 24584 19292
rect 24578 19252 24584 19264
rect 24636 19252 24642 19304
rect 28460 19236 28488 19323
rect 28813 19295 28871 19301
rect 28813 19261 28825 19295
rect 28859 19292 28871 19295
rect 29196 19292 29224 19332
rect 29457 19329 29469 19332
rect 29503 19329 29515 19363
rect 29457 19323 29515 19329
rect 28859 19264 29224 19292
rect 28859 19261 28871 19264
rect 28813 19255 28871 19261
rect 29270 19252 29276 19304
rect 29328 19292 29334 19304
rect 32048 19292 32076 19468
rect 33594 19456 33600 19468
rect 33652 19456 33658 19508
rect 45465 19499 45523 19505
rect 45465 19465 45477 19499
rect 45511 19496 45523 19499
rect 47486 19496 47492 19508
rect 45511 19468 47492 19496
rect 45511 19465 45523 19468
rect 45465 19459 45523 19465
rect 47486 19456 47492 19468
rect 47544 19456 47550 19508
rect 47670 19496 47676 19508
rect 47631 19468 47676 19496
rect 47670 19456 47676 19468
rect 47728 19456 47734 19508
rect 32214 19388 32220 19440
rect 32272 19428 32278 19440
rect 32309 19431 32367 19437
rect 32309 19428 32321 19431
rect 32272 19400 32321 19428
rect 32272 19388 32278 19400
rect 32309 19397 32321 19400
rect 32355 19397 32367 19431
rect 46290 19428 46296 19440
rect 46251 19400 46296 19428
rect 32309 19391 32367 19397
rect 46290 19388 46296 19400
rect 46348 19388 46354 19440
rect 46477 19431 46535 19437
rect 46477 19397 46489 19431
rect 46523 19428 46535 19431
rect 47118 19428 47124 19440
rect 46523 19400 47124 19428
rect 46523 19397 46535 19400
rect 46477 19391 46535 19397
rect 47118 19388 47124 19400
rect 47176 19388 47182 19440
rect 36538 19320 36544 19372
rect 36596 19360 36602 19372
rect 43073 19363 43131 19369
rect 43073 19360 43085 19363
rect 36596 19332 43085 19360
rect 36596 19320 36602 19332
rect 43073 19329 43085 19332
rect 43119 19360 43131 19363
rect 45002 19360 45008 19372
rect 43119 19332 45008 19360
rect 43119 19329 43131 19332
rect 43073 19323 43131 19329
rect 45002 19320 45008 19332
rect 45060 19320 45066 19372
rect 45646 19360 45652 19372
rect 45607 19332 45652 19360
rect 45646 19320 45652 19332
rect 45704 19320 45710 19372
rect 46198 19320 46204 19372
rect 46256 19360 46262 19372
rect 46385 19363 46443 19369
rect 46385 19360 46397 19363
rect 46256 19332 46397 19360
rect 46256 19320 46262 19332
rect 46385 19329 46397 19332
rect 46431 19329 46443 19363
rect 46385 19323 46443 19329
rect 47394 19320 47400 19372
rect 47452 19360 47458 19372
rect 47581 19363 47639 19369
rect 47581 19360 47593 19363
rect 47452 19332 47593 19360
rect 47452 19320 47458 19332
rect 47581 19329 47593 19332
rect 47627 19329 47639 19363
rect 47581 19323 47639 19329
rect 32217 19295 32275 19301
rect 32217 19292 32229 19295
rect 29328 19264 29373 19292
rect 32048 19264 32229 19292
rect 29328 19252 29334 19264
rect 32217 19261 32229 19264
rect 32263 19261 32275 19295
rect 32217 19255 32275 19261
rect 32493 19295 32551 19301
rect 32493 19261 32505 19295
rect 32539 19292 32551 19295
rect 34146 19292 34152 19304
rect 32539 19264 34152 19292
rect 32539 19261 32551 19264
rect 32493 19255 32551 19261
rect 28442 19224 28448 19236
rect 21131 19196 21956 19224
rect 25608 19196 27200 19224
rect 28355 19196 28448 19224
rect 21131 19193 21143 19196
rect 21085 19187 21143 19193
rect 13173 19159 13231 19165
rect 13173 19125 13185 19159
rect 13219 19156 13231 19159
rect 13630 19156 13636 19168
rect 13219 19128 13636 19156
rect 13219 19125 13231 19128
rect 13173 19119 13231 19125
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 24394 19116 24400 19168
rect 24452 19156 24458 19168
rect 25608 19156 25636 19196
rect 27062 19156 27068 19168
rect 24452 19128 25636 19156
rect 27023 19128 27068 19156
rect 24452 19116 24458 19128
rect 27062 19116 27068 19128
rect 27120 19116 27126 19168
rect 27172 19156 27200 19196
rect 28442 19184 28448 19196
rect 28500 19224 28506 19236
rect 32508 19224 32536 19255
rect 34146 19252 34152 19264
rect 34204 19252 34210 19304
rect 35526 19252 35532 19304
rect 35584 19292 35590 19304
rect 37550 19292 37556 19304
rect 35584 19264 37556 19292
rect 35584 19252 35590 19264
rect 37550 19252 37556 19264
rect 37608 19252 37614 19304
rect 46661 19295 46719 19301
rect 46661 19261 46673 19295
rect 46707 19292 46719 19295
rect 46934 19292 46940 19304
rect 46707 19264 46940 19292
rect 46707 19261 46719 19264
rect 46661 19255 46719 19261
rect 46934 19252 46940 19264
rect 46992 19252 46998 19304
rect 33594 19224 33600 19236
rect 28500 19196 32536 19224
rect 33507 19196 33600 19224
rect 28500 19184 28506 19196
rect 33594 19184 33600 19196
rect 33652 19224 33658 19236
rect 35544 19224 35572 19252
rect 33652 19196 35572 19224
rect 33652 19184 33658 19196
rect 41322 19184 41328 19236
rect 41380 19224 41386 19236
rect 46109 19227 46167 19233
rect 46109 19224 46121 19227
rect 41380 19196 46121 19224
rect 41380 19184 41386 19196
rect 46109 19193 46121 19196
rect 46155 19224 46167 19227
rect 47026 19224 47032 19236
rect 46155 19196 47032 19224
rect 46155 19193 46167 19196
rect 46109 19187 46167 19193
rect 47026 19184 47032 19196
rect 47084 19184 47090 19236
rect 31386 19156 31392 19168
rect 27172 19128 31392 19156
rect 31386 19116 31392 19128
rect 31444 19116 31450 19168
rect 42794 19116 42800 19168
rect 42852 19156 42858 19168
rect 43165 19159 43223 19165
rect 43165 19156 43177 19159
rect 42852 19128 43177 19156
rect 42852 19116 42858 19128
rect 43165 19125 43177 19128
rect 43211 19125 43223 19159
rect 43165 19119 43223 19125
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 16942 18952 16948 18964
rect 2225 18915 2283 18921
rect 14476 18924 16528 18952
rect 16903 18924 16948 18952
rect 12710 18884 12716 18896
rect 11716 18856 12716 18884
rect 11716 18825 11744 18856
rect 12710 18844 12716 18856
rect 12768 18844 12774 18896
rect 11701 18819 11759 18825
rect 11701 18785 11713 18819
rect 11747 18785 11759 18819
rect 11701 18779 11759 18785
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12492 18788 12537 18816
rect 12492 18776 12498 18788
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 2188 18720 6914 18748
rect 2188 18708 2194 18720
rect 6886 18612 6914 18720
rect 11882 18680 11888 18692
rect 11843 18652 11888 18680
rect 11882 18640 11888 18652
rect 11940 18640 11946 18692
rect 13538 18612 13544 18624
rect 6886 18584 13544 18612
rect 13538 18572 13544 18584
rect 13596 18612 13602 18624
rect 14476 18612 14504 18924
rect 16500 18884 16528 18924
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 21453 18955 21511 18961
rect 21453 18921 21465 18955
rect 21499 18952 21511 18955
rect 21818 18952 21824 18964
rect 21499 18924 21824 18952
rect 21499 18921 21511 18924
rect 21453 18915 21511 18921
rect 21818 18912 21824 18924
rect 21876 18912 21882 18964
rect 23477 18955 23535 18961
rect 23477 18921 23489 18955
rect 23523 18952 23535 18955
rect 24578 18952 24584 18964
rect 23523 18924 24584 18952
rect 23523 18921 23535 18924
rect 23477 18915 23535 18921
rect 24578 18912 24584 18924
rect 24636 18912 24642 18964
rect 24854 18952 24860 18964
rect 24815 18924 24860 18952
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 27157 18955 27215 18961
rect 27157 18952 27169 18955
rect 24964 18924 27169 18952
rect 24394 18884 24400 18896
rect 16500 18856 24400 18884
rect 24394 18844 24400 18856
rect 24452 18844 24458 18896
rect 24762 18844 24768 18896
rect 24820 18884 24826 18896
rect 24964 18884 24992 18924
rect 27157 18921 27169 18924
rect 27203 18921 27215 18955
rect 33134 18952 33140 18964
rect 33095 18924 33140 18952
rect 27157 18915 27215 18921
rect 33134 18912 33140 18924
rect 33192 18912 33198 18964
rect 33410 18952 33416 18964
rect 33371 18924 33416 18952
rect 33410 18912 33416 18924
rect 33468 18912 33474 18964
rect 41138 18912 41144 18964
rect 41196 18952 41202 18964
rect 41196 18924 41414 18952
rect 41196 18912 41202 18924
rect 24820 18856 24992 18884
rect 24820 18844 24826 18856
rect 25406 18844 25412 18896
rect 25464 18844 25470 18896
rect 41386 18884 41414 18924
rect 47210 18912 47216 18964
rect 47268 18952 47274 18964
rect 48041 18955 48099 18961
rect 48041 18952 48053 18955
rect 47268 18924 48053 18952
rect 47268 18912 47274 18924
rect 48041 18921 48053 18924
rect 48087 18921 48099 18955
rect 48041 18915 48099 18921
rect 41386 18856 45508 18884
rect 15470 18816 15476 18828
rect 14752 18788 15476 18816
rect 14752 18757 14780 18788
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 23017 18819 23075 18825
rect 23017 18785 23029 18819
rect 23063 18816 23075 18819
rect 24302 18816 24308 18828
rect 23063 18788 24308 18816
rect 23063 18785 23075 18788
rect 23017 18779 23075 18785
rect 24302 18776 24308 18788
rect 24360 18776 24366 18828
rect 25424 18816 25452 18844
rect 25685 18819 25743 18825
rect 25685 18816 25697 18819
rect 25424 18788 25697 18816
rect 25685 18785 25697 18788
rect 25731 18785 25743 18819
rect 25685 18779 25743 18785
rect 28534 18776 28540 18828
rect 28592 18816 28598 18828
rect 29641 18819 29699 18825
rect 29641 18816 29653 18819
rect 28592 18788 29653 18816
rect 28592 18776 28598 18788
rect 29641 18785 29653 18788
rect 29687 18785 29699 18819
rect 29641 18779 29699 18785
rect 30101 18819 30159 18825
rect 30101 18785 30113 18819
rect 30147 18816 30159 18819
rect 30374 18816 30380 18828
rect 30147 18788 30380 18816
rect 30147 18785 30159 18788
rect 30101 18779 30159 18785
rect 30374 18776 30380 18788
rect 30432 18776 30438 18828
rect 42794 18816 42800 18828
rect 42755 18788 42800 18816
rect 42794 18776 42800 18788
rect 42852 18776 42858 18828
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 15194 18748 15200 18760
rect 15155 18720 15200 18748
rect 14737 18711 14795 18717
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18748 21511 18751
rect 22002 18748 22008 18760
rect 21499 18720 22008 18748
rect 21499 18717 21511 18720
rect 21453 18711 21511 18717
rect 22002 18708 22008 18720
rect 22060 18748 22066 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22060 18720 22937 18748
rect 22060 18708 22066 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 23474 18748 23480 18760
rect 23435 18720 23480 18748
rect 22925 18711 22983 18717
rect 15473 18683 15531 18689
rect 15473 18649 15485 18683
rect 15519 18649 15531 18683
rect 16758 18680 16764 18692
rect 16698 18652 16764 18680
rect 15473 18643 15531 18649
rect 13596 18584 14504 18612
rect 14553 18615 14611 18621
rect 13596 18572 13602 18584
rect 14553 18581 14565 18615
rect 14599 18612 14611 18615
rect 15488 18612 15516 18643
rect 16758 18640 16764 18652
rect 16816 18640 16822 18692
rect 22940 18680 22968 18711
rect 23474 18708 23480 18720
rect 23532 18708 23538 18760
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 23842 18748 23848 18760
rect 23707 18720 23848 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24670 18680 24676 18692
rect 22940 18652 24676 18680
rect 24670 18640 24676 18652
rect 24728 18640 24734 18692
rect 14599 18584 15516 18612
rect 24780 18612 24808 18711
rect 25314 18708 25320 18760
rect 25372 18748 25378 18760
rect 25409 18751 25467 18757
rect 25409 18748 25421 18751
rect 25372 18720 25421 18748
rect 25372 18708 25378 18720
rect 25409 18717 25421 18720
rect 25455 18717 25467 18751
rect 28442 18748 28448 18760
rect 28403 18720 28448 18748
rect 25409 18711 25467 18717
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 28626 18748 28632 18760
rect 28587 18720 28632 18748
rect 28626 18708 28632 18720
rect 28684 18708 28690 18760
rect 29733 18751 29791 18757
rect 29733 18717 29745 18751
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 27062 18680 27068 18692
rect 26910 18652 27068 18680
rect 27062 18640 27068 18652
rect 27120 18640 27126 18692
rect 28537 18683 28595 18689
rect 28537 18649 28549 18683
rect 28583 18680 28595 18683
rect 29270 18680 29276 18692
rect 28583 18652 29276 18680
rect 28583 18649 28595 18652
rect 28537 18643 28595 18649
rect 29270 18640 29276 18652
rect 29328 18680 29334 18692
rect 29748 18680 29776 18711
rect 29914 18708 29920 18760
rect 29972 18748 29978 18760
rect 30653 18751 30711 18757
rect 30653 18748 30665 18751
rect 29972 18720 30665 18748
rect 29972 18708 29978 18720
rect 30653 18717 30665 18720
rect 30699 18717 30711 18751
rect 30653 18711 30711 18717
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32953 18751 33011 18757
rect 32953 18748 32965 18751
rect 32272 18720 32965 18748
rect 32272 18708 32278 18720
rect 32953 18717 32965 18720
rect 32999 18717 33011 18751
rect 32953 18711 33011 18717
rect 42613 18751 42671 18757
rect 42613 18717 42625 18751
rect 42659 18717 42671 18751
rect 45186 18748 45192 18760
rect 45147 18720 45192 18748
rect 42613 18711 42671 18717
rect 29328 18652 29776 18680
rect 30837 18683 30895 18689
rect 29328 18640 29334 18652
rect 30837 18649 30849 18683
rect 30883 18680 30895 18683
rect 32030 18680 32036 18692
rect 30883 18652 32036 18680
rect 30883 18649 30895 18652
rect 30837 18643 30895 18649
rect 32030 18640 32036 18652
rect 32088 18640 32094 18692
rect 32122 18640 32128 18692
rect 32180 18680 32186 18692
rect 32493 18683 32551 18689
rect 32493 18680 32505 18683
rect 32180 18652 32505 18680
rect 32180 18640 32186 18652
rect 32493 18649 32505 18652
rect 32539 18680 32551 18683
rect 32858 18680 32864 18692
rect 32539 18652 32864 18680
rect 32539 18649 32551 18652
rect 32493 18643 32551 18649
rect 32858 18640 32864 18652
rect 32916 18640 32922 18692
rect 42628 18680 42656 18711
rect 45186 18708 45192 18720
rect 45244 18708 45250 18760
rect 45370 18748 45376 18760
rect 45331 18720 45376 18748
rect 45370 18708 45376 18720
rect 45428 18708 45434 18760
rect 45480 18748 45508 18856
rect 45833 18819 45891 18825
rect 45833 18785 45845 18819
rect 45879 18816 45891 18819
rect 47118 18816 47124 18828
rect 45879 18788 47124 18816
rect 45879 18785 45891 18788
rect 45833 18779 45891 18785
rect 47118 18776 47124 18788
rect 47176 18776 47182 18828
rect 46198 18748 46204 18760
rect 45480 18720 46204 18748
rect 46198 18708 46204 18720
rect 46256 18708 46262 18760
rect 46382 18708 46388 18760
rect 46440 18748 46446 18760
rect 46477 18751 46535 18757
rect 46477 18748 46489 18751
rect 46440 18720 46489 18748
rect 46440 18708 46446 18720
rect 46477 18717 46489 18720
rect 46523 18717 46535 18751
rect 46477 18711 46535 18717
rect 46845 18751 46903 18757
rect 46845 18717 46857 18751
rect 46891 18748 46903 18751
rect 47026 18748 47032 18760
rect 46891 18720 47032 18748
rect 46891 18717 46903 18720
rect 46845 18711 46903 18717
rect 47026 18708 47032 18720
rect 47084 18708 47090 18760
rect 47302 18748 47308 18760
rect 47263 18720 47308 18748
rect 47302 18708 47308 18720
rect 47360 18708 47366 18760
rect 47949 18751 48007 18757
rect 47949 18717 47961 18751
rect 47995 18748 48007 18751
rect 48038 18748 48044 18760
rect 47995 18720 48044 18748
rect 47995 18717 48007 18720
rect 47949 18711 48007 18717
rect 48038 18708 48044 18720
rect 48096 18708 48102 18760
rect 44082 18680 44088 18692
rect 42628 18652 44088 18680
rect 44082 18640 44088 18652
rect 44140 18640 44146 18692
rect 44450 18680 44456 18692
rect 44411 18652 44456 18680
rect 44450 18640 44456 18652
rect 44508 18640 44514 18692
rect 46106 18680 46112 18692
rect 46067 18652 46112 18680
rect 46106 18640 46112 18652
rect 46164 18640 46170 18692
rect 26418 18612 26424 18624
rect 24780 18584 26424 18612
rect 14599 18581 14611 18584
rect 14553 18575 14611 18581
rect 26418 18572 26424 18584
rect 26476 18572 26482 18624
rect 44358 18572 44364 18624
rect 44416 18612 44422 18624
rect 45281 18615 45339 18621
rect 45281 18612 45293 18615
rect 44416 18584 45293 18612
rect 44416 18572 44422 18584
rect 45281 18581 45293 18584
rect 45327 18581 45339 18615
rect 45281 18575 45339 18581
rect 46474 18572 46480 18624
rect 46532 18612 46538 18624
rect 47397 18615 47455 18621
rect 47397 18612 47409 18615
rect 46532 18584 47409 18612
rect 46532 18572 46538 18584
rect 47397 18581 47409 18584
rect 47443 18581 47455 18615
rect 47397 18575 47455 18581
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 44818 18408 44824 18420
rect 3476 18380 31064 18408
rect 3476 18368 3482 18380
rect 11882 18340 11888 18352
rect 11843 18312 11888 18340
rect 11882 18300 11888 18312
rect 11940 18300 11946 18352
rect 13630 18340 13636 18352
rect 13591 18312 13636 18340
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 14366 18300 14372 18352
rect 14424 18300 14430 18352
rect 15194 18300 15200 18352
rect 15252 18340 15258 18352
rect 15933 18343 15991 18349
rect 15933 18340 15945 18343
rect 15252 18312 15945 18340
rect 15252 18300 15258 18312
rect 15933 18309 15945 18312
rect 15979 18309 15991 18343
rect 16758 18340 16764 18352
rect 16719 18312 16764 18340
rect 15933 18303 15991 18309
rect 16758 18300 16764 18312
rect 16816 18300 16822 18352
rect 18598 18300 18604 18352
rect 18656 18300 18662 18352
rect 22833 18343 22891 18349
rect 22833 18309 22845 18343
rect 22879 18340 22891 18343
rect 23569 18343 23627 18349
rect 23569 18340 23581 18343
rect 22879 18312 23581 18340
rect 22879 18309 22891 18312
rect 22833 18303 22891 18309
rect 23569 18309 23581 18312
rect 23615 18309 23627 18343
rect 27982 18340 27988 18352
rect 23569 18303 23627 18309
rect 27908 18312 27988 18340
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 11790 18272 11796 18284
rect 11751 18244 11796 18272
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 15654 18272 15660 18284
rect 15615 18244 15660 18272
rect 15654 18232 15660 18244
rect 15712 18232 15718 18284
rect 16666 18272 16672 18284
rect 16627 18244 16672 18272
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 22741 18275 22799 18281
rect 22741 18241 22753 18275
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18272 27675 18275
rect 27706 18272 27712 18284
rect 27663 18244 27712 18272
rect 27663 18241 27675 18244
rect 27617 18235 27675 18241
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18204 13415 18207
rect 13998 18204 14004 18216
rect 13403 18176 14004 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 13998 18164 14004 18176
rect 14056 18164 14062 18216
rect 17678 18204 17684 18216
rect 17639 18176 17684 18204
rect 17678 18164 17684 18176
rect 17736 18164 17742 18216
rect 17957 18207 18015 18213
rect 17957 18173 17969 18207
rect 18003 18204 18015 18207
rect 19794 18204 19800 18216
rect 18003 18176 19800 18204
rect 18003 18173 18015 18176
rect 17957 18167 18015 18173
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 15378 18136 15384 18148
rect 14660 18108 15384 18136
rect 1949 18071 2007 18077
rect 1949 18037 1961 18071
rect 1995 18068 2007 18071
rect 14660 18068 14688 18108
rect 15378 18096 15384 18108
rect 15436 18096 15442 18148
rect 19426 18136 19432 18148
rect 19387 18108 19432 18136
rect 19426 18096 19432 18108
rect 19484 18096 19490 18148
rect 22756 18136 22784 18235
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 27908 18281 27936 18312
rect 27982 18300 27988 18312
rect 28040 18300 28046 18352
rect 28074 18300 28080 18352
rect 28132 18340 28138 18352
rect 31036 18340 31064 18380
rect 31864 18380 44824 18408
rect 28132 18312 28225 18340
rect 31036 18312 31156 18340
rect 28132 18300 28138 18312
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18241 27951 18275
rect 28092 18272 28120 18300
rect 28721 18275 28779 18281
rect 28721 18272 28733 18275
rect 28092 18244 28733 18272
rect 27893 18235 27951 18241
rect 28721 18241 28733 18244
rect 28767 18241 28779 18275
rect 28721 18235 28779 18241
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 24762 18204 24768 18216
rect 23431 18176 24768 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25314 18204 25320 18216
rect 25271 18176 25320 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 27985 18207 28043 18213
rect 27985 18173 27997 18207
rect 28031 18173 28043 18207
rect 27985 18167 28043 18173
rect 23014 18136 23020 18148
rect 22756 18108 23020 18136
rect 23014 18096 23020 18108
rect 23072 18136 23078 18148
rect 28000 18136 28028 18167
rect 28166 18164 28172 18216
rect 28224 18204 28230 18216
rect 28537 18207 28595 18213
rect 28537 18204 28549 18207
rect 28224 18176 28549 18204
rect 28224 18164 28230 18176
rect 28537 18173 28549 18176
rect 28583 18173 28595 18207
rect 28537 18167 28595 18173
rect 29733 18207 29791 18213
rect 29733 18173 29745 18207
rect 29779 18173 29791 18207
rect 29914 18204 29920 18216
rect 29875 18176 29920 18204
rect 29733 18167 29791 18173
rect 28442 18136 28448 18148
rect 23072 18108 27936 18136
rect 28000 18108 28448 18136
rect 23072 18096 23078 18108
rect 1995 18040 14688 18068
rect 1995 18037 2007 18040
rect 1949 18031 2007 18037
rect 14918 18028 14924 18080
rect 14976 18068 14982 18080
rect 15102 18068 15108 18080
rect 14976 18040 15108 18068
rect 14976 18028 14982 18040
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 27709 18071 27767 18077
rect 27709 18037 27721 18071
rect 27755 18068 27767 18071
rect 27798 18068 27804 18080
rect 27755 18040 27804 18068
rect 27755 18037 27767 18040
rect 27709 18031 27767 18037
rect 27798 18028 27804 18040
rect 27856 18028 27862 18080
rect 27908 18068 27936 18108
rect 28442 18096 28448 18108
rect 28500 18096 28506 18148
rect 29748 18136 29776 18167
rect 29914 18164 29920 18176
rect 29972 18164 29978 18216
rect 31128 18213 31156 18312
rect 31113 18207 31171 18213
rect 31113 18173 31125 18207
rect 31159 18173 31171 18207
rect 31113 18167 31171 18173
rect 30374 18136 30380 18148
rect 28552 18108 29684 18136
rect 29748 18108 30380 18136
rect 28552 18068 28580 18108
rect 27908 18040 28580 18068
rect 28905 18071 28963 18077
rect 28905 18037 28917 18071
rect 28951 18068 28963 18071
rect 29178 18068 29184 18080
rect 28951 18040 29184 18068
rect 28951 18037 28963 18040
rect 28905 18031 28963 18037
rect 29178 18028 29184 18040
rect 29236 18028 29242 18080
rect 29656 18068 29684 18108
rect 30374 18096 30380 18108
rect 30432 18136 30438 18148
rect 31018 18136 31024 18148
rect 30432 18108 31024 18136
rect 30432 18096 30438 18108
rect 31018 18096 31024 18108
rect 31076 18096 31082 18148
rect 31864 18068 31892 18380
rect 44818 18368 44824 18380
rect 44876 18368 44882 18420
rect 45186 18368 45192 18420
rect 45244 18408 45250 18420
rect 47949 18411 48007 18417
rect 47949 18408 47961 18411
rect 45244 18380 47961 18408
rect 45244 18368 45250 18380
rect 47949 18377 47961 18380
rect 47995 18377 48007 18411
rect 47949 18371 48007 18377
rect 32214 18300 32220 18352
rect 32272 18340 32278 18352
rect 41322 18340 41328 18352
rect 32272 18312 41328 18340
rect 32272 18300 32278 18312
rect 41322 18300 41328 18312
rect 41380 18340 41386 18352
rect 45373 18343 45431 18349
rect 41380 18312 41460 18340
rect 41380 18300 41386 18312
rect 32030 18232 32036 18284
rect 32088 18272 32094 18284
rect 32125 18275 32183 18281
rect 32125 18272 32137 18275
rect 32088 18244 32137 18272
rect 32088 18232 32094 18244
rect 32125 18241 32137 18244
rect 32171 18272 32183 18275
rect 33229 18275 33287 18281
rect 32171 18244 32536 18272
rect 32171 18241 32183 18244
rect 32125 18235 32183 18241
rect 32508 18136 32536 18244
rect 33229 18241 33241 18275
rect 33275 18241 33287 18275
rect 33229 18235 33287 18241
rect 32585 18207 32643 18213
rect 32585 18173 32597 18207
rect 32631 18204 32643 18207
rect 33244 18204 33272 18235
rect 41138 18232 41144 18284
rect 41196 18272 41202 18284
rect 41432 18281 41460 18312
rect 45373 18309 45385 18343
rect 45419 18340 45431 18343
rect 46106 18340 46112 18352
rect 45419 18312 46112 18340
rect 45419 18309 45431 18312
rect 45373 18303 45431 18309
rect 46106 18300 46112 18312
rect 46164 18300 46170 18352
rect 47486 18300 47492 18352
rect 47544 18340 47550 18352
rect 47765 18343 47823 18349
rect 47765 18340 47777 18343
rect 47544 18312 47777 18340
rect 47544 18300 47550 18312
rect 47765 18309 47777 18312
rect 47811 18309 47823 18343
rect 47765 18303 47823 18309
rect 44364 18284 44416 18290
rect 41233 18275 41291 18281
rect 41233 18272 41245 18275
rect 41196 18244 41245 18272
rect 41196 18232 41202 18244
rect 41233 18241 41245 18244
rect 41279 18241 41291 18275
rect 41233 18235 41291 18241
rect 41417 18275 41475 18281
rect 41417 18241 41429 18275
rect 41463 18241 41475 18275
rect 41417 18235 41475 18241
rect 41693 18275 41751 18281
rect 41693 18241 41705 18275
rect 41739 18241 41751 18275
rect 43714 18272 43720 18284
rect 43675 18244 43720 18272
rect 41693 18235 41751 18241
rect 41708 18204 41736 18235
rect 43714 18232 43720 18244
rect 43772 18232 43778 18284
rect 46750 18232 46756 18284
rect 46808 18272 46814 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 46808 18244 47593 18272
rect 46808 18232 46814 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 44364 18226 44416 18232
rect 44637 18207 44695 18213
rect 32631 18176 33272 18204
rect 41386 18176 43944 18204
rect 32631 18173 32643 18176
rect 32585 18167 32643 18173
rect 41386 18136 41414 18176
rect 41598 18136 41604 18148
rect 32508 18108 41414 18136
rect 41559 18108 41604 18136
rect 41598 18096 41604 18108
rect 41656 18096 41662 18148
rect 32214 18068 32220 18080
rect 29656 18040 31892 18068
rect 32175 18040 32220 18068
rect 32214 18028 32220 18040
rect 32272 18028 32278 18080
rect 32398 18028 32404 18080
rect 32456 18068 32462 18080
rect 33045 18071 33103 18077
rect 33045 18068 33057 18071
rect 32456 18040 33057 18068
rect 32456 18028 32462 18040
rect 33045 18037 33057 18040
rect 33091 18037 33103 18071
rect 43916 18068 43944 18176
rect 44637 18173 44649 18207
rect 44683 18204 44695 18207
rect 45189 18207 45247 18213
rect 45189 18204 45201 18207
rect 44683 18176 45201 18204
rect 44683 18173 44695 18176
rect 44637 18167 44695 18173
rect 45189 18173 45201 18176
rect 45235 18173 45247 18207
rect 45646 18204 45652 18216
rect 45607 18176 45652 18204
rect 45189 18167 45247 18173
rect 44358 18096 44364 18148
rect 44416 18136 44422 18148
rect 44652 18136 44680 18167
rect 45646 18164 45652 18176
rect 45704 18164 45710 18216
rect 44416 18108 44680 18136
rect 44416 18096 44422 18108
rect 46382 18068 46388 18080
rect 43916 18040 46388 18068
rect 33045 18031 33103 18037
rect 46382 18028 46388 18040
rect 46440 18028 46446 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 12434 17864 12440 17876
rect 3108 17836 12440 17864
rect 3108 17824 3114 17836
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 14366 17864 14372 17876
rect 14327 17836 14372 17864
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 17497 17867 17555 17873
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 17678 17864 17684 17876
rect 17543 17836 17684 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 18598 17864 18604 17876
rect 18559 17836 18604 17864
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 19794 17864 19800 17876
rect 19755 17836 19800 17864
rect 19794 17824 19800 17836
rect 19852 17824 19858 17876
rect 23106 17824 23112 17876
rect 23164 17864 23170 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 23164 17836 23305 17864
rect 23164 17824 23170 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 29914 17824 29920 17876
rect 29972 17864 29978 17876
rect 30193 17867 30251 17873
rect 30193 17864 30205 17867
rect 29972 17836 30205 17864
rect 29972 17824 29978 17836
rect 30193 17833 30205 17836
rect 30239 17833 30251 17867
rect 42610 17864 42616 17876
rect 30193 17827 30251 17833
rect 31726 17836 42616 17864
rect 12802 17796 12808 17808
rect 11716 17768 12808 17796
rect 11716 17737 11744 17768
rect 12802 17756 12808 17768
rect 12860 17796 12866 17808
rect 15102 17796 15108 17808
rect 12860 17768 15108 17796
rect 12860 17756 12866 17768
rect 15102 17756 15108 17768
rect 15160 17756 15166 17808
rect 24026 17756 24032 17808
rect 24084 17796 24090 17808
rect 31726 17796 31754 17836
rect 42610 17824 42616 17836
rect 42668 17824 42674 17876
rect 44174 17824 44180 17876
rect 44232 17864 44238 17876
rect 45649 17867 45707 17873
rect 45649 17864 45661 17867
rect 44232 17836 45661 17864
rect 44232 17824 44238 17836
rect 45649 17833 45661 17836
rect 45695 17833 45707 17867
rect 45649 17827 45707 17833
rect 24084 17768 31754 17796
rect 24084 17756 24090 17768
rect 36538 17756 36544 17808
rect 36596 17796 36602 17808
rect 36596 17768 44128 17796
rect 36596 17756 36602 17768
rect 11701 17731 11759 17737
rect 11701 17697 11713 17731
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 16666 17728 16672 17740
rect 12492 17700 12537 17728
rect 14292 17700 16672 17728
rect 12492 17688 12498 17700
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 14292 17669 14320 17700
rect 16666 17688 16672 17700
rect 16724 17688 16730 17740
rect 18690 17688 18696 17740
rect 18748 17728 18754 17740
rect 19337 17731 19395 17737
rect 19337 17728 19349 17731
rect 18748 17700 19349 17728
rect 18748 17688 18754 17700
rect 19337 17697 19349 17700
rect 19383 17697 19395 17731
rect 38746 17728 38752 17740
rect 19337 17691 19395 17697
rect 30116 17700 38752 17728
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 13780 17632 14289 17660
rect 13780 17620 13786 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 16574 17660 16580 17672
rect 15712 17632 16580 17660
rect 15712 17620 15718 17632
rect 16574 17620 16580 17632
rect 16632 17660 16638 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 16632 17632 17325 17660
rect 16632 17620 16638 17632
rect 17313 17629 17325 17632
rect 17359 17660 17371 17663
rect 17494 17660 17500 17672
rect 17359 17632 17500 17660
rect 17359 17629 17371 17632
rect 17313 17623 17371 17629
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 19150 17660 19156 17672
rect 18555 17632 19156 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 19150 17620 19156 17632
rect 19208 17620 19214 17672
rect 19426 17660 19432 17672
rect 19387 17632 19432 17660
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 20438 17620 20444 17672
rect 20496 17660 20502 17672
rect 20533 17663 20591 17669
rect 20533 17660 20545 17663
rect 20496 17632 20545 17660
rect 20496 17620 20502 17632
rect 20533 17629 20545 17632
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17660 27123 17663
rect 27798 17660 27804 17672
rect 27111 17632 27804 17660
rect 27111 17629 27123 17632
rect 27065 17623 27123 17629
rect 27798 17620 27804 17632
rect 27856 17620 27862 17672
rect 30116 17669 30144 17700
rect 38746 17688 38752 17700
rect 38804 17688 38810 17740
rect 41414 17688 41420 17740
rect 41472 17728 41478 17740
rect 41598 17728 41604 17740
rect 41472 17700 41517 17728
rect 41559 17700 41604 17728
rect 41472 17688 41478 17700
rect 41598 17688 41604 17700
rect 41656 17688 41662 17740
rect 41874 17728 41880 17740
rect 41835 17700 41880 17728
rect 41874 17688 41880 17700
rect 41932 17688 41938 17740
rect 27893 17663 27951 17669
rect 27893 17629 27905 17663
rect 27939 17660 27951 17663
rect 30101 17663 30159 17669
rect 27939 17632 29868 17660
rect 27939 17629 27951 17632
rect 27893 17623 27951 17629
rect 11882 17592 11888 17604
rect 11843 17564 11888 17592
rect 11882 17552 11888 17564
rect 11940 17552 11946 17604
rect 23109 17595 23167 17601
rect 23109 17561 23121 17595
rect 23155 17592 23167 17595
rect 23198 17592 23204 17604
rect 23155 17564 23204 17592
rect 23155 17561 23167 17564
rect 23109 17555 23167 17561
rect 23198 17552 23204 17564
rect 23256 17552 23262 17604
rect 23325 17595 23383 17601
rect 23325 17561 23337 17595
rect 23371 17592 23383 17595
rect 23842 17592 23848 17604
rect 23371 17564 23848 17592
rect 23371 17561 23383 17564
rect 23325 17555 23383 17561
rect 23842 17552 23848 17564
rect 23900 17552 23906 17604
rect 27249 17595 27307 17601
rect 27249 17561 27261 17595
rect 27295 17592 27307 17595
rect 27338 17592 27344 17604
rect 27295 17564 27344 17592
rect 27295 17561 27307 17564
rect 27249 17555 27307 17561
rect 27338 17552 27344 17564
rect 27396 17592 27402 17604
rect 27706 17592 27712 17604
rect 27396 17564 27712 17592
rect 27396 17552 27402 17564
rect 27706 17552 27712 17564
rect 27764 17552 27770 17604
rect 28074 17592 28080 17604
rect 28035 17564 28080 17592
rect 28074 17552 28080 17564
rect 28132 17552 28138 17604
rect 28442 17592 28448 17604
rect 28403 17564 28448 17592
rect 28442 17552 28448 17564
rect 28500 17552 28506 17604
rect 17310 17484 17316 17536
rect 17368 17524 17374 17536
rect 20162 17524 20168 17536
rect 17368 17496 20168 17524
rect 17368 17484 17374 17496
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 20625 17527 20683 17533
rect 20625 17493 20637 17527
rect 20671 17524 20683 17527
rect 20806 17524 20812 17536
rect 20671 17496 20812 17524
rect 20671 17493 20683 17496
rect 20625 17487 20683 17493
rect 20806 17484 20812 17496
rect 20864 17484 20870 17536
rect 23474 17524 23480 17536
rect 23435 17496 23480 17524
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 27433 17527 27491 17533
rect 27433 17493 27445 17527
rect 27479 17524 27491 17527
rect 27890 17524 27896 17536
rect 27479 17496 27896 17524
rect 27479 17493 27491 17496
rect 27433 17487 27491 17493
rect 27890 17484 27896 17496
rect 27948 17484 27954 17536
rect 28166 17524 28172 17536
rect 28127 17496 28172 17524
rect 28166 17484 28172 17496
rect 28224 17484 28230 17536
rect 28258 17484 28264 17536
rect 28316 17524 28322 17536
rect 29840 17524 29868 17632
rect 30101 17629 30113 17663
rect 30147 17629 30159 17663
rect 31018 17660 31024 17672
rect 30979 17632 31024 17660
rect 30101 17623 30159 17629
rect 31018 17620 31024 17632
rect 31076 17620 31082 17672
rect 44100 17669 44128 17768
rect 45005 17731 45063 17737
rect 45005 17697 45017 17731
rect 45051 17728 45063 17731
rect 45186 17728 45192 17740
rect 45051 17700 45192 17728
rect 45051 17697 45063 17700
rect 45005 17691 45063 17697
rect 45186 17688 45192 17700
rect 45244 17688 45250 17740
rect 46293 17731 46351 17737
rect 46293 17697 46305 17731
rect 46339 17728 46351 17731
rect 47486 17728 47492 17740
rect 46339 17700 47492 17728
rect 46339 17697 46351 17700
rect 46293 17691 46351 17697
rect 47486 17688 47492 17700
rect 47544 17688 47550 17740
rect 44085 17663 44143 17669
rect 44085 17629 44097 17663
rect 44131 17629 44143 17663
rect 45370 17660 45376 17672
rect 45331 17632 45376 17660
rect 44085 17623 44143 17629
rect 45370 17620 45376 17632
rect 45428 17620 45434 17672
rect 45465 17663 45523 17669
rect 45465 17629 45477 17663
rect 45511 17629 45523 17663
rect 45465 17623 45523 17629
rect 31205 17595 31263 17601
rect 31205 17561 31217 17595
rect 31251 17592 31263 17595
rect 32398 17592 32404 17604
rect 31251 17564 32404 17592
rect 31251 17561 31263 17564
rect 31205 17555 31263 17561
rect 32398 17552 32404 17564
rect 32456 17552 32462 17604
rect 32858 17592 32864 17604
rect 32819 17564 32864 17592
rect 32858 17552 32864 17564
rect 32916 17552 32922 17604
rect 45480 17592 45508 17623
rect 43732 17564 45508 17592
rect 46477 17595 46535 17601
rect 43732 17536 43760 17564
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 47670 17592 47676 17604
rect 46523 17564 47676 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 47670 17552 47676 17564
rect 47728 17552 47734 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 43714 17524 43720 17536
rect 28316 17496 28361 17524
rect 29840 17496 43720 17524
rect 28316 17484 28322 17496
rect 43714 17484 43720 17496
rect 43772 17484 43778 17536
rect 44177 17527 44235 17533
rect 44177 17493 44189 17527
rect 44223 17524 44235 17527
rect 44266 17524 44272 17536
rect 44223 17496 44272 17524
rect 44223 17493 44235 17496
rect 44177 17487 44235 17493
rect 44266 17484 44272 17496
rect 44324 17484 44330 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 4706 17280 4712 17332
rect 4764 17320 4770 17332
rect 11882 17320 11888 17332
rect 4764 17292 6914 17320
rect 11843 17292 11888 17320
rect 4764 17280 4770 17292
rect 6886 17252 6914 17292
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 27249 17323 27307 17329
rect 12406 17292 27108 17320
rect 12406 17252 12434 17292
rect 13998 17252 14004 17264
rect 6886 17224 12434 17252
rect 13959 17224 14004 17252
rect 13998 17212 14004 17224
rect 14056 17212 14062 17264
rect 19426 17212 19432 17264
rect 19484 17212 19490 17264
rect 20346 17252 20352 17264
rect 20307 17224 20352 17252
rect 20346 17212 20352 17224
rect 20404 17212 20410 17264
rect 20565 17255 20623 17261
rect 20565 17221 20577 17255
rect 20611 17252 20623 17255
rect 20714 17252 20720 17264
rect 20611 17224 20720 17252
rect 20611 17221 20623 17224
rect 20565 17215 20623 17221
rect 20714 17212 20720 17224
rect 20772 17252 20778 17264
rect 20990 17252 20996 17264
rect 20772 17224 20996 17252
rect 20772 17212 20778 17224
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 22554 17212 22560 17264
rect 22612 17212 22618 17264
rect 27080 17196 27108 17292
rect 27249 17289 27261 17323
rect 27295 17320 27307 17323
rect 28258 17320 28264 17332
rect 27295 17292 28264 17320
rect 27295 17289 27307 17292
rect 27249 17283 27307 17289
rect 28258 17280 28264 17292
rect 28316 17280 28322 17332
rect 29730 17280 29736 17332
rect 29788 17320 29794 17332
rect 36538 17320 36544 17332
rect 29788 17292 36544 17320
rect 29788 17280 29794 17292
rect 36538 17280 36544 17292
rect 36596 17280 36602 17332
rect 41892 17292 45324 17320
rect 41892 17264 41920 17292
rect 28442 17252 28448 17264
rect 28092 17224 28448 17252
rect 28092 17196 28120 17224
rect 28442 17212 28448 17224
rect 28500 17212 28506 17264
rect 32858 17212 32864 17264
rect 32916 17252 32922 17264
rect 41874 17252 41880 17264
rect 32916 17224 41880 17252
rect 32916 17212 32922 17224
rect 41874 17212 41880 17224
rect 41932 17212 41938 17264
rect 44266 17252 44272 17264
rect 44227 17224 44272 17252
rect 44266 17212 44272 17224
rect 44324 17212 44330 17264
rect 45296 17252 45324 17292
rect 45370 17280 45376 17332
rect 45428 17320 45434 17332
rect 46845 17323 46903 17329
rect 46845 17320 46857 17323
rect 45428 17292 46857 17320
rect 45428 17280 45434 17292
rect 46845 17289 46857 17292
rect 46891 17289 46903 17323
rect 47670 17320 47676 17332
rect 47631 17292 47676 17320
rect 46845 17283 46903 17289
rect 47670 17280 47676 17292
rect 47728 17280 47734 17332
rect 45646 17252 45652 17264
rect 45296 17224 45652 17252
rect 45646 17212 45652 17224
rect 45704 17212 45710 17264
rect 11790 17184 11796 17196
rect 11751 17156 11796 17184
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 13909 17187 13967 17193
rect 13909 17153 13921 17187
rect 13955 17184 13967 17187
rect 15654 17184 15660 17196
rect 13955 17156 15660 17184
rect 13955 17153 13967 17156
rect 13909 17147 13967 17153
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 15930 17184 15936 17196
rect 15887 17156 15936 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 17494 17184 17500 17196
rect 17455 17156 17500 17184
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17184 24271 17187
rect 24670 17184 24676 17196
rect 24259 17156 24676 17184
rect 24259 17153 24271 17156
rect 24213 17147 24271 17153
rect 24670 17144 24676 17156
rect 24728 17184 24734 17196
rect 25225 17187 25283 17193
rect 25225 17184 25237 17187
rect 24728 17156 25237 17184
rect 24728 17144 24734 17156
rect 25225 17153 25237 17156
rect 25271 17153 25283 17187
rect 25225 17147 25283 17153
rect 25961 17187 26019 17193
rect 25961 17153 25973 17187
rect 26007 17184 26019 17187
rect 26418 17184 26424 17196
rect 26007 17156 26424 17184
rect 26007 17153 26019 17156
rect 25961 17147 26019 17153
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 27062 17184 27068 17196
rect 26975 17156 27068 17184
rect 27062 17144 27068 17156
rect 27120 17144 27126 17196
rect 27154 17144 27160 17196
rect 27212 17184 27218 17196
rect 27249 17187 27307 17193
rect 27249 17184 27261 17187
rect 27212 17156 27261 17184
rect 27212 17144 27218 17156
rect 27249 17153 27261 17156
rect 27295 17153 27307 17187
rect 27982 17184 27988 17196
rect 27943 17156 27988 17184
rect 27249 17147 27307 17153
rect 27982 17144 27988 17156
rect 28040 17144 28046 17196
rect 28074 17144 28080 17196
rect 28132 17184 28138 17196
rect 28261 17187 28319 17193
rect 28132 17156 28177 17184
rect 28132 17144 28138 17156
rect 28261 17153 28273 17187
rect 28307 17184 28319 17187
rect 28813 17187 28871 17193
rect 28813 17184 28825 17187
rect 28307 17156 28825 17184
rect 28307 17153 28319 17156
rect 28261 17147 28319 17153
rect 28813 17153 28825 17156
rect 28859 17153 28871 17187
rect 29178 17184 29184 17196
rect 29139 17156 29184 17184
rect 28813 17147 28871 17153
rect 29178 17144 29184 17156
rect 29236 17144 29242 17196
rect 46750 17184 46756 17196
rect 46711 17156 46756 17184
rect 46750 17144 46756 17156
rect 46808 17144 46814 17196
rect 46937 17187 46995 17193
rect 46937 17153 46949 17187
rect 46983 17184 46995 17187
rect 47394 17184 47400 17196
rect 46983 17156 47400 17184
rect 46983 17153 46995 17156
rect 46937 17147 46995 17153
rect 47394 17144 47400 17156
rect 47452 17144 47458 17196
rect 47581 17187 47639 17193
rect 47581 17153 47593 17187
rect 47627 17184 47639 17187
rect 47670 17184 47676 17196
rect 47627 17156 47676 17184
rect 47627 17153 47639 17156
rect 47581 17147 47639 17153
rect 47670 17144 47676 17156
rect 47728 17144 47734 17196
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17116 17647 17119
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17635 17088 18153 17116
rect 17635 17085 17647 17088
rect 17589 17079 17647 17085
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17116 18475 17119
rect 18506 17116 18512 17128
rect 18463 17088 18512 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 18782 17076 18788 17128
rect 18840 17116 18846 17128
rect 21818 17116 21824 17128
rect 18840 17088 20760 17116
rect 21779 17088 21824 17116
rect 18840 17076 18846 17088
rect 19518 17008 19524 17060
rect 19576 17048 19582 17060
rect 19889 17051 19947 17057
rect 19889 17048 19901 17051
rect 19576 17020 19901 17048
rect 19576 17008 19582 17020
rect 19889 17017 19901 17020
rect 19935 17048 19947 17051
rect 20346 17048 20352 17060
rect 19935 17020 20352 17048
rect 19935 17017 19947 17020
rect 19889 17011 19947 17017
rect 20346 17008 20352 17020
rect 20404 17008 20410 17060
rect 20732 17057 20760 17088
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 44085 17119 44143 17125
rect 22152 17088 22197 17116
rect 22152 17076 22158 17088
rect 44085 17085 44097 17119
rect 44131 17116 44143 17119
rect 44358 17116 44364 17128
rect 44131 17088 44364 17116
rect 44131 17085 44143 17088
rect 44085 17079 44143 17085
rect 44358 17076 44364 17088
rect 44416 17076 44422 17128
rect 44542 17116 44548 17128
rect 44503 17088 44548 17116
rect 44542 17076 44548 17088
rect 44600 17076 44606 17128
rect 20717 17051 20775 17057
rect 20717 17017 20729 17051
rect 20763 17017 20775 17051
rect 20717 17011 20775 17017
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 15838 16940 15844 16992
rect 15896 16980 15902 16992
rect 15933 16983 15991 16989
rect 15933 16980 15945 16983
rect 15896 16952 15945 16980
rect 15896 16940 15902 16952
rect 15933 16949 15945 16952
rect 15979 16949 15991 16983
rect 15933 16943 15991 16949
rect 19702 16940 19708 16992
rect 19760 16980 19766 16992
rect 20530 16980 20536 16992
rect 19760 16952 20536 16980
rect 19760 16940 19766 16952
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 23566 16980 23572 16992
rect 23527 16952 23572 16980
rect 23566 16940 23572 16952
rect 23624 16940 23630 16992
rect 24213 16983 24271 16989
rect 24213 16949 24225 16983
rect 24259 16980 24271 16983
rect 24394 16980 24400 16992
rect 24259 16952 24400 16980
rect 24259 16949 24271 16952
rect 24213 16943 24271 16949
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 25222 16980 25228 16992
rect 25183 16952 25228 16980
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 26050 16980 26056 16992
rect 26011 16952 26056 16980
rect 26050 16940 26056 16952
rect 26108 16940 26114 16992
rect 30653 16983 30711 16989
rect 30653 16949 30665 16983
rect 30699 16980 30711 16983
rect 41414 16980 41420 16992
rect 30699 16952 41420 16980
rect 30699 16949 30711 16952
rect 30653 16943 30711 16949
rect 41414 16940 41420 16952
rect 41472 16980 41478 16992
rect 42242 16980 42248 16992
rect 41472 16952 42248 16980
rect 41472 16940 41478 16952
rect 42242 16940 42248 16952
rect 42300 16940 42306 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 18506 16776 18512 16788
rect 18467 16748 18512 16776
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 18616 16748 19656 16776
rect 17310 16708 17316 16720
rect 15672 16680 17316 16708
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 15672 16649 15700 16680
rect 17310 16668 17316 16680
rect 17368 16668 17374 16720
rect 17402 16668 17408 16720
rect 17460 16708 17466 16720
rect 18616 16708 18644 16748
rect 17460 16680 18644 16708
rect 19521 16711 19579 16717
rect 17460 16668 17466 16680
rect 19521 16677 19533 16711
rect 19567 16677 19579 16711
rect 19628 16708 19656 16748
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 22925 16779 22983 16785
rect 22925 16776 22937 16779
rect 22152 16748 22937 16776
rect 22152 16736 22158 16748
rect 22925 16745 22937 16748
rect 22971 16745 22983 16779
rect 44542 16776 44548 16788
rect 22925 16739 22983 16745
rect 24504 16748 44548 16776
rect 24504 16708 24532 16748
rect 44542 16736 44548 16748
rect 44600 16736 44606 16788
rect 19628 16680 24532 16708
rect 19521 16671 19579 16677
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16609 15715 16643
rect 15838 16640 15844 16652
rect 15799 16612 15844 16640
rect 15657 16603 15715 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 19536 16640 19564 16671
rect 27338 16668 27344 16720
rect 27396 16708 27402 16720
rect 27396 16680 27936 16708
rect 27396 16668 27402 16680
rect 20990 16640 20996 16652
rect 18524 16612 19564 16640
rect 19812 16612 20996 16640
rect 18524 16581 18552 16612
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18690 16572 18696 16584
rect 18651 16544 18696 16572
rect 18509 16535 18567 16541
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 19702 16572 19708 16584
rect 19663 16544 19708 16572
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19812 16581 19840 16612
rect 20990 16600 20996 16612
rect 21048 16640 21054 16652
rect 24394 16640 24400 16652
rect 21048 16612 22094 16640
rect 24355 16612 24400 16640
rect 21048 16600 21054 16612
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 20404 16544 20637 16572
rect 20404 16532 20410 16544
rect 20625 16541 20637 16544
rect 20671 16541 20683 16575
rect 22066 16572 22094 16612
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 24673 16643 24731 16649
rect 24673 16609 24685 16643
rect 24719 16640 24731 16643
rect 25406 16640 25412 16652
rect 24719 16612 25412 16640
rect 24719 16609 24731 16612
rect 24673 16603 24731 16609
rect 25406 16600 25412 16612
rect 25464 16600 25470 16652
rect 26142 16640 26148 16652
rect 26103 16612 26148 16640
rect 26142 16600 26148 16612
rect 26200 16600 26206 16652
rect 26418 16600 26424 16652
rect 26476 16640 26482 16652
rect 27908 16640 27936 16680
rect 27982 16668 27988 16720
rect 28040 16708 28046 16720
rect 28537 16711 28595 16717
rect 28537 16708 28549 16711
rect 28040 16680 28549 16708
rect 28040 16668 28046 16680
rect 28537 16677 28549 16680
rect 28583 16677 28595 16711
rect 38654 16708 38660 16720
rect 28537 16671 28595 16677
rect 31220 16680 38660 16708
rect 26476 16612 26648 16640
rect 27908 16612 28028 16640
rect 26476 16600 26482 16612
rect 23109 16575 23167 16581
rect 23109 16572 23121 16575
rect 22066 16544 23121 16572
rect 20625 16535 20683 16541
rect 23109 16541 23121 16544
rect 23155 16541 23167 16575
rect 23109 16535 23167 16541
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 23474 16572 23480 16584
rect 23431 16544 23480 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 23566 16532 23572 16584
rect 23624 16572 23630 16584
rect 26620 16581 26648 16612
rect 26605 16575 26663 16581
rect 23624 16544 23669 16572
rect 23624 16532 23630 16544
rect 26605 16541 26617 16575
rect 26651 16541 26663 16575
rect 26605 16535 26663 16541
rect 27798 16532 27804 16584
rect 27856 16572 27862 16584
rect 28000 16581 28028 16612
rect 28258 16600 28264 16652
rect 28316 16640 28322 16652
rect 28316 16612 28488 16640
rect 28316 16600 28322 16612
rect 28460 16581 28488 16612
rect 31220 16581 31248 16680
rect 38654 16668 38660 16680
rect 38712 16708 38718 16720
rect 39114 16708 39120 16720
rect 38712 16680 39120 16708
rect 38712 16668 38718 16680
rect 39114 16668 39120 16680
rect 39172 16668 39178 16720
rect 45002 16708 45008 16720
rect 44915 16680 45008 16708
rect 45002 16668 45008 16680
rect 45060 16708 45066 16720
rect 46934 16708 46940 16720
rect 45060 16680 46940 16708
rect 45060 16668 45066 16680
rect 46934 16668 46940 16680
rect 46992 16668 46998 16720
rect 42610 16640 42616 16652
rect 42571 16612 42616 16640
rect 42610 16600 42616 16612
rect 42668 16600 42674 16652
rect 45020 16581 45048 16668
rect 46293 16643 46351 16649
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47762 16640 47768 16652
rect 46339 16612 47768 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47762 16600 47768 16612
rect 47820 16600 47826 16652
rect 27985 16575 28043 16581
rect 27856 16544 27901 16572
rect 27856 16532 27862 16544
rect 27985 16541 27997 16575
rect 28031 16541 28043 16575
rect 27985 16535 28043 16541
rect 28445 16575 28503 16581
rect 28445 16541 28457 16575
rect 28491 16541 28503 16575
rect 28445 16535 28503 16541
rect 31205 16575 31263 16581
rect 31205 16541 31217 16575
rect 31251 16541 31263 16575
rect 31205 16535 31263 16541
rect 45005 16575 45063 16581
rect 45005 16541 45017 16575
rect 45051 16541 45063 16575
rect 45005 16535 45063 16541
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 17494 16504 17500 16516
rect 17455 16476 17500 16504
rect 17494 16464 17500 16476
rect 17552 16464 17558 16516
rect 19518 16504 19524 16516
rect 19479 16476 19524 16504
rect 19518 16464 19524 16476
rect 19576 16464 19582 16516
rect 20806 16504 20812 16516
rect 20767 16476 20812 16504
rect 20806 16464 20812 16476
rect 20864 16464 20870 16516
rect 22465 16507 22523 16513
rect 22465 16473 22477 16507
rect 22511 16473 22523 16507
rect 26050 16504 26056 16516
rect 25898 16476 26056 16504
rect 22465 16467 22523 16473
rect 22480 16436 22508 16467
rect 26050 16464 26056 16476
rect 26108 16464 26114 16516
rect 42797 16507 42855 16513
rect 26160 16476 31754 16504
rect 26160 16436 26188 16476
rect 26694 16436 26700 16448
rect 22480 16408 26188 16436
rect 26655 16408 26700 16436
rect 26694 16396 26700 16408
rect 26752 16396 26758 16448
rect 27985 16439 28043 16445
rect 27985 16405 27997 16439
rect 28031 16436 28043 16439
rect 28166 16436 28172 16448
rect 28031 16408 28172 16436
rect 28031 16405 28043 16408
rect 27985 16399 28043 16405
rect 28166 16396 28172 16408
rect 28224 16396 28230 16448
rect 30558 16396 30564 16448
rect 30616 16436 30622 16448
rect 31297 16439 31355 16445
rect 31297 16436 31309 16439
rect 30616 16408 31309 16436
rect 30616 16396 30622 16408
rect 31297 16405 31309 16408
rect 31343 16405 31355 16439
rect 31726 16436 31754 16476
rect 42797 16473 42809 16507
rect 42843 16504 42855 16507
rect 42886 16504 42892 16516
rect 42843 16476 42892 16504
rect 42843 16473 42855 16476
rect 42797 16467 42855 16473
rect 42886 16464 42892 16476
rect 42944 16464 42950 16516
rect 44453 16507 44511 16513
rect 44453 16473 44465 16507
rect 44499 16504 44511 16507
rect 46014 16504 46020 16516
rect 44499 16476 46020 16504
rect 44499 16473 44511 16476
rect 44453 16467 44511 16473
rect 46014 16464 46020 16476
rect 46072 16464 46078 16516
rect 46474 16504 46480 16516
rect 46435 16476 46480 16504
rect 46474 16464 46480 16476
rect 46532 16464 46538 16516
rect 48130 16504 48136 16516
rect 48091 16476 48136 16504
rect 48130 16464 48136 16476
rect 48188 16464 48194 16516
rect 43714 16436 43720 16448
rect 31726 16408 43720 16436
rect 31297 16399 31355 16405
rect 43714 16396 43720 16408
rect 43772 16396 43778 16448
rect 44082 16396 44088 16448
rect 44140 16436 44146 16448
rect 45097 16439 45155 16445
rect 45097 16436 45109 16439
rect 44140 16408 45109 16436
rect 44140 16396 44146 16408
rect 45097 16405 45109 16408
rect 45143 16405 45155 16439
rect 45097 16399 45155 16405
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 19337 16235 19395 16241
rect 12406 16204 19288 16232
rect 12406 16164 12434 16204
rect 6886 16136 12434 16164
rect 16025 16167 16083 16173
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16096 2099 16099
rect 6886 16096 6914 16136
rect 16025 16133 16037 16167
rect 16071 16164 16083 16167
rect 16853 16167 16911 16173
rect 16853 16164 16865 16167
rect 16071 16136 16865 16164
rect 16071 16133 16083 16136
rect 16025 16127 16083 16133
rect 16853 16133 16865 16136
rect 16899 16133 16911 16167
rect 19260 16164 19288 16204
rect 19337 16201 19349 16235
rect 19383 16232 19395 16235
rect 19426 16232 19432 16244
rect 19383 16204 19432 16232
rect 19383 16201 19395 16204
rect 19337 16195 19395 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 21818 16192 21824 16244
rect 21876 16232 21882 16244
rect 22005 16235 22063 16241
rect 22005 16232 22017 16235
rect 21876 16204 22017 16232
rect 21876 16192 21882 16204
rect 22005 16201 22017 16204
rect 22051 16201 22063 16235
rect 22005 16195 22063 16201
rect 25406 16192 25412 16244
rect 25464 16232 25470 16244
rect 25593 16235 25651 16241
rect 25593 16232 25605 16235
rect 25464 16204 25605 16232
rect 25464 16192 25470 16204
rect 25593 16201 25605 16204
rect 25639 16201 25651 16235
rect 25593 16195 25651 16201
rect 27157 16235 27215 16241
rect 27157 16201 27169 16235
rect 27203 16232 27215 16235
rect 28074 16232 28080 16244
rect 27203 16204 28080 16232
rect 27203 16201 27215 16204
rect 27157 16195 27215 16201
rect 28074 16192 28080 16204
rect 28132 16192 28138 16244
rect 28534 16232 28540 16244
rect 28495 16204 28540 16232
rect 28534 16192 28540 16204
rect 28592 16192 28598 16244
rect 42886 16232 42892 16244
rect 42847 16204 42892 16232
rect 42886 16192 42892 16204
rect 42944 16192 42950 16244
rect 43714 16192 43720 16244
rect 43772 16232 43778 16244
rect 45646 16232 45652 16244
rect 43772 16204 45652 16232
rect 43772 16192 43778 16204
rect 45646 16192 45652 16204
rect 45704 16192 45710 16244
rect 20898 16164 20904 16176
rect 19260 16136 20904 16164
rect 16853 16127 16911 16133
rect 20898 16124 20904 16136
rect 20956 16124 20962 16176
rect 28166 16124 28172 16176
rect 28224 16164 28230 16176
rect 44082 16164 44088 16176
rect 28224 16136 28580 16164
rect 44043 16136 44088 16164
rect 28224 16124 28230 16136
rect 15930 16096 15936 16108
rect 2087 16068 6914 16096
rect 15891 16068 15936 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 19150 16056 19156 16108
rect 19208 16096 19214 16108
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 19208 16068 19257 16096
rect 19208 16056 19214 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 19245 16059 19303 16065
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16096 25283 16099
rect 26142 16096 26148 16108
rect 25271 16068 26148 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 16666 16028 16672 16040
rect 16627 16000 16672 16028
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 17129 16031 17187 16037
rect 17129 15997 17141 16031
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 22741 16031 22799 16037
rect 22741 15997 22753 16031
rect 22787 15997 22799 16031
rect 22741 15991 22799 15997
rect 22925 16031 22983 16037
rect 22925 15997 22937 16031
rect 22971 16028 22983 16031
rect 23382 16028 23388 16040
rect 22971 16000 23388 16028
rect 22971 15997 22983 16000
rect 22925 15991 22983 15997
rect 3234 15920 3240 15972
rect 3292 15960 3298 15972
rect 3292 15932 6914 15960
rect 3292 15920 3298 15932
rect 6886 15892 6914 15932
rect 17144 15892 17172 15991
rect 22756 15960 22784 15991
rect 23382 15988 23388 16000
rect 23440 15988 23446 16040
rect 24302 16028 24308 16040
rect 24263 16000 24308 16028
rect 24302 15988 24308 16000
rect 24360 15988 24366 16040
rect 25130 16028 25136 16040
rect 25091 16000 25136 16028
rect 25130 15988 25136 16000
rect 25188 15988 25194 16040
rect 23198 15960 23204 15972
rect 22756 15932 23204 15960
rect 23198 15920 23204 15932
rect 23256 15960 23262 15972
rect 25240 15960 25268 16059
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 27062 16096 27068 16108
rect 27023 16068 27068 16096
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27249 16099 27307 16105
rect 27249 16096 27261 16099
rect 27212 16068 27261 16096
rect 27212 16056 27218 16068
rect 27249 16065 27261 16068
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 27890 16056 27896 16108
rect 27948 16096 27954 16108
rect 28552 16105 28580 16136
rect 44082 16124 44088 16136
rect 44140 16124 44146 16176
rect 28353 16099 28411 16105
rect 28353 16096 28365 16099
rect 27948 16068 28365 16096
rect 27948 16056 27954 16068
rect 28353 16065 28365 16068
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 28537 16099 28595 16105
rect 28537 16065 28549 16099
rect 28583 16065 28595 16099
rect 28537 16059 28595 16065
rect 38654 16056 38660 16108
rect 38712 16096 38718 16108
rect 42797 16099 42855 16105
rect 42797 16096 42809 16099
rect 38712 16068 42809 16096
rect 38712 16056 38718 16068
rect 42797 16065 42809 16068
rect 42843 16065 42855 16099
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 42797 16059 42855 16065
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 42242 15988 42248 16040
rect 42300 16028 42306 16040
rect 43901 16031 43959 16037
rect 43901 16028 43913 16031
rect 42300 16000 43913 16028
rect 42300 15988 42306 16000
rect 43901 15997 43913 16000
rect 43947 15997 43959 16031
rect 45094 16028 45100 16040
rect 45055 16000 45100 16028
rect 43901 15991 43959 15997
rect 45094 15988 45100 16000
rect 45152 15988 45158 16040
rect 23256 15932 25268 15960
rect 23256 15920 23262 15932
rect 6886 15864 17172 15892
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 21821 15691 21879 15697
rect 21821 15657 21833 15691
rect 21867 15688 21879 15691
rect 22554 15688 22560 15700
rect 21867 15660 22560 15688
rect 21867 15657 21879 15660
rect 21821 15651 21879 15657
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 23198 15688 23204 15700
rect 23159 15660 23204 15688
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 23290 15648 23296 15700
rect 23348 15688 23354 15700
rect 23385 15691 23443 15697
rect 23385 15688 23397 15691
rect 23348 15660 23397 15688
rect 23348 15648 23354 15660
rect 23385 15657 23397 15660
rect 23431 15657 23443 15691
rect 23385 15651 23443 15657
rect 24489 15691 24547 15697
rect 24489 15657 24501 15691
rect 24535 15688 24547 15691
rect 25130 15688 25136 15700
rect 24535 15660 25136 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 25130 15648 25136 15660
rect 25188 15648 25194 15700
rect 47486 15648 47492 15700
rect 47544 15688 47550 15700
rect 47673 15691 47731 15697
rect 47673 15688 47685 15691
rect 47544 15660 47685 15688
rect 47544 15648 47550 15660
rect 47673 15657 47685 15660
rect 47719 15657 47731 15691
rect 47673 15651 47731 15657
rect 24596 15592 25452 15620
rect 24596 15496 24624 15592
rect 25222 15512 25228 15564
rect 25280 15552 25286 15564
rect 25317 15555 25375 15561
rect 25317 15552 25329 15555
rect 25280 15524 25329 15552
rect 25280 15512 25286 15524
rect 25317 15521 25329 15524
rect 25363 15521 25375 15555
rect 25424 15552 25452 15592
rect 27065 15555 27123 15561
rect 27065 15552 27077 15555
rect 25424 15524 27077 15552
rect 25317 15515 25375 15521
rect 27065 15521 27077 15524
rect 27111 15552 27123 15555
rect 30377 15555 30435 15561
rect 30377 15552 30389 15555
rect 27111 15524 30389 15552
rect 27111 15521 27123 15524
rect 27065 15515 27123 15521
rect 30377 15521 30389 15524
rect 30423 15521 30435 15555
rect 30558 15552 30564 15564
rect 30519 15524 30564 15552
rect 30377 15515 30435 15521
rect 30558 15512 30564 15524
rect 30616 15512 30622 15564
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 21729 15487 21787 15493
rect 21729 15484 21741 15487
rect 19208 15456 21741 15484
rect 19208 15444 19214 15456
rect 21729 15453 21741 15456
rect 21775 15453 21787 15487
rect 21729 15447 21787 15453
rect 23842 15444 23848 15496
rect 23900 15484 23906 15496
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 23900 15456 24409 15484
rect 23900 15444 23906 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 24397 15447 24455 15453
rect 24578 15444 24584 15496
rect 24636 15484 24642 15496
rect 24636 15456 24729 15484
rect 24636 15444 24642 15456
rect 26694 15444 26700 15496
rect 26752 15444 26758 15496
rect 16666 15376 16672 15428
rect 16724 15416 16730 15428
rect 23017 15419 23075 15425
rect 23017 15416 23029 15419
rect 16724 15388 23029 15416
rect 16724 15376 16730 15388
rect 23017 15385 23029 15388
rect 23063 15416 23075 15419
rect 23566 15416 23572 15428
rect 23063 15388 23572 15416
rect 23063 15385 23075 15388
rect 23017 15379 23075 15385
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 25590 15416 25596 15428
rect 25551 15388 25596 15416
rect 25590 15376 25596 15388
rect 25648 15376 25654 15428
rect 32214 15416 32220 15428
rect 32175 15388 32220 15416
rect 32214 15376 32220 15388
rect 32272 15376 32278 15428
rect 23106 15308 23112 15360
rect 23164 15348 23170 15360
rect 23227 15351 23285 15357
rect 23227 15348 23239 15351
rect 23164 15320 23239 15348
rect 23164 15308 23170 15320
rect 23227 15317 23239 15320
rect 23273 15348 23285 15351
rect 24578 15348 24584 15360
rect 23273 15320 24584 15348
rect 23273 15317 23285 15320
rect 23227 15311 23285 15317
rect 24578 15308 24584 15320
rect 24636 15308 24642 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 23382 15144 23388 15156
rect 23343 15116 23388 15144
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 23014 14968 23020 15020
rect 23072 15008 23078 15020
rect 23293 15011 23351 15017
rect 23293 15008 23305 15011
rect 23072 14980 23305 15008
rect 23072 14968 23078 14980
rect 23293 14977 23305 14980
rect 23339 14977 23351 15011
rect 23293 14971 23351 14977
rect 24397 15011 24455 15017
rect 24397 14977 24409 15011
rect 24443 15008 24455 15011
rect 24578 15008 24584 15020
rect 24443 14980 24584 15008
rect 24443 14977 24455 14980
rect 24397 14971 24455 14977
rect 24578 14968 24584 14980
rect 24636 14968 24642 15020
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2314 14940 2320 14952
rect 1995 14912 2320 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 23842 14900 23848 14952
rect 23900 14940 23906 14952
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 23900 14912 24317 14940
rect 23900 14900 23906 14912
rect 24305 14909 24317 14912
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24765 14943 24823 14949
rect 24765 14909 24777 14943
rect 24811 14940 24823 14943
rect 25590 14940 25596 14952
rect 24811 14912 25596 14940
rect 24811 14909 24823 14912
rect 24765 14903 24823 14909
rect 25590 14900 25596 14912
rect 25648 14900 25654 14952
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 23014 14872 23020 14884
rect 22796 14844 23020 14872
rect 22796 14832 22802 14844
rect 23014 14832 23020 14844
rect 23072 14832 23078 14884
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2314 14600 2320 14612
rect 2275 14572 2320 14600
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2682 14396 2688 14408
rect 2271 14368 2688 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 25774 14396 25780 14408
rect 2740 14368 25780 14396
rect 2740 14356 2746 14368
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 15286 13784 15292 13796
rect 3476 13756 15292 13784
rect 3476 13744 3482 13756
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 22005 13379 22063 13385
rect 22005 13345 22017 13379
rect 22051 13376 22063 13379
rect 22830 13376 22836 13388
rect 22051 13348 22836 13376
rect 22051 13345 22063 13348
rect 22005 13339 22063 13345
rect 22830 13336 22836 13348
rect 22888 13336 22894 13388
rect 23658 13376 23664 13388
rect 23619 13348 23664 13376
rect 23658 13336 23664 13348
rect 23716 13336 23722 13388
rect 47670 13308 47676 13320
rect 47631 13280 47676 13308
rect 47670 13268 47676 13280
rect 47728 13268 47734 13320
rect 22189 13243 22247 13249
rect 22189 13209 22201 13243
rect 22235 13240 22247 13243
rect 22462 13240 22468 13252
rect 22235 13212 22468 13240
rect 22235 13209 22247 13212
rect 22189 13203 22247 13209
rect 22462 13200 22468 13212
rect 22520 13200 22526 13252
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 22462 12968 22468 12980
rect 22423 12940 22468 12968
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 22370 12832 22376 12844
rect 22283 12804 22376 12832
rect 22370 12792 22376 12804
rect 22428 12832 22434 12844
rect 47302 12832 47308 12844
rect 22428 12804 47308 12832
rect 22428 12792 22434 12804
rect 47302 12792 47308 12804
rect 47360 12792 47366 12844
rect 30006 12696 30012 12708
rect 6886 12668 30012 12696
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 6886 12628 6914 12668
rect 30006 12656 30012 12668
rect 30064 12656 30070 12708
rect 47762 12628 47768 12640
rect 1627 12600 6914 12628
rect 47723 12600 47768 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 47762 12588 47768 12600
rect 47820 12588 47826 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 46293 12291 46351 12297
rect 46293 12257 46305 12291
rect 46339 12288 46351 12291
rect 47670 12288 47676 12300
rect 46339 12260 47676 12288
rect 46339 12257 46351 12260
rect 46293 12251 46351 12257
rect 47670 12248 47676 12260
rect 47728 12248 47734 12300
rect 48130 12288 48136 12300
rect 48091 12260 48136 12288
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 46477 12155 46535 12161
rect 46477 12121 46489 12155
rect 46523 12152 46535 12155
rect 47670 12152 47676 12164
rect 46523 12124 47676 12152
rect 46523 12121 46535 12124
rect 46477 12115 46535 12121
rect 47670 12112 47676 12124
rect 47728 12112 47734 12164
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 47670 11880 47676 11892
rect 47631 11852 47676 11880
rect 47670 11840 47676 11852
rect 47728 11840 47734 11892
rect 41506 11704 41512 11756
rect 41564 11744 41570 11756
rect 46661 11747 46719 11753
rect 46661 11744 46673 11747
rect 41564 11716 46673 11744
rect 41564 11704 41570 11716
rect 46661 11713 46673 11716
rect 46707 11713 46719 11747
rect 46661 11707 46719 11713
rect 46934 11704 46940 11756
rect 46992 11744 46998 11756
rect 47581 11747 47639 11753
rect 47581 11744 47593 11747
rect 46992 11716 47593 11744
rect 46992 11704 46998 11716
rect 47581 11713 47593 11716
rect 47627 11713 47639 11747
rect 47581 11707 47639 11713
rect 46474 11500 46480 11552
rect 46532 11540 46538 11552
rect 46753 11543 46811 11549
rect 46753 11540 46765 11543
rect 46532 11512 46765 11540
rect 46532 11500 46538 11512
rect 46753 11509 46765 11512
rect 46799 11509 46811 11543
rect 46753 11503 46811 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 47762 11268 47768 11280
rect 46308 11240 47768 11268
rect 46308 11209 46336 11240
rect 47762 11228 47768 11240
rect 47820 11228 47826 11280
rect 46293 11203 46351 11209
rect 46293 11169 46305 11203
rect 46339 11169 46351 11203
rect 46474 11200 46480 11212
rect 46435 11172 46480 11200
rect 46293 11163 46351 11169
rect 46474 11160 46480 11172
rect 46532 11160 46538 11212
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 12434 10996 12440 11008
rect 4120 10968 12440 10996
rect 4120 10956 4126 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 47486 10616 47492 10668
rect 47544 10656 47550 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 47544 10628 47593 10656
rect 47544 10616 47550 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 47029 10455 47087 10461
rect 47029 10452 47041 10455
rect 46348 10424 47041 10452
rect 46348 10412 46354 10424
rect 47029 10421 47041 10424
rect 47075 10421 47087 10455
rect 47670 10452 47676 10464
rect 47631 10424 47676 10452
rect 47029 10415 47087 10421
rect 47670 10412 47676 10424
rect 47728 10412 47734 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 46477 10115 46535 10121
rect 46477 10081 46489 10115
rect 46523 10112 46535 10115
rect 47670 10112 47676 10124
rect 46523 10084 47676 10112
rect 46523 10081 46535 10084
rect 46477 10075 46535 10081
rect 47670 10072 47676 10084
rect 47728 10072 47734 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 47854 9568 47860 9580
rect 47815 9540 47860 9568
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 48041 9435 48099 9441
rect 48041 9401 48053 9435
rect 48087 9432 48099 9435
rect 48222 9432 48228 9444
rect 48087 9404 48228 9432
rect 48087 9401 48099 9404
rect 48041 9395 48099 9401
rect 48222 9392 48228 9404
rect 48280 9392 48286 9444
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47762 8888 47768 8900
rect 47723 8860 47768 8888
rect 47762 8848 47768 8860
rect 47820 8848 47826 8900
rect 27522 8780 27528 8832
rect 27580 8820 27586 8832
rect 47857 8823 47915 8829
rect 47857 8820 47869 8823
rect 27580 8792 47869 8820
rect 27580 8780 27586 8792
rect 47857 8789 47869 8792
rect 47903 8789 47915 8823
rect 47857 8783 47915 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 48130 8480 48136 8492
rect 48091 8452 48136 8480
rect 48130 8440 48136 8452
rect 48188 8440 48194 8492
rect 47118 8236 47124 8288
rect 47176 8276 47182 8288
rect 47949 8279 48007 8285
rect 47949 8276 47961 8279
rect 47176 8248 47961 8276
rect 47176 8236 47182 8248
rect 47949 8245 47961 8248
rect 47995 8245 48007 8279
rect 47949 8239 48007 8245
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 46768 7976 47440 8004
rect 46768 7948 46796 7976
rect 45554 7936 45560 7948
rect 45515 7908 45560 7936
rect 45554 7896 45560 7908
rect 45612 7896 45618 7948
rect 46569 7939 46627 7945
rect 46569 7905 46581 7939
rect 46615 7936 46627 7939
rect 46750 7936 46756 7948
rect 46615 7908 46756 7936
rect 46615 7905 46627 7908
rect 46569 7899 46627 7905
rect 46750 7896 46756 7908
rect 46808 7896 46814 7948
rect 47118 7936 47124 7948
rect 47079 7908 47124 7936
rect 47118 7896 47124 7908
rect 47176 7896 47182 7948
rect 47412 7945 47440 7976
rect 47397 7939 47455 7945
rect 47397 7905 47409 7939
rect 47443 7905 47455 7939
rect 47397 7899 47455 7905
rect 45649 7803 45707 7809
rect 45649 7769 45661 7803
rect 45695 7800 45707 7803
rect 47213 7803 47271 7809
rect 45695 7772 46336 7800
rect 45695 7769 45707 7772
rect 45649 7763 45707 7769
rect 46308 7744 46336 7772
rect 47213 7769 47225 7803
rect 47259 7800 47271 7803
rect 47578 7800 47584 7812
rect 47259 7772 47584 7800
rect 47259 7769 47271 7772
rect 47213 7763 47271 7769
rect 47578 7760 47584 7772
rect 47636 7760 47642 7812
rect 46290 7692 46296 7744
rect 46348 7692 46354 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 47578 7528 47584 7540
rect 47539 7500 47584 7528
rect 47578 7488 47584 7500
rect 47636 7488 47642 7540
rect 46290 7392 46296 7404
rect 46251 7364 46296 7392
rect 46290 7352 46296 7364
rect 46348 7352 46354 7404
rect 47765 7395 47823 7401
rect 47765 7392 47777 7395
rect 46768 7364 47777 7392
rect 46768 7333 46796 7364
rect 47765 7361 47777 7364
rect 47811 7361 47823 7395
rect 47765 7355 47823 7361
rect 46753 7327 46811 7333
rect 46753 7293 46765 7327
rect 46799 7293 46811 7327
rect 46753 7287 46811 7293
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 45925 7259 45983 7265
rect 45925 7256 45937 7259
rect 2096 7228 45937 7256
rect 2096 7216 2102 7228
rect 45925 7225 45937 7228
rect 45971 7256 45983 7259
rect 45971 7228 46428 7256
rect 45971 7225 45983 7228
rect 45925 7219 45983 7225
rect 46400 7197 46428 7228
rect 46385 7191 46443 7197
rect 46385 7157 46397 7191
rect 46431 7157 46443 7191
rect 46385 7151 46443 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 17494 6848 17500 6860
rect 4120 6820 17500 6848
rect 4120 6808 4126 6820
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 41785 6851 41843 6857
rect 41785 6817 41797 6851
rect 41831 6848 41843 6851
rect 43530 6848 43536 6860
rect 41831 6820 43536 6848
rect 41831 6817 41843 6820
rect 41785 6811 41843 6817
rect 43530 6808 43536 6820
rect 43588 6808 43594 6860
rect 47302 6848 47308 6860
rect 47263 6820 47308 6848
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 47394 6808 47400 6860
rect 47452 6848 47458 6860
rect 47581 6851 47639 6857
rect 47581 6848 47593 6851
rect 47452 6820 47593 6848
rect 47452 6808 47458 6820
rect 47581 6817 47593 6820
rect 47627 6817 47639 6851
rect 47581 6811 47639 6817
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 40313 6715 40371 6721
rect 40313 6712 40325 6715
rect 4028 6684 40325 6712
rect 4028 6672 4034 6684
rect 40313 6681 40325 6684
rect 40359 6712 40371 6715
rect 40773 6715 40831 6721
rect 40773 6712 40785 6715
rect 40359 6684 40785 6712
rect 40359 6681 40371 6684
rect 40313 6675 40371 6681
rect 40773 6681 40785 6684
rect 40819 6681 40831 6715
rect 40773 6675 40831 6681
rect 40862 6672 40868 6724
rect 40920 6712 40926 6724
rect 40920 6684 40965 6712
rect 40920 6672 40926 6684
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 40681 6443 40739 6449
rect 40681 6409 40693 6443
rect 40727 6440 40739 6443
rect 40862 6440 40868 6452
rect 40727 6412 40868 6440
rect 40727 6409 40739 6412
rect 40681 6403 40739 6409
rect 40862 6400 40868 6412
rect 40920 6400 40926 6452
rect 44634 6400 44640 6452
rect 44692 6440 44698 6452
rect 48041 6443 48099 6449
rect 48041 6440 48053 6443
rect 44692 6412 48053 6440
rect 44692 6400 44698 6412
rect 48041 6409 48053 6412
rect 48087 6409 48099 6443
rect 48041 6403 48099 6409
rect 40862 6304 40868 6316
rect 40823 6276 40868 6304
rect 40862 6264 40868 6276
rect 40920 6264 40926 6316
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 45554 5828 45560 5840
rect 41892 5800 45560 5828
rect 41892 5772 41920 5800
rect 45554 5788 45560 5800
rect 45612 5788 45618 5840
rect 41874 5760 41880 5772
rect 41787 5732 41880 5760
rect 41874 5720 41880 5732
rect 41932 5720 41938 5772
rect 42705 5763 42763 5769
rect 42705 5729 42717 5763
rect 42751 5760 42763 5763
rect 43530 5760 43536 5772
rect 42751 5732 43536 5760
rect 42751 5729 42763 5732
rect 42705 5723 42763 5729
rect 43530 5720 43536 5732
rect 43588 5720 43594 5772
rect 41966 5584 41972 5636
rect 42024 5624 42030 5636
rect 42024 5596 42069 5624
rect 42024 5584 42030 5596
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 40681 5355 40739 5361
rect 40681 5321 40693 5355
rect 40727 5352 40739 5355
rect 40862 5352 40868 5364
rect 40727 5324 40868 5352
rect 40727 5321 40739 5324
rect 40681 5315 40739 5321
rect 40862 5312 40868 5324
rect 40920 5312 40926 5364
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5216 21879 5219
rect 22094 5216 22100 5228
rect 21867 5188 22100 5216
rect 21867 5185 21879 5188
rect 21821 5179 21879 5185
rect 22094 5176 22100 5188
rect 22152 5176 22158 5228
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5216 22523 5219
rect 23842 5216 23848 5228
rect 22511 5188 23848 5216
rect 22511 5185 22523 5188
rect 22465 5179 22523 5185
rect 23842 5176 23848 5188
rect 23900 5176 23906 5228
rect 40221 5219 40279 5225
rect 40221 5185 40233 5219
rect 40267 5216 40279 5219
rect 41966 5216 41972 5228
rect 40267 5188 41972 5216
rect 40267 5185 40279 5188
rect 40221 5179 40279 5185
rect 41966 5176 41972 5188
rect 42024 5176 42030 5228
rect 47762 5216 47768 5228
rect 47723 5188 47768 5216
rect 47762 5176 47768 5188
rect 47820 5176 47826 5228
rect 19058 5108 19064 5160
rect 19116 5148 19122 5160
rect 32030 5148 32036 5160
rect 19116 5120 32036 5148
rect 19116 5108 19122 5120
rect 32030 5108 32036 5120
rect 32088 5108 32094 5160
rect 21913 5083 21971 5089
rect 21913 5049 21925 5083
rect 21959 5080 21971 5083
rect 23106 5080 23112 5092
rect 21959 5052 23112 5080
rect 21959 5049 21971 5052
rect 21913 5043 21971 5049
rect 23106 5040 23112 5052
rect 23164 5040 23170 5092
rect 47949 5083 48007 5089
rect 47949 5080 47961 5083
rect 31726 5052 47961 5080
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 22557 5015 22615 5021
rect 22557 5012 22569 5015
rect 22336 4984 22569 5012
rect 22336 4972 22342 4984
rect 22557 4981 22569 4984
rect 22603 4981 22615 5015
rect 22557 4975 22615 4981
rect 22922 4972 22928 5024
rect 22980 5012 22986 5024
rect 31726 5012 31754 5052
rect 47949 5049 47961 5052
rect 47995 5049 48007 5083
rect 47949 5043 48007 5049
rect 40310 5012 40316 5024
rect 22980 4984 31754 5012
rect 40271 4984 40316 5012
rect 22980 4972 22986 4984
rect 40310 4972 40316 4984
rect 40368 4972 40374 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 32306 4808 32312 4820
rect 19392 4780 32312 4808
rect 19392 4768 19398 4780
rect 32306 4768 32312 4780
rect 32364 4768 32370 4820
rect 22370 4740 22376 4752
rect 12406 4712 22376 4740
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 12406 4604 12434 4712
rect 22370 4700 22376 4712
rect 22428 4700 22434 4752
rect 31754 4700 31760 4752
rect 31812 4740 31818 4752
rect 40310 4740 40316 4752
rect 31812 4712 40316 4740
rect 31812 4700 31818 4712
rect 40310 4700 40316 4712
rect 40368 4700 40374 4752
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 22741 4675 22799 4681
rect 22152 4644 22197 4672
rect 22152 4632 22158 4644
rect 22741 4641 22753 4675
rect 22787 4672 22799 4675
rect 23750 4672 23756 4684
rect 22787 4644 23756 4672
rect 22787 4641 22799 4644
rect 22741 4635 22799 4641
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 37921 4675 37979 4681
rect 37921 4641 37933 4675
rect 37967 4672 37979 4675
rect 38562 4672 38568 4684
rect 37967 4644 38568 4672
rect 37967 4641 37979 4644
rect 37921 4635 37979 4641
rect 38562 4632 38568 4644
rect 38620 4632 38626 4684
rect 46290 4632 46296 4684
rect 46348 4672 46354 4684
rect 47581 4675 47639 4681
rect 47581 4672 47593 4675
rect 46348 4644 47593 4672
rect 46348 4632 46354 4644
rect 47581 4641 47593 4644
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 7423 4576 12434 4604
rect 20717 4607 20775 4613
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 20717 4573 20729 4607
rect 20763 4604 20775 4607
rect 21082 4604 21088 4616
rect 20763 4576 21088 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 21358 4604 21364 4616
rect 21319 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 22370 4604 22376 4616
rect 22051 4576 22376 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 22646 4604 22652 4616
rect 22607 4576 22652 4604
rect 22646 4564 22652 4576
rect 22704 4564 22710 4616
rect 23474 4604 23480 4616
rect 23435 4576 23480 4604
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 39945 4607 40003 4613
rect 39945 4573 39957 4607
rect 39991 4604 40003 4607
rect 40494 4604 40500 4616
rect 39991 4576 40500 4604
rect 39991 4573 40003 4576
rect 39945 4567 40003 4573
rect 40494 4564 40500 4576
rect 40552 4564 40558 4616
rect 40589 4607 40647 4613
rect 40589 4573 40601 4607
rect 40635 4573 40647 4607
rect 40589 4567 40647 4573
rect 46661 4607 46719 4613
rect 46661 4573 46673 4607
rect 46707 4573 46719 4607
rect 46661 4567 46719 4573
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 36541 4539 36599 4545
rect 36541 4536 36553 4539
rect 6696 4508 36553 4536
rect 6696 4496 6702 4508
rect 36541 4505 36553 4508
rect 36587 4536 36599 4539
rect 36909 4539 36967 4545
rect 36909 4536 36921 4539
rect 36587 4508 36921 4536
rect 36587 4505 36599 4508
rect 36541 4499 36599 4505
rect 36909 4505 36921 4508
rect 36955 4505 36967 4539
rect 36909 4499 36967 4505
rect 36998 4496 37004 4548
rect 37056 4536 37062 4548
rect 37056 4508 37101 4536
rect 37056 4496 37062 4508
rect 38654 4496 38660 4548
rect 38712 4536 38718 4548
rect 40604 4536 40632 4567
rect 38712 4508 40632 4536
rect 46676 4536 46704 4567
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47305 4607 47363 4613
rect 47305 4604 47317 4607
rect 46900 4576 47317 4604
rect 46900 4564 46906 4576
rect 47305 4573 47317 4576
rect 47351 4573 47363 4607
rect 47305 4567 47363 4573
rect 47486 4536 47492 4548
rect 46676 4508 47492 4536
rect 38712 4496 38718 4508
rect 47486 4496 47492 4508
rect 47544 4496 47550 4548
rect 7466 4468 7472 4480
rect 7427 4440 7472 4468
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 20806 4468 20812 4480
rect 20767 4440 20812 4468
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 21453 4471 21511 4477
rect 21453 4437 21465 4471
rect 21499 4468 21511 4471
rect 22462 4468 22468 4480
rect 21499 4440 22468 4468
rect 21499 4437 21511 4440
rect 21453 4431 21511 4437
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 23293 4471 23351 4477
rect 23293 4437 23305 4471
rect 23339 4468 23351 4471
rect 25314 4468 25320 4480
rect 23339 4440 25320 4468
rect 23339 4437 23351 4440
rect 23293 4431 23351 4437
rect 25314 4428 25320 4440
rect 25372 4428 25378 4480
rect 40034 4468 40040 4480
rect 39995 4440 40040 4468
rect 40034 4428 40040 4440
rect 40092 4428 40098 4480
rect 40126 4428 40132 4480
rect 40184 4468 40190 4480
rect 40681 4471 40739 4477
rect 40681 4468 40693 4471
rect 40184 4440 40693 4468
rect 40184 4428 40190 4440
rect 40681 4437 40693 4440
rect 40727 4437 40739 4471
rect 46750 4468 46756 4480
rect 46711 4440 46756 4468
rect 40681 4431 40739 4437
rect 46750 4428 46756 4440
rect 46808 4428 46814 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 20898 4264 20904 4276
rect 19260 4236 20904 4264
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4128 12127 4131
rect 13446 4128 13452 4140
rect 12115 4100 13452 4128
rect 12115 4097 12127 4100
rect 12069 4091 12127 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13596 4100 13737 4128
rect 13596 4088 13602 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 17218 4128 17224 4140
rect 16715 4100 17224 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17644 4100 17693 4128
rect 17644 4088 17650 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 18322 4128 18328 4140
rect 18283 4100 18328 4128
rect 17681 4091 17739 4097
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4060 6975 4063
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 6963 4032 7389 4060
rect 6963 4029 6975 4032
rect 6917 4023 6975 4029
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 7561 4063 7619 4069
rect 7561 4029 7573 4063
rect 7607 4060 7619 4063
rect 8294 4060 8300 4072
rect 7607 4032 8300 4060
rect 7607 4029 7619 4032
rect 7561 4023 7619 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1636 3896 2145 3924
rect 1636 3884 1642 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2832 3896 2881 3924
rect 2832 3884 2838 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 2869 3887 2927 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 8404 3924 8432 4023
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 17310 4060 17316 4072
rect 9180 4032 17316 4060
rect 9180 4020 9186 4032
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 19260 4060 19288 4236
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 21913 4267 21971 4273
rect 21913 4264 21925 4267
rect 21416 4236 21925 4264
rect 21416 4224 21422 4236
rect 21913 4233 21925 4236
rect 21959 4233 21971 4267
rect 21913 4227 21971 4233
rect 22646 4224 22652 4276
rect 22704 4264 22710 4276
rect 23201 4267 23259 4273
rect 23201 4264 23213 4267
rect 22704 4236 23213 4264
rect 22704 4224 22710 4236
rect 23201 4233 23213 4236
rect 23247 4233 23259 4267
rect 25682 4264 25688 4276
rect 23201 4227 23259 4233
rect 25240 4236 25688 4264
rect 20162 4156 20168 4208
rect 20220 4156 20226 4208
rect 22296 4168 22600 4196
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19392 4100 19441 4128
rect 19392 4088 19398 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 20070 4128 20076 4140
rect 20031 4100 20076 4128
rect 19429 4091 19487 4097
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20180 4128 20208 4156
rect 20346 4128 20352 4140
rect 20180 4100 20352 4128
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20717 4131 20775 4137
rect 20717 4097 20729 4131
rect 20763 4097 20775 4131
rect 20717 4091 20775 4097
rect 17420 4032 19288 4060
rect 19521 4063 19579 4069
rect 17420 3992 17448 4032
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 20162 4060 20168 4072
rect 19567 4032 20168 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 20732 4060 20760 4091
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 20864 4100 21833 4128
rect 20864 4088 20870 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22296 4128 22324 4168
rect 22462 4128 22468 4140
rect 22152 4100 22324 4128
rect 22423 4100 22468 4128
rect 22152 4088 22158 4100
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 22572 4128 22600 4168
rect 22738 4156 22744 4208
rect 22796 4196 22802 4208
rect 22796 4168 23244 4196
rect 22796 4156 22802 4168
rect 23216 4140 23244 4168
rect 23106 4128 23112 4140
rect 22572 4100 22692 4128
rect 23067 4100 23112 4128
rect 21266 4060 21272 4072
rect 20732 4032 21272 4060
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 21358 4020 21364 4072
rect 21416 4060 21422 4072
rect 21416 4032 22324 4060
rect 21416 4020 21422 4032
rect 10428 3964 17448 3992
rect 17773 3995 17831 4001
rect 7156 3896 8432 3924
rect 7156 3884 7162 3896
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9272 3896 9873 3924
rect 9272 3884 9278 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10428 3924 10456 3964
rect 17773 3961 17785 3995
rect 17819 3992 17831 3995
rect 18230 3992 18236 4004
rect 17819 3964 18236 3992
rect 17819 3961 17831 3964
rect 17773 3955 17831 3961
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 18782 3952 18788 4004
rect 18840 3992 18846 4004
rect 22002 3992 22008 4004
rect 18840 3964 22008 3992
rect 18840 3952 18846 3964
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 22296 3992 22324 4032
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 22557 4063 22615 4069
rect 22557 4060 22569 4063
rect 22428 4032 22569 4060
rect 22428 4020 22434 4032
rect 22557 4029 22569 4032
rect 22603 4029 22615 4063
rect 22664 4060 22692 4100
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23198 4088 23204 4140
rect 23256 4088 23262 4140
rect 23750 4128 23756 4140
rect 23711 4100 23756 4128
rect 23750 4088 23756 4100
rect 23808 4088 23814 4140
rect 23842 4088 23848 4140
rect 23900 4128 23906 4140
rect 24581 4131 24639 4137
rect 23900 4100 23945 4128
rect 23900 4088 23906 4100
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 24854 4128 24860 4140
rect 24627 4100 24860 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 24854 4088 24860 4100
rect 24912 4128 24918 4140
rect 25240 4128 25268 4236
rect 25682 4224 25688 4236
rect 25740 4224 25746 4276
rect 36541 4267 36599 4273
rect 36541 4233 36553 4267
rect 36587 4264 36599 4267
rect 36998 4264 37004 4276
rect 36587 4236 37004 4264
rect 36587 4233 36599 4236
rect 36541 4227 36599 4233
rect 36998 4224 37004 4236
rect 37056 4224 37062 4276
rect 39316 4236 41460 4264
rect 25501 4199 25559 4205
rect 25501 4165 25513 4199
rect 25547 4196 25559 4199
rect 25590 4196 25596 4208
rect 25547 4168 25596 4196
rect 25547 4165 25559 4168
rect 25501 4159 25559 4165
rect 25590 4156 25596 4168
rect 25648 4156 25654 4208
rect 37642 4196 37648 4208
rect 37603 4168 37648 4196
rect 37642 4156 37648 4168
rect 37700 4156 37706 4208
rect 38562 4196 38568 4208
rect 38523 4168 38568 4196
rect 38562 4156 38568 4168
rect 38620 4156 38626 4208
rect 36722 4128 36728 4140
rect 24912 4100 25268 4128
rect 26344 4100 31754 4128
rect 36683 4100 36728 4128
rect 24912 4088 24918 4100
rect 25222 4060 25228 4072
rect 22664 4032 25228 4060
rect 22557 4023 22615 4029
rect 25222 4020 25228 4032
rect 25280 4020 25286 4072
rect 25406 4060 25412 4072
rect 25319 4032 25412 4060
rect 25406 4020 25412 4032
rect 25464 4060 25470 4072
rect 26344 4060 26372 4100
rect 25464 4032 26372 4060
rect 26421 4063 26479 4069
rect 25464 4020 25470 4032
rect 26421 4029 26433 4063
rect 26467 4060 26479 4063
rect 27798 4060 27804 4072
rect 26467 4032 27804 4060
rect 26467 4029 26479 4032
rect 26421 4023 26479 4029
rect 27798 4020 27804 4032
rect 27856 4020 27862 4072
rect 31726 4060 31754 4100
rect 36722 4088 36728 4100
rect 36780 4088 36786 4140
rect 37550 4060 37556 4072
rect 31726 4032 37556 4060
rect 37550 4020 37556 4032
rect 37608 4020 37614 4072
rect 39316 4060 39344 4236
rect 40034 4156 40040 4208
rect 40092 4156 40098 4208
rect 39393 4131 39451 4137
rect 39393 4097 39405 4131
rect 39439 4128 39451 4131
rect 40052 4128 40080 4156
rect 39439 4100 40080 4128
rect 39439 4097 39451 4100
rect 39393 4091 39451 4097
rect 40034 4060 40040 4072
rect 38304 4032 39344 4060
rect 39995 4032 40040 4060
rect 22296 3964 24808 3992
rect 10008 3896 10456 3924
rect 10008 3884 10014 3896
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11756 3896 12173 3924
rect 11756 3884 11762 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 13998 3924 14004 3936
rect 13863 3896 14004 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 16761 3927 16819 3933
rect 16761 3893 16773 3927
rect 16807 3924 16819 3927
rect 17678 3924 17684 3936
rect 16807 3896 17684 3924
rect 16807 3893 16819 3896
rect 16761 3887 16819 3893
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 17920 3896 18429 3924
rect 17920 3884 17926 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18417 3887 18475 3893
rect 20165 3927 20223 3933
rect 20165 3893 20177 3927
rect 20211 3924 20223 3927
rect 20714 3924 20720 3936
rect 20211 3896 20720 3924
rect 20211 3893 20223 3896
rect 20165 3887 20223 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 20809 3927 20867 3933
rect 20809 3893 20821 3927
rect 20855 3924 20867 3927
rect 21818 3924 21824 3936
rect 20855 3896 21824 3924
rect 20855 3893 20867 3896
rect 20809 3887 20867 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 24302 3924 24308 3936
rect 21968 3896 24308 3924
rect 21968 3884 21974 3896
rect 24302 3884 24308 3896
rect 24360 3884 24366 3936
rect 24670 3924 24676 3936
rect 24631 3896 24676 3924
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 24780 3924 24808 3964
rect 25498 3952 25504 4004
rect 25556 3992 25562 4004
rect 38304 3992 38332 4032
rect 40034 4020 40040 4032
rect 40092 4020 40098 4072
rect 40221 4063 40279 4069
rect 40221 4029 40233 4063
rect 40267 4060 40279 4063
rect 40310 4060 40316 4072
rect 40267 4032 40316 4060
rect 40267 4029 40279 4032
rect 40221 4023 40279 4029
rect 40310 4020 40316 4032
rect 40368 4020 40374 4072
rect 40494 4060 40500 4072
rect 40455 4032 40500 4060
rect 40494 4020 40500 4032
rect 40552 4020 40558 4072
rect 41432 4060 41460 4236
rect 46382 4156 46388 4208
rect 46440 4196 46446 4208
rect 46569 4199 46627 4205
rect 46569 4196 46581 4199
rect 46440 4168 46581 4196
rect 46440 4156 46446 4168
rect 46569 4165 46581 4168
rect 46615 4165 46627 4199
rect 46569 4159 46627 4165
rect 46658 4156 46664 4208
rect 46716 4196 46722 4208
rect 47765 4199 47823 4205
rect 47765 4196 47777 4199
rect 46716 4168 47777 4196
rect 46716 4156 46722 4168
rect 47765 4165 47777 4168
rect 47811 4165 47823 4199
rect 47765 4159 47823 4165
rect 42981 4131 43039 4137
rect 42981 4097 42993 4131
rect 43027 4128 43039 4131
rect 44910 4128 44916 4140
rect 43027 4100 44916 4128
rect 43027 4097 43039 4100
rect 42981 4091 43039 4097
rect 44910 4088 44916 4100
rect 44968 4088 44974 4140
rect 48041 4063 48099 4069
rect 48041 4060 48053 4063
rect 41432 4032 48053 4060
rect 48041 4029 48053 4032
rect 48087 4029 48099 4063
rect 48041 4023 48099 4029
rect 39574 3992 39580 4004
rect 25556 3964 38332 3992
rect 38396 3964 39580 3992
rect 25556 3952 25562 3964
rect 27430 3924 27436 3936
rect 24780 3896 27436 3924
rect 27430 3884 27436 3896
rect 27488 3884 27494 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 38396 3924 38424 3964
rect 39574 3952 39580 3964
rect 39632 3952 39638 4004
rect 39758 3952 39764 4004
rect 39816 3992 39822 4004
rect 46753 3995 46811 4001
rect 46753 3992 46765 3995
rect 39816 3964 40540 3992
rect 39816 3952 39822 3964
rect 27764 3896 38424 3924
rect 27764 3884 27770 3896
rect 38470 3884 38476 3936
rect 38528 3924 38534 3936
rect 39485 3927 39543 3933
rect 39485 3924 39497 3927
rect 38528 3896 39497 3924
rect 38528 3884 38534 3896
rect 39485 3893 39497 3896
rect 39531 3893 39543 3927
rect 40512 3924 40540 3964
rect 41386 3964 46765 3992
rect 41386 3924 41414 3964
rect 46753 3961 46765 3964
rect 46799 3961 46811 3995
rect 46753 3955 46811 3961
rect 40512 3896 41414 3924
rect 39485 3887 39543 3893
rect 42794 3884 42800 3936
rect 42852 3924 42858 3936
rect 43073 3927 43131 3933
rect 43073 3924 43085 3927
rect 42852 3896 43085 3924
rect 42852 3884 42858 3896
rect 43073 3893 43085 3896
rect 43119 3893 43131 3927
rect 43806 3924 43812 3936
rect 43767 3896 43812 3924
rect 43073 3887 43131 3893
rect 43806 3884 43812 3896
rect 43864 3884 43870 3936
rect 46017 3927 46075 3933
rect 46017 3893 46029 3927
rect 46063 3924 46075 3927
rect 46290 3924 46296 3936
rect 46063 3896 46296 3924
rect 46063 3893 46075 3896
rect 46017 3887 46075 3893
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 8294 3720 8300 3732
rect 8255 3692 8300 3720
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 17218 3720 17224 3732
rect 17179 3692 17224 3720
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 22738 3720 22744 3732
rect 17368 3692 22744 3720
rect 17368 3680 17374 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 22848 3692 23152 3720
rect 22848 3652 22876 3692
rect 7576 3624 22876 3652
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 1912 3556 3985 3584
rect 1912 3544 1918 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 3973 3547 4031 3553
rect 2682 3516 2688 3528
rect 2643 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7282 3516 7288 3528
rect 7147 3488 7288 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7576 3525 7604 3624
rect 22922 3612 22928 3664
rect 22980 3652 22986 3664
rect 23017 3655 23075 3661
rect 23017 3652 23029 3655
rect 22980 3624 23029 3652
rect 22980 3612 22986 3624
rect 23017 3621 23029 3624
rect 23063 3621 23075 3655
rect 23124 3652 23152 3692
rect 23198 3680 23204 3732
rect 23256 3720 23262 3732
rect 24949 3723 25007 3729
rect 24949 3720 24961 3723
rect 23256 3692 24961 3720
rect 23256 3680 23262 3692
rect 24949 3689 24961 3692
rect 24995 3689 25007 3723
rect 32858 3720 32864 3732
rect 24949 3683 25007 3689
rect 25056 3692 32864 3720
rect 24854 3652 24860 3664
rect 23124 3624 24860 3652
rect 23017 3615 23075 3621
rect 24854 3612 24860 3624
rect 24912 3612 24918 3664
rect 9214 3584 9220 3596
rect 9175 3556 9220 3584
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9456 3556 9689 3584
rect 9456 3544 9462 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 12400 3556 14933 3584
rect 12400 3544 12406 3556
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 14921 3547 14979 3553
rect 15381 3587 15439 3593
rect 15381 3553 15393 3587
rect 15427 3584 15439 3587
rect 15427 3556 15884 3584
rect 15427 3553 15439 3556
rect 15381 3547 15439 3553
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 9122 3516 9128 3528
rect 8251 3488 9128 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11572 3488 11713 3516
rect 11572 3476 11578 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 15856 3525 15884 3556
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 20990 3584 20996 3596
rect 16448 3556 20996 3584
rect 16448 3544 16454 3556
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 21082 3544 21088 3596
rect 21140 3584 21146 3596
rect 21913 3587 21971 3593
rect 21913 3584 21925 3587
rect 21140 3556 21925 3584
rect 21140 3544 21146 3556
rect 21913 3553 21925 3556
rect 21959 3553 21971 3587
rect 21913 3547 21971 3553
rect 22002 3544 22008 3596
rect 22060 3584 22066 3596
rect 25056 3584 25084 3692
rect 32858 3680 32864 3692
rect 32916 3720 32922 3732
rect 38565 3723 38623 3729
rect 32916 3692 35894 3720
rect 32916 3680 32922 3692
rect 22060 3556 25084 3584
rect 25148 3624 29868 3652
rect 22060 3544 22066 3556
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13872 3488 14289 3516
rect 13872 3476 13878 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 15013 3519 15071 3525
rect 15013 3485 15025 3519
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 15979 3488 16497 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16485 3485 16497 3488
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1360 3420 1869 3448
rect 1360 3408 1366 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 1857 3411 1915 3417
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 9401 3451 9459 3457
rect 2271 3420 7788 3448
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2777 3383 2835 3389
rect 2777 3380 2789 3383
rect 2096 3352 2789 3380
rect 2096 3340 2102 3352
rect 2777 3349 2789 3352
rect 2823 3349 2835 3383
rect 2777 3343 2835 3349
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7653 3383 7711 3389
rect 7653 3380 7665 3383
rect 6972 3352 7665 3380
rect 6972 3340 6978 3352
rect 7653 3349 7665 3352
rect 7699 3349 7711 3383
rect 7760 3380 7788 3420
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 10134 3448 10140 3460
rect 9447 3420 10140 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 15028 3448 15056 3479
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 16816 3488 17141 3516
rect 16816 3476 16822 3488
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 17678 3476 17684 3528
rect 17736 3516 17742 3528
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17736 3488 17785 3516
rect 17736 3476 17742 3488
rect 17773 3485 17785 3488
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18012 3488 18521 3516
rect 18012 3476 18018 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 18656 3488 19257 3516
rect 18656 3476 18662 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 19484 3488 20085 3516
rect 19484 3476 19490 3488
rect 20073 3485 20085 3488
rect 20119 3485 20131 3519
rect 20073 3479 20131 3485
rect 20533 3519 20591 3525
rect 20533 3485 20545 3519
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 18782 3448 18788 3460
rect 15028 3420 18788 3448
rect 18782 3408 18788 3420
rect 18840 3408 18846 3460
rect 20548 3448 20576 3479
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21177 3519 21235 3525
rect 21177 3516 21189 3519
rect 20772 3488 21189 3516
rect 20772 3476 20778 3488
rect 21177 3485 21189 3488
rect 21223 3485 21235 3519
rect 21177 3479 21235 3485
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3516 21327 3519
rect 21450 3516 21456 3528
rect 21315 3488 21456 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 21818 3516 21824 3528
rect 21779 3488 21824 3516
rect 21818 3476 21824 3488
rect 21876 3476 21882 3528
rect 23842 3516 23848 3528
rect 22066 3512 22876 3516
rect 23124 3512 23244 3516
rect 22066 3488 23244 3512
rect 23803 3488 23848 3516
rect 22066 3448 22094 3488
rect 22848 3484 23152 3488
rect 20548 3420 22094 3448
rect 23216 3448 23244 3488
rect 23842 3476 23848 3488
rect 23900 3476 23906 3528
rect 25148 3518 25176 3624
rect 25222 3544 25228 3596
rect 25280 3584 25286 3596
rect 29730 3584 29736 3596
rect 25280 3556 29736 3584
rect 25280 3544 25286 3556
rect 29730 3544 29736 3556
rect 29788 3544 29794 3596
rect 25056 3516 25176 3518
rect 27246 3516 27252 3528
rect 24412 3490 25176 3516
rect 24412 3488 25084 3490
rect 27207 3488 27252 3516
rect 24412 3448 24440 3488
rect 27246 3476 27252 3488
rect 27304 3476 27310 3528
rect 29840 3516 29868 3624
rect 30926 3612 30932 3664
rect 30984 3652 30990 3664
rect 32214 3652 32220 3664
rect 30984 3624 32220 3652
rect 30984 3612 30990 3624
rect 32214 3612 32220 3624
rect 32272 3612 32278 3664
rect 31478 3516 31484 3528
rect 29840 3488 31484 3516
rect 31478 3476 31484 3488
rect 31536 3476 31542 3528
rect 32214 3476 32220 3528
rect 32272 3516 32278 3528
rect 32401 3519 32459 3525
rect 32401 3516 32413 3519
rect 32272 3488 32413 3516
rect 32272 3476 32278 3488
rect 32401 3485 32413 3488
rect 32447 3485 32459 3519
rect 32401 3479 32459 3485
rect 23216 3420 24440 3448
rect 24486 3408 24492 3460
rect 24544 3448 24550 3460
rect 24857 3451 24915 3457
rect 24857 3448 24869 3451
rect 24544 3420 24869 3448
rect 24544 3408 24550 3420
rect 24857 3417 24869 3420
rect 24903 3417 24915 3451
rect 24857 3411 24915 3417
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 25593 3451 25651 3457
rect 25593 3448 25605 3451
rect 25372 3420 25605 3448
rect 25372 3408 25378 3420
rect 25593 3417 25605 3420
rect 25639 3417 25651 3451
rect 25593 3411 25651 3417
rect 25685 3451 25743 3457
rect 25685 3417 25697 3451
rect 25731 3417 25743 3451
rect 25685 3411 25743 3417
rect 26605 3451 26663 3457
rect 26605 3417 26617 3451
rect 26651 3448 26663 3451
rect 27798 3448 27804 3460
rect 26651 3420 27804 3448
rect 26651 3417 26663 3420
rect 26605 3411 26663 3417
rect 16390 3380 16396 3392
rect 7760 3352 16396 3380
rect 7653 3343 7711 3349
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 16577 3383 16635 3389
rect 16577 3349 16589 3383
rect 16623 3380 16635 3383
rect 16666 3380 16672 3392
rect 16623 3352 16672 3380
rect 16623 3349 16635 3352
rect 16577 3343 16635 3349
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 17828 3352 17877 3380
rect 17828 3340 17834 3352
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 17865 3343 17923 3349
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18564 3352 18613 3380
rect 18564 3340 18570 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 19337 3383 19395 3389
rect 19337 3349 19349 3383
rect 19383 3380 19395 3383
rect 19978 3380 19984 3392
rect 19383 3352 19984 3380
rect 19383 3349 19395 3352
rect 19337 3343 19395 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 20622 3380 20628 3392
rect 20583 3352 20628 3380
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 22830 3380 22836 3392
rect 20772 3352 22836 3380
rect 20772 3340 20778 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 25700 3380 25728 3411
rect 27798 3408 27804 3420
rect 27856 3408 27862 3460
rect 35866 3448 35894 3692
rect 38565 3689 38577 3723
rect 38611 3720 38623 3723
rect 38654 3720 38660 3732
rect 38611 3692 38660 3720
rect 38611 3689 38623 3692
rect 38565 3683 38623 3689
rect 38654 3680 38660 3692
rect 38712 3680 38718 3732
rect 39390 3680 39396 3732
rect 39448 3720 39454 3732
rect 39448 3692 45692 3720
rect 39448 3680 39454 3692
rect 39117 3655 39175 3661
rect 39117 3621 39129 3655
rect 39163 3652 39175 3655
rect 40310 3652 40316 3664
rect 39163 3624 40316 3652
rect 39163 3621 39175 3624
rect 39117 3615 39175 3621
rect 40310 3612 40316 3624
rect 40368 3612 40374 3664
rect 40497 3655 40555 3661
rect 40497 3621 40509 3655
rect 40543 3652 40555 3655
rect 40586 3652 40592 3664
rect 40543 3624 40592 3652
rect 40543 3621 40555 3624
rect 40497 3615 40555 3621
rect 40586 3612 40592 3624
rect 40644 3612 40650 3664
rect 43806 3652 43812 3664
rect 42628 3624 43812 3652
rect 37550 3544 37556 3596
rect 37608 3584 37614 3596
rect 40957 3587 41015 3593
rect 40957 3584 40969 3587
rect 37608 3556 40969 3584
rect 37608 3544 37614 3556
rect 38470 3516 38476 3528
rect 38431 3488 38476 3516
rect 38470 3476 38476 3488
rect 38528 3476 38534 3528
rect 39298 3516 39304 3528
rect 39259 3488 39304 3516
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 39868 3525 39896 3556
rect 40957 3553 40969 3556
rect 41003 3584 41015 3587
rect 41874 3584 41880 3596
rect 41003 3556 41880 3584
rect 41003 3553 41015 3556
rect 40957 3547 41015 3553
rect 41874 3544 41880 3556
rect 41932 3544 41938 3596
rect 42628 3593 42656 3624
rect 43806 3612 43812 3624
rect 43864 3612 43870 3664
rect 42613 3587 42671 3593
rect 42613 3553 42625 3587
rect 42659 3553 42671 3587
rect 42794 3584 42800 3596
rect 42755 3556 42800 3584
rect 42613 3547 42671 3553
rect 42794 3544 42800 3556
rect 42852 3544 42858 3596
rect 43162 3584 43168 3596
rect 43123 3556 43168 3584
rect 43162 3544 43168 3556
rect 43220 3544 43226 3596
rect 39853 3519 39911 3525
rect 39853 3485 39865 3519
rect 39899 3485 39911 3519
rect 39853 3479 39911 3485
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 40000 3488 40049 3516
rect 40000 3476 40006 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 41141 3519 41199 3525
rect 41141 3485 41153 3519
rect 41187 3516 41199 3519
rect 41782 3516 41788 3528
rect 41187 3488 41788 3516
rect 41187 3485 41199 3488
rect 41141 3479 41199 3485
rect 41782 3476 41788 3488
rect 41840 3476 41846 3528
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45664 3525 45692 3692
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 40494 3448 40500 3460
rect 35866 3420 40500 3448
rect 40494 3408 40500 3420
rect 40552 3408 40558 3460
rect 42518 3408 42524 3460
rect 42576 3448 42582 3460
rect 43990 3448 43996 3460
rect 42576 3420 43996 3448
rect 42576 3408 42582 3420
rect 43990 3408 43996 3420
rect 44048 3408 44054 3460
rect 45741 3451 45799 3457
rect 45741 3417 45753 3451
rect 45787 3448 45799 3451
rect 46477 3451 46535 3457
rect 46477 3448 46489 3451
rect 45787 3420 46489 3448
rect 45787 3417 45799 3420
rect 45741 3411 45799 3417
rect 46477 3417 46489 3420
rect 46523 3417 46535 3451
rect 46477 3411 46535 3417
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 27065 3383 27123 3389
rect 27065 3380 27077 3383
rect 25700 3352 27077 3380
rect 27065 3349 27077 3352
rect 27111 3349 27123 3383
rect 27065 3343 27123 3349
rect 27430 3340 27436 3392
rect 27488 3380 27494 3392
rect 31110 3380 31116 3392
rect 27488 3352 31116 3380
rect 27488 3340 27494 3352
rect 31110 3340 31116 3352
rect 31168 3340 31174 3392
rect 31573 3383 31631 3389
rect 31573 3349 31585 3383
rect 31619 3380 31631 3383
rect 32398 3380 32404 3392
rect 31619 3352 32404 3380
rect 31619 3349 31631 3352
rect 31573 3343 31631 3349
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 37642 3340 37648 3392
rect 37700 3380 37706 3392
rect 41414 3380 41420 3392
rect 37700 3352 41420 3380
rect 37700 3340 37706 3352
rect 41414 3340 41420 3352
rect 41472 3340 41478 3392
rect 41601 3383 41659 3389
rect 41601 3349 41613 3383
rect 41647 3380 41659 3383
rect 42426 3380 42432 3392
rect 41647 3352 42432 3380
rect 41647 3349 41659 3352
rect 41601 3343 41659 3349
rect 42426 3340 42432 3352
rect 42484 3340 42490 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 9950 3176 9956 3188
rect 4120 3148 9956 3176
rect 4120 3136 4126 3148
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 16758 3176 16764 3188
rect 10060 3148 14136 3176
rect 16719 3148 16764 3176
rect 2038 3108 2044 3120
rect 1999 3080 2044 3108
rect 2038 3068 2044 3080
rect 2096 3068 2102 3120
rect 7466 3108 7472 3120
rect 7427 3080 7472 3108
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 10060 3049 10088 3148
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 11698 3108 11704 3120
rect 10192 3080 10237 3108
rect 11659 3080 11704 3108
rect 10192 3068 10198 3080
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 13998 3108 14004 3120
rect 13959 3080 14004 3108
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 14108 3108 14136 3148
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 17954 3176 17960 3188
rect 17915 3148 17960 3176
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18598 3176 18604 3188
rect 18559 3148 18604 3176
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 20714 3176 20720 3188
rect 18708 3148 20720 3176
rect 18708 3108 18736 3148
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 20864 3148 22094 3176
rect 20864 3136 20870 3148
rect 14108 3080 18736 3108
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 20622 3108 20628 3120
rect 19659 3080 20628 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 22066 3108 22094 3148
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 26145 3179 26203 3185
rect 22244 3148 25820 3176
rect 22244 3136 22250 3148
rect 22554 3108 22560 3120
rect 22066 3080 22560 3108
rect 22554 3068 22560 3080
rect 22612 3068 22618 3120
rect 25590 3108 25596 3120
rect 22664 3080 25596 3108
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3009 10103 3043
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 10045 3003 10103 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17862 3040 17868 3052
rect 17823 3012 17868 3040
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 19426 3040 19432 3052
rect 19387 3012 19432 3040
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 22189 3043 22247 3049
rect 22189 3040 22201 3043
rect 21968 3012 22201 3040
rect 21968 3000 21974 3012
rect 22189 3009 22201 3012
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2317 2975 2375 2981
rect 2317 2972 2329 2975
rect 716 2944 2329 2972
rect 716 2932 722 2944
rect 2317 2941 2329 2944
rect 2363 2941 2375 2975
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 2317 2935 2375 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11992 2904 12020 2935
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 19702 2972 19708 2984
rect 14884 2944 19708 2972
rect 14884 2932 14890 2944
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 19886 2972 19892 2984
rect 19847 2944 19892 2972
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 19978 2932 19984 2984
rect 20036 2972 20042 2984
rect 20162 2972 20168 2984
rect 20036 2944 20168 2972
rect 20036 2932 20042 2944
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 20346 2932 20352 2984
rect 20404 2972 20410 2984
rect 22664 2972 22692 3080
rect 25590 3068 25596 3080
rect 25648 3108 25654 3120
rect 25792 3108 25820 3148
rect 26145 3145 26157 3179
rect 26191 3176 26203 3179
rect 27246 3176 27252 3188
rect 26191 3148 27252 3176
rect 26191 3145 26203 3148
rect 26145 3139 26203 3145
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 27338 3136 27344 3188
rect 27396 3176 27402 3188
rect 27525 3179 27583 3185
rect 27525 3176 27537 3179
rect 27396 3148 27537 3176
rect 27396 3136 27402 3148
rect 27525 3145 27537 3148
rect 27571 3145 27583 3179
rect 36722 3176 36728 3188
rect 36683 3148 36728 3176
rect 27525 3139 27583 3145
rect 36722 3136 36728 3148
rect 36780 3136 36786 3188
rect 39298 3136 39304 3188
rect 39356 3176 39362 3188
rect 39945 3179 40003 3185
rect 39945 3176 39957 3179
rect 39356 3148 39957 3176
rect 39356 3136 39362 3148
rect 39945 3145 39957 3148
rect 39991 3145 40003 3179
rect 39945 3139 40003 3145
rect 40402 3136 40408 3188
rect 40460 3136 40466 3188
rect 40957 3179 41015 3185
rect 40957 3145 40969 3179
rect 41003 3176 41015 3179
rect 41003 3148 41644 3176
rect 41003 3145 41015 3148
rect 40957 3139 41015 3145
rect 27706 3108 27712 3120
rect 25648 3080 25728 3108
rect 25792 3080 27712 3108
rect 25648 3068 25654 3080
rect 22830 3040 22836 3052
rect 22791 3012 22836 3040
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 25700 3049 25728 3080
rect 27706 3068 27712 3080
rect 27764 3068 27770 3120
rect 32122 3108 32128 3120
rect 31726 3080 32128 3108
rect 25685 3043 25743 3049
rect 25685 3009 25697 3043
rect 25731 3009 25743 3043
rect 25685 3003 25743 3009
rect 25774 3000 25780 3052
rect 25832 3040 25838 3052
rect 26234 3040 26240 3052
rect 25832 3012 26240 3040
rect 25832 3000 25838 3012
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 27062 3000 27068 3052
rect 27120 3040 27126 3052
rect 27433 3043 27491 3049
rect 27433 3040 27445 3043
rect 27120 3012 27445 3040
rect 27120 3000 27126 3012
rect 27433 3009 27445 3012
rect 27479 3009 27491 3043
rect 27433 3003 27491 3009
rect 20404 2944 22692 2972
rect 23017 2975 23075 2981
rect 20404 2932 20410 2944
rect 23017 2941 23029 2975
rect 23063 2972 23075 2975
rect 23566 2972 23572 2984
rect 23063 2944 23428 2972
rect 23527 2944 23572 2972
rect 23063 2941 23075 2944
rect 23017 2935 23075 2941
rect 22186 2904 22192 2916
rect 11020 2876 12020 2904
rect 12406 2876 22192 2904
rect 11020 2864 11026 2876
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 12406 2836 12434 2876
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 22370 2904 22376 2916
rect 22331 2876 22376 2904
rect 22370 2864 22376 2876
rect 22428 2864 22434 2916
rect 23400 2904 23428 2944
rect 23566 2932 23572 2944
rect 23624 2932 23630 2984
rect 27614 2972 27620 2984
rect 25792 2944 27620 2972
rect 25792 2904 25820 2944
rect 27614 2932 27620 2944
rect 27672 2932 27678 2984
rect 23400 2876 25820 2904
rect 26234 2864 26240 2916
rect 26292 2904 26298 2916
rect 31726 2904 31754 3080
rect 32122 3068 32128 3080
rect 32180 3068 32186 3120
rect 32398 3108 32404 3120
rect 32359 3080 32404 3108
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 39577 3111 39635 3117
rect 39577 3077 39589 3111
rect 39623 3108 39635 3111
rect 40420 3108 40448 3136
rect 39623 3080 40448 3108
rect 39623 3077 39635 3080
rect 39577 3071 39635 3077
rect 41616 3073 41644 3148
rect 47026 3136 47032 3188
rect 47084 3176 47090 3188
rect 47857 3179 47915 3185
rect 47857 3176 47869 3179
rect 47084 3148 47869 3176
rect 47084 3136 47090 3148
rect 47857 3145 47869 3148
rect 47903 3145 47915 3179
rect 47857 3139 47915 3145
rect 41601 3067 41659 3073
rect 41690 3068 41696 3120
rect 41748 3108 41754 3120
rect 44450 3108 44456 3120
rect 41748 3080 44456 3108
rect 41748 3068 41754 3080
rect 44450 3068 44456 3080
rect 44508 3068 44514 3120
rect 45373 3111 45431 3117
rect 45373 3077 45385 3111
rect 45419 3108 45431 3111
rect 46750 3108 46756 3120
rect 45419 3080 46756 3108
rect 45419 3077 45431 3080
rect 45373 3071 45431 3077
rect 46750 3068 46756 3080
rect 46808 3068 46814 3120
rect 32214 3040 32220 3052
rect 32175 3012 32220 3040
rect 32214 3000 32220 3012
rect 32272 3000 32278 3052
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3040 36323 3043
rect 37642 3040 37648 3052
rect 36311 3012 37648 3040
rect 36311 3009 36323 3012
rect 36265 3003 36323 3009
rect 37642 3000 37648 3012
rect 37700 3000 37706 3052
rect 39114 3000 39120 3052
rect 39172 3040 39178 3052
rect 39761 3043 39819 3049
rect 39761 3040 39773 3043
rect 39172 3012 39773 3040
rect 39172 3000 39178 3012
rect 39761 3009 39773 3012
rect 39807 3040 39819 3043
rect 39942 3040 39948 3052
rect 39807 3012 39948 3040
rect 39807 3009 39819 3012
rect 39761 3003 39819 3009
rect 39942 3000 39948 3012
rect 40000 3040 40006 3052
rect 40405 3044 40463 3049
rect 41506 3044 41512 3052
rect 40328 3043 40463 3044
rect 40328 3040 40417 3043
rect 40000 3016 40417 3040
rect 40000 3012 40356 3016
rect 40000 3000 40006 3012
rect 40405 3009 40417 3016
rect 40451 3009 40463 3043
rect 41432 3040 41512 3044
rect 40405 3003 40463 3009
rect 40604 3016 41512 3040
rect 40604 3012 41460 3016
rect 33413 2975 33471 2981
rect 33413 2941 33425 2975
rect 33459 2972 33471 2975
rect 40604 2972 40632 3012
rect 41506 3000 41512 3016
rect 41564 3000 41570 3052
rect 41601 3033 41613 3067
rect 41647 3033 41659 3067
rect 42426 3040 42432 3052
rect 41601 3027 41659 3033
rect 42387 3012 42432 3040
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3040 47823 3043
rect 48314 3040 48320 3052
rect 47811 3012 48320 3040
rect 47811 3009 47823 3012
rect 47765 3003 47823 3009
rect 48314 3000 48320 3012
rect 48372 3000 48378 3052
rect 33459 2944 33548 2972
rect 33459 2941 33471 2944
rect 33413 2935 33471 2941
rect 33520 2916 33548 2944
rect 35866 2944 40632 2972
rect 40681 2975 40739 2981
rect 26292 2876 31754 2904
rect 26292 2864 26298 2876
rect 33502 2864 33508 2916
rect 33560 2864 33566 2916
rect 3936 2808 12434 2836
rect 3936 2796 3942 2808
rect 13446 2796 13452 2848
rect 13504 2836 13510 2848
rect 20806 2836 20812 2848
rect 13504 2808 20812 2836
rect 13504 2796 13510 2808
rect 20806 2796 20812 2808
rect 20864 2796 20870 2848
rect 20898 2796 20904 2848
rect 20956 2836 20962 2848
rect 22094 2836 22100 2848
rect 20956 2808 22100 2836
rect 20956 2796 20962 2808
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 25774 2836 25780 2848
rect 25735 2808 25780 2836
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 26142 2796 26148 2848
rect 26200 2836 26206 2848
rect 35866 2836 35894 2944
rect 40681 2941 40693 2975
rect 40727 2972 40739 2975
rect 41782 2972 41788 2984
rect 40727 2944 41788 2972
rect 40727 2941 40739 2944
rect 40681 2935 40739 2941
rect 41782 2932 41788 2944
rect 41840 2932 41846 2984
rect 42613 2975 42671 2981
rect 42613 2941 42625 2975
rect 42659 2941 42671 2975
rect 42613 2935 42671 2941
rect 42889 2975 42947 2981
rect 42889 2941 42901 2975
rect 42935 2941 42947 2975
rect 42889 2935 42947 2941
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 41417 2907 41475 2913
rect 41417 2873 41429 2907
rect 41463 2904 41475 2907
rect 42628 2904 42656 2935
rect 41463 2876 42656 2904
rect 41463 2873 41475 2876
rect 41417 2867 41475 2873
rect 26200 2808 35894 2836
rect 26200 2796 26206 2808
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 36357 2839 36415 2845
rect 36357 2836 36369 2839
rect 36228 2808 36369 2836
rect 36228 2796 36234 2808
rect 36357 2805 36369 2808
rect 36403 2805 36415 2839
rect 36357 2799 36415 2805
rect 40402 2796 40408 2848
rect 40460 2836 40466 2848
rect 40497 2839 40555 2845
rect 40497 2836 40509 2839
rect 40460 2808 40509 2836
rect 40460 2796 40466 2808
rect 40497 2805 40509 2808
rect 40543 2805 40555 2839
rect 40497 2799 40555 2805
rect 40586 2796 40592 2848
rect 40644 2836 40650 2848
rect 42904 2836 42932 2935
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 40644 2808 42932 2836
rect 40644 2796 40650 2808
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5307 2604 9536 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 2774 2564 2780 2576
rect 1412 2536 2780 2564
rect 1412 2505 1440 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 6638 2524 6644 2576
rect 6696 2564 6702 2576
rect 9508 2564 9536 2604
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 9640 2604 17540 2632
rect 9640 2592 9646 2604
rect 12342 2564 12348 2576
rect 6696 2536 7052 2564
rect 9508 2536 12348 2564
rect 6696 2524 6702 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2866 2496 2872 2508
rect 2827 2468 2872 2496
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 6454 2456 6460 2508
rect 6512 2496 6518 2508
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 6512 2468 6561 2496
rect 6512 2456 6518 2468
rect 6549 2465 6561 2468
rect 6595 2465 6607 2499
rect 6549 2459 6607 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6914 2496 6920 2508
rect 6779 2468 6920 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7024 2505 7052 2536
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 16482 2524 16488 2576
rect 16540 2564 16546 2576
rect 17313 2567 17371 2573
rect 17313 2564 17325 2567
rect 16540 2536 17325 2564
rect 16540 2524 16546 2536
rect 17313 2533 17325 2536
rect 17359 2533 17371 2567
rect 17512 2564 17540 2604
rect 17586 2592 17592 2644
rect 17644 2632 17650 2644
rect 17865 2635 17923 2641
rect 17865 2632 17877 2635
rect 17644 2604 17877 2632
rect 17644 2592 17650 2604
rect 17865 2601 17877 2604
rect 17911 2601 17923 2635
rect 17865 2595 17923 2601
rect 18322 2592 18328 2644
rect 18380 2632 18386 2644
rect 18509 2635 18567 2641
rect 18509 2632 18521 2635
rect 18380 2604 18521 2632
rect 18380 2592 18386 2604
rect 18509 2601 18521 2604
rect 18555 2601 18567 2635
rect 18509 2595 18567 2601
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 19702 2632 19708 2644
rect 19383 2604 19708 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 19702 2592 19708 2604
rect 19760 2592 19766 2644
rect 19981 2635 20039 2641
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 20070 2632 20076 2644
rect 20027 2604 20076 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20254 2592 20260 2644
rect 20312 2632 20318 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20312 2604 20913 2632
rect 20312 2592 20318 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 23658 2632 23664 2644
rect 20901 2595 20959 2601
rect 21008 2604 23664 2632
rect 21008 2564 21036 2604
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 26050 2592 26056 2644
rect 26108 2632 26114 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 26108 2604 28641 2632
rect 26108 2592 26114 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 28629 2595 28687 2601
rect 29733 2635 29791 2641
rect 29733 2601 29745 2635
rect 29779 2632 29791 2635
rect 31754 2632 31760 2644
rect 29779 2604 31760 2632
rect 29779 2601 29791 2604
rect 29733 2595 29791 2601
rect 31754 2592 31760 2604
rect 31812 2592 31818 2644
rect 32122 2592 32128 2644
rect 32180 2632 32186 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 32180 2604 35541 2632
rect 32180 2592 32186 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 36354 2632 36360 2644
rect 36315 2604 36360 2632
rect 35529 2595 35587 2601
rect 36354 2592 36360 2604
rect 36412 2592 36418 2644
rect 39114 2632 39120 2644
rect 39075 2604 39120 2632
rect 39114 2592 39120 2604
rect 39172 2592 39178 2644
rect 41693 2635 41751 2641
rect 41693 2601 41705 2635
rect 41739 2632 41751 2635
rect 41782 2632 41788 2644
rect 41739 2604 41788 2632
rect 41739 2601 41751 2604
rect 41693 2595 41751 2601
rect 41782 2592 41788 2604
rect 41840 2592 41846 2644
rect 17512 2536 21036 2564
rect 22005 2567 22063 2573
rect 17313 2527 17371 2533
rect 22005 2533 22017 2567
rect 22051 2564 22063 2567
rect 25406 2564 25412 2576
rect 22051 2536 25412 2564
rect 22051 2533 22063 2536
rect 22005 2527 22063 2533
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 22020 2496 22048 2527
rect 25406 2524 25412 2536
rect 25464 2524 25470 2576
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 45557 2567 45615 2573
rect 45557 2564 45569 2567
rect 28960 2536 45569 2564
rect 28960 2524 28966 2536
rect 45557 2533 45569 2536
rect 45603 2533 45615 2567
rect 45557 2527 45615 2533
rect 11756 2468 22048 2496
rect 11756 2456 11762 2468
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22336 2468 22876 2496
rect 22336 2456 22342 2468
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2792 2400 3801 2428
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2792 2360 2820 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 15010 2428 15016 2440
rect 5445 2391 5503 2397
rect 8312 2400 15016 2428
rect 8312 2360 8340 2400
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15470 2428 15476 2440
rect 15335 2400 15476 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 17770 2428 17776 2440
rect 15620 2400 15665 2428
rect 17731 2400 17776 2428
rect 15620 2388 15626 2400
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 18230 2388 18236 2440
rect 18288 2428 18294 2440
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18288 2400 18429 2428
rect 18288 2388 18294 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19794 2428 19800 2440
rect 19291 2400 19800 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 19794 2388 19800 2400
rect 19852 2388 19858 2440
rect 19889 2431 19947 2437
rect 19889 2397 19901 2431
rect 19935 2428 19947 2431
rect 20070 2428 20076 2440
rect 19935 2400 20076 2428
rect 19935 2397 19947 2400
rect 19889 2391 19947 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 22370 2428 22376 2440
rect 22331 2400 22376 2428
rect 22370 2388 22376 2400
rect 22428 2388 22434 2440
rect 22848 2437 22876 2468
rect 23842 2456 23848 2508
rect 23900 2496 23906 2508
rect 24489 2499 24547 2505
rect 24489 2496 24501 2499
rect 23900 2468 24501 2496
rect 23900 2456 23906 2468
rect 24489 2465 24501 2468
rect 24535 2465 24547 2499
rect 24670 2496 24676 2508
rect 24631 2468 24676 2496
rect 24489 2459 24547 2465
rect 24670 2456 24676 2468
rect 24728 2456 24734 2508
rect 25130 2496 25136 2508
rect 25091 2468 25136 2496
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 27154 2456 27160 2508
rect 27212 2496 27218 2508
rect 27249 2499 27307 2505
rect 27249 2496 27261 2499
rect 27212 2468 27261 2496
rect 27212 2456 27218 2468
rect 27249 2465 27261 2468
rect 27295 2465 27307 2499
rect 27249 2459 27307 2465
rect 33134 2456 33140 2508
rect 33192 2496 33198 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 33192 2468 40509 2496
rect 33192 2456 33198 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 41966 2456 41972 2508
rect 42024 2496 42030 2508
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 42024 2468 46489 2496
rect 42024 2456 42030 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 46477 2459 46535 2465
rect 46566 2456 46572 2508
rect 46624 2496 46630 2508
rect 47857 2499 47915 2505
rect 47857 2496 47869 2499
rect 46624 2468 47869 2496
rect 46624 2456 46630 2468
rect 47857 2465 47869 2468
rect 47903 2465 47915 2499
rect 47857 2459 47915 2465
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 38068 2400 38117 2428
rect 38068 2388 38074 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39301 2431 39359 2437
rect 39301 2397 39313 2431
rect 39347 2428 39359 2431
rect 39942 2428 39948 2440
rect 39347 2400 39948 2428
rect 39347 2397 39359 2400
rect 39301 2391 39359 2397
rect 39942 2388 39948 2400
rect 40000 2388 40006 2440
rect 41230 2388 41236 2440
rect 41288 2428 41294 2440
rect 41877 2431 41935 2437
rect 41877 2428 41889 2431
rect 41288 2400 41889 2428
rect 41288 2388 41294 2400
rect 41877 2397 41889 2400
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 46201 2431 46259 2437
rect 46201 2397 46213 2431
rect 46247 2428 46259 2431
rect 47026 2428 47032 2440
rect 46247 2400 47032 2428
rect 46247 2397 46259 2400
rect 46201 2391 46259 2397
rect 2648 2332 2820 2360
rect 3988 2332 8340 2360
rect 2648 2320 2654 2332
rect 3988 2301 4016 2332
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8444 2332 9413 2360
rect 8444 2320 8450 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16172 2332 17141 2360
rect 16172 2320 16178 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 39390 2320 39396 2372
rect 39448 2360 39454 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39448 2332 40325 2360
rect 39448 2320 39454 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41049 2363 41107 2369
rect 41049 2360 41061 2363
rect 40644 2332 41061 2360
rect 40644 2320 40650 2332
rect 41049 2329 41061 2332
rect 41095 2329 41107 2363
rect 41049 2323 41107 2329
rect 41414 2320 41420 2372
rect 41472 2360 41478 2372
rect 43916 2360 43944 2391
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 47673 2431 47731 2437
rect 47673 2397 47685 2431
rect 47719 2428 47731 2431
rect 48038 2428 48044 2440
rect 47719 2400 48044 2428
rect 47719 2397 47731 2400
rect 47673 2391 47731 2397
rect 48038 2388 48044 2400
rect 48096 2388 48102 2440
rect 41472 2332 43944 2360
rect 45373 2363 45431 2369
rect 41472 2320 41478 2332
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46750 2360 46756 2372
rect 45419 2332 46756 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46750 2320 46756 2332
rect 46808 2320 46814 2372
rect 3973 2295 4031 2301
rect 3973 2261 3985 2295
rect 4019 2261 4031 2295
rect 9674 2292 9680 2304
rect 9635 2264 9680 2292
rect 3973 2255 4031 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 31846 2252 31852 2304
rect 31904 2292 31910 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 31904 2264 38301 2292
rect 31904 2252 31910 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 38289 2255 38347 2261
rect 41141 2295 41199 2301
rect 41141 2261 41153 2295
rect 41187 2292 41199 2295
rect 43254 2292 43260 2304
rect 41187 2264 43260 2292
rect 41187 2261 41199 2264
rect 41141 2255 41199 2261
rect 43254 2252 43260 2264
rect 43312 2252 43318 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 3510 2048 3516 2100
rect 3568 2088 3574 2100
rect 9582 2088 9588 2100
rect 3568 2060 9588 2088
rect 3568 2048 3574 2060
rect 9582 2048 9588 2060
rect 9640 2048 9646 2100
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 23934 2088 23940 2100
rect 9732 2060 23940 2088
rect 9732 2048 9738 2060
rect 23934 2048 23940 2060
rect 23992 2048 23998 2100
rect 2958 1980 2964 2032
rect 3016 2020 3022 2032
rect 11698 2020 11704 2032
rect 3016 1992 11704 2020
rect 3016 1980 3022 1992
rect 11698 1980 11704 1992
rect 11756 1980 11762 2032
rect 15562 1980 15568 2032
rect 15620 2020 15626 2032
rect 36170 2020 36176 2032
rect 15620 1992 36176 2020
rect 15620 1980 15626 1992
rect 36170 1980 36176 1992
rect 36228 1980 36234 2032
rect 22554 1368 22560 1420
rect 22612 1408 22618 1420
rect 23566 1408 23572 1420
rect 22612 1380 23572 1408
rect 22612 1368 22618 1380
rect 23566 1368 23572 1380
rect 23624 1368 23630 1420
<< via1 >>
rect 15936 47540 15988 47592
rect 20076 47540 20128 47592
rect 20260 47540 20312 47592
rect 28264 47540 28316 47592
rect 3056 47472 3108 47524
rect 35440 47472 35492 47524
rect 2044 47404 2096 47456
rect 40132 47404 40184 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 3056 47243 3108 47252
rect 3056 47209 3065 47243
rect 3065 47209 3099 47243
rect 3099 47209 3108 47243
rect 3056 47200 3108 47209
rect 3332 47200 3384 47252
rect 21824 47200 21876 47252
rect 29000 47200 29052 47252
rect 30196 47200 30248 47252
rect 41696 47200 41748 47252
rect 46848 47200 46900 47252
rect 20260 47132 20312 47184
rect 20352 47132 20404 47184
rect 2044 47107 2096 47116
rect 2044 47073 2053 47107
rect 2053 47073 2087 47107
rect 2087 47073 2096 47107
rect 2044 47064 2096 47073
rect 11612 47064 11664 47116
rect 1952 46996 2004 47048
rect 3240 46996 3292 47048
rect 4804 47039 4856 47048
rect 4804 47005 4813 47039
rect 4813 47005 4847 47039
rect 4847 47005 4856 47039
rect 4804 46996 4856 47005
rect 5816 46996 5868 47048
rect 7380 47039 7432 47048
rect 7380 47005 7389 47039
rect 7389 47005 7423 47039
rect 7423 47005 7432 47039
rect 7380 46996 7432 47005
rect 9036 46996 9088 47048
rect 12900 46996 12952 47048
rect 13820 47064 13872 47116
rect 17408 47064 17460 47116
rect 20076 47064 20128 47116
rect 47860 47132 47912 47184
rect 14464 46996 14516 47048
rect 16580 46996 16632 47048
rect 18604 46996 18656 47048
rect 21088 47039 21140 47048
rect 21088 47005 21097 47039
rect 21097 47005 21131 47039
rect 21131 47005 21140 47039
rect 21088 46996 21140 47005
rect 22008 47039 22060 47048
rect 22008 47005 22017 47039
rect 22017 47005 22051 47039
rect 22051 47005 22060 47039
rect 22008 46996 22060 47005
rect 4068 46971 4120 46980
rect 2596 46860 2648 46912
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 6644 46971 6696 46980
rect 6644 46937 6653 46971
rect 6653 46937 6687 46971
rect 6687 46937 6696 46971
rect 6644 46928 6696 46937
rect 7472 46928 7524 46980
rect 9496 46928 9548 46980
rect 19432 46928 19484 46980
rect 16120 46860 16172 46912
rect 16580 46860 16632 46912
rect 18696 46860 18748 46912
rect 19984 46928 20036 46980
rect 24584 46996 24636 47048
rect 25504 47039 25556 47048
rect 25504 47005 25513 47039
rect 25513 47005 25547 47039
rect 25547 47005 25556 47039
rect 25504 46996 25556 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 30932 46996 30984 47048
rect 38108 46996 38160 47048
rect 42708 47039 42760 47048
rect 42708 47005 42717 47039
rect 42717 47005 42751 47039
rect 42751 47005 42760 47039
rect 42708 46996 42760 47005
rect 44456 47064 44508 47116
rect 48320 47064 48372 47116
rect 43812 46996 43864 47048
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 20168 46860 20220 46912
rect 27804 46928 27856 46980
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 43352 46928 43404 46980
rect 45468 46928 45520 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 3884 46588 3936 46640
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 22008 46588 22060 46640
rect 24584 46563 24636 46572
rect 24584 46529 24593 46563
rect 24593 46529 24627 46563
rect 24627 46529 24636 46563
rect 24584 46520 24636 46529
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 47952 46563 48004 46572
rect 47952 46529 47961 46563
rect 47961 46529 47995 46563
rect 47995 46529 48004 46563
rect 47952 46520 48004 46529
rect 3976 46495 4028 46504
rect 3976 46461 3985 46495
rect 3985 46461 4019 46495
rect 4019 46461 4028 46495
rect 3976 46452 4028 46461
rect 5080 46452 5132 46504
rect 12072 46452 12124 46504
rect 13544 46452 13596 46504
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 14280 46452 14332 46461
rect 20076 46452 20128 46504
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32312 46495 32364 46504
rect 32312 46461 32321 46495
rect 32321 46461 32355 46495
rect 32355 46461 32364 46495
rect 32312 46452 32364 46461
rect 38292 46495 38344 46504
rect 32220 46384 32272 46436
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 45376 46495 45428 46504
rect 42524 46384 42576 46436
rect 45376 46461 45385 46495
rect 45385 46461 45419 46495
rect 45419 46461 45428 46495
rect 45376 46452 45428 46461
rect 46756 46495 46808 46504
rect 46756 46461 46765 46495
rect 46765 46461 46799 46495
rect 46799 46461 46808 46495
rect 46756 46452 46808 46461
rect 45652 46384 45704 46436
rect 1676 46316 1728 46368
rect 10968 46316 11020 46368
rect 41328 46316 41380 46368
rect 48044 46359 48096 46368
rect 48044 46325 48053 46359
rect 48053 46325 48087 46359
rect 48087 46325 48096 46359
rect 48044 46316 48096 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3976 46112 4028 46164
rect 5080 46155 5132 46164
rect 5080 46121 5089 46155
rect 5089 46121 5123 46155
rect 5123 46121 5132 46155
rect 5080 46112 5132 46121
rect 13544 46155 13596 46164
rect 13544 46121 13553 46155
rect 13553 46121 13587 46155
rect 13587 46121 13596 46155
rect 13544 46112 13596 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 20076 46155 20128 46164
rect 20076 46121 20085 46155
rect 20085 46121 20119 46155
rect 20119 46121 20128 46155
rect 20076 46112 20128 46121
rect 24768 46112 24820 46164
rect 32312 46112 32364 46164
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 42616 46112 42668 46164
rect 45376 46112 45428 46164
rect 1768 45908 1820 45960
rect 21088 45976 21140 46028
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 12256 45908 12308 45960
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 20628 45908 20680 45960
rect 39948 46044 40000 46096
rect 25504 45976 25556 46028
rect 25780 46019 25832 46028
rect 25780 45985 25789 46019
rect 25789 45985 25823 46019
rect 25823 45985 25832 46019
rect 25780 45976 25832 45985
rect 41328 46019 41380 46028
rect 41328 45985 41337 46019
rect 41337 45985 41371 46019
rect 41371 45985 41380 46019
rect 41328 45976 41380 45985
rect 41880 46019 41932 46028
rect 41880 45985 41889 46019
rect 41889 45985 41923 46019
rect 41923 45985 41932 46019
rect 41880 45976 41932 45985
rect 31760 45951 31812 45960
rect 21088 45840 21140 45892
rect 12348 45815 12400 45824
rect 12348 45781 12357 45815
rect 12357 45781 12391 45815
rect 12391 45781 12400 45815
rect 12348 45772 12400 45781
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 31760 45917 31769 45951
rect 31769 45917 31803 45951
rect 31803 45917 31812 45951
rect 31760 45908 31812 45917
rect 39948 45908 40000 45960
rect 45744 45976 45796 46028
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 46296 45951 46348 45960
rect 41512 45883 41564 45892
rect 41512 45849 41521 45883
rect 41521 45849 41555 45883
rect 41555 45849 41564 45883
rect 41512 45840 41564 45849
rect 46296 45917 46305 45951
rect 46305 45917 46339 45951
rect 46339 45917 46348 45951
rect 46296 45908 46348 45917
rect 45376 45840 45428 45892
rect 45836 45883 45888 45892
rect 45836 45849 45845 45883
rect 45845 45849 45879 45883
rect 45879 45849 45888 45883
rect 45836 45840 45888 45849
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 45100 45772 45152 45824
rect 45560 45772 45612 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 12072 45611 12124 45620
rect 12072 45577 12081 45611
rect 12081 45577 12115 45611
rect 12115 45577 12124 45611
rect 12072 45568 12124 45577
rect 21088 45611 21140 45620
rect 21088 45577 21097 45611
rect 21097 45577 21131 45611
rect 21131 45577 21140 45611
rect 21088 45568 21140 45577
rect 25412 45611 25464 45620
rect 25412 45577 25421 45611
rect 25421 45577 25455 45611
rect 25455 45577 25464 45611
rect 25412 45568 25464 45577
rect 41512 45611 41564 45620
rect 41512 45577 41521 45611
rect 41521 45577 41555 45611
rect 41555 45577 41564 45611
rect 41512 45568 41564 45577
rect 46388 45568 46440 45620
rect 42800 45500 42852 45552
rect 1768 45475 1820 45484
rect 1768 45441 1777 45475
rect 1777 45441 1811 45475
rect 1811 45441 1820 45475
rect 1768 45432 1820 45441
rect 11980 45475 12032 45484
rect 11980 45441 11989 45475
rect 11989 45441 12023 45475
rect 12023 45441 12032 45475
rect 11980 45432 12032 45441
rect 31024 45432 31076 45484
rect 41420 45475 41472 45484
rect 41420 45441 41429 45475
rect 41429 45441 41463 45475
rect 41463 45441 41472 45475
rect 41420 45432 41472 45441
rect 2228 45364 2280 45416
rect 2780 45407 2832 45416
rect 2780 45373 2789 45407
rect 2789 45373 2823 45407
rect 2823 45373 2832 45407
rect 2780 45364 2832 45373
rect 42800 45407 42852 45416
rect 42800 45373 42809 45407
rect 42809 45373 42843 45407
rect 42843 45373 42852 45407
rect 42800 45364 42852 45373
rect 44088 45407 44140 45416
rect 44088 45373 44097 45407
rect 44097 45373 44131 45407
rect 44131 45373 44140 45407
rect 44088 45364 44140 45373
rect 45100 45407 45152 45416
rect 45100 45373 45109 45407
rect 45109 45373 45143 45407
rect 45143 45373 45152 45407
rect 45100 45364 45152 45373
rect 45652 45407 45704 45416
rect 45652 45373 45661 45407
rect 45661 45373 45695 45407
rect 45695 45373 45704 45407
rect 45652 45364 45704 45373
rect 43536 45296 43588 45348
rect 27252 45271 27304 45280
rect 27252 45237 27261 45271
rect 27261 45237 27295 45271
rect 27295 45237 27304 45271
rect 27252 45228 27304 45237
rect 47492 45228 47544 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 2228 45067 2280 45076
rect 2228 45033 2237 45067
rect 2237 45033 2271 45067
rect 2271 45033 2280 45067
rect 2228 45024 2280 45033
rect 42800 45067 42852 45076
rect 42800 45033 42809 45067
rect 42809 45033 42843 45067
rect 42843 45033 42852 45067
rect 42800 45024 42852 45033
rect 43536 45067 43588 45076
rect 43536 45033 43545 45067
rect 43545 45033 43579 45067
rect 43579 45033 43588 45067
rect 43536 45024 43588 45033
rect 45100 45024 45152 45076
rect 46480 45024 46532 45076
rect 46296 44956 46348 45008
rect 27252 44931 27304 44940
rect 27252 44897 27261 44931
rect 27261 44897 27295 44931
rect 27295 44897 27304 44931
rect 27252 44888 27304 44897
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 2320 44820 2372 44872
rect 27068 44863 27120 44872
rect 27068 44829 27077 44863
rect 27077 44829 27111 44863
rect 27111 44829 27120 44863
rect 27068 44820 27120 44829
rect 38660 44752 38712 44804
rect 45008 44820 45060 44872
rect 45376 44820 45428 44872
rect 46204 44752 46256 44804
rect 46480 44795 46532 44804
rect 46480 44761 46489 44795
rect 46489 44761 46523 44795
rect 46523 44761 46532 44795
rect 46480 44752 46532 44761
rect 47032 44684 47084 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 27068 44523 27120 44532
rect 27068 44489 27077 44523
rect 27077 44489 27111 44523
rect 27111 44489 27120 44523
rect 27068 44480 27120 44489
rect 46480 44480 46532 44532
rect 45468 44412 45520 44464
rect 25136 44344 25188 44396
rect 45192 44344 45244 44396
rect 45744 44387 45796 44396
rect 45744 44353 45753 44387
rect 45753 44353 45787 44387
rect 45787 44353 45796 44387
rect 45744 44344 45796 44353
rect 47584 44387 47636 44396
rect 41420 44276 41472 44328
rect 47584 44353 47593 44387
rect 47593 44353 47627 44387
rect 47627 44353 47636 44387
rect 47584 44344 47636 44353
rect 46940 44183 46992 44192
rect 46940 44149 46949 44183
rect 46949 44149 46983 44183
rect 46983 44149 46992 44183
rect 46940 44140 46992 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 46940 43800 46992 43852
rect 48228 43800 48280 43852
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 41236 43188 41288 43240
rect 47768 43095 47820 43104
rect 47768 43061 47777 43095
rect 47777 43061 47811 43095
rect 47811 43061 47820 43095
rect 47768 43052 47820 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47768 42712 47820 42764
rect 46940 42576 46992 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 46940 42347 46992 42356
rect 46940 42313 46949 42347
rect 46949 42313 46983 42347
rect 46983 42313 46992 42347
rect 46940 42304 46992 42313
rect 44364 42236 44416 42288
rect 45376 42236 45428 42288
rect 46204 42168 46256 42220
rect 46664 42168 46716 42220
rect 1400 41964 1452 42016
rect 46480 41964 46532 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 46480 41667 46532 41676
rect 46480 41633 46489 41667
rect 46489 41633 46523 41667
rect 46523 41633 46532 41667
rect 46480 41624 46532 41633
rect 48136 41599 48188 41608
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 47676 41488 47728 41540
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 14096 41080 14148 41132
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 47308 40876 47360 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 22928 40468 22980 40520
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 10324 40332 10376 40384
rect 22100 40375 22152 40384
rect 22100 40341 22109 40375
rect 22109 40341 22143 40375
rect 22143 40341 22152 40375
rect 22100 40332 22152 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 22928 40171 22980 40180
rect 22928 40137 22937 40171
rect 22937 40137 22971 40171
rect 22971 40137 22980 40171
rect 22928 40128 22980 40137
rect 20352 40103 20404 40112
rect 20352 40069 20361 40103
rect 20361 40069 20395 40103
rect 20395 40069 20404 40103
rect 20352 40060 20404 40069
rect 20536 40103 20588 40112
rect 20536 40069 20545 40103
rect 20545 40069 20579 40103
rect 20579 40069 20588 40103
rect 20536 40060 20588 40069
rect 45836 40060 45888 40112
rect 23112 39924 23164 39976
rect 20536 39856 20588 39908
rect 20352 39788 20404 39840
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 22100 39448 22152 39500
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 19984 39380 20036 39432
rect 21364 39423 21416 39432
rect 21364 39389 21373 39423
rect 21373 39389 21407 39423
rect 21407 39389 21416 39423
rect 21364 39380 21416 39389
rect 45008 39423 45060 39432
rect 45008 39389 45017 39423
rect 45017 39389 45051 39423
rect 45051 39389 45060 39423
rect 45008 39380 45060 39389
rect 22100 39312 22152 39364
rect 46940 39312 46992 39364
rect 20260 39244 20312 39296
rect 22928 39244 22980 39296
rect 45192 39244 45244 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 22100 39040 22152 39092
rect 23112 39083 23164 39092
rect 23112 39049 23121 39083
rect 23121 39049 23155 39083
rect 23155 39049 23164 39083
rect 23112 39040 23164 39049
rect 45192 39015 45244 39024
rect 19340 38904 19392 38956
rect 19984 38904 20036 38956
rect 20260 38904 20312 38956
rect 20444 38768 20496 38820
rect 45192 38981 45201 39015
rect 45201 38981 45235 39015
rect 45235 38981 45244 39015
rect 45192 38972 45244 38981
rect 46848 39015 46900 39024
rect 46848 38981 46857 39015
rect 46857 38981 46891 39015
rect 46891 38981 46900 39015
rect 46848 38972 46900 38981
rect 22928 38904 22980 38956
rect 22560 38836 22612 38888
rect 28816 38904 28868 38956
rect 43628 38947 43680 38956
rect 43628 38913 43637 38947
rect 43637 38913 43671 38947
rect 43671 38913 43680 38947
rect 43628 38904 43680 38913
rect 47768 38947 47820 38956
rect 47768 38913 47777 38947
rect 47777 38913 47811 38947
rect 47811 38913 47820 38947
rect 47768 38904 47820 38913
rect 44364 38879 44416 38888
rect 44364 38845 44373 38879
rect 44373 38845 44407 38879
rect 44407 38845 44416 38879
rect 44364 38836 44416 38845
rect 44640 38836 44692 38888
rect 23480 38700 23532 38752
rect 27896 38743 27948 38752
rect 27896 38709 27905 38743
rect 27905 38709 27939 38743
rect 27939 38709 27948 38743
rect 27896 38700 27948 38709
rect 47032 38700 47084 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 12348 38292 12400 38344
rect 16488 38335 16540 38344
rect 16488 38301 16497 38335
rect 16497 38301 16531 38335
rect 16531 38301 16540 38335
rect 16488 38292 16540 38301
rect 11980 38224 12032 38276
rect 27344 38496 27396 38548
rect 46940 38539 46992 38548
rect 46940 38505 46949 38539
rect 46949 38505 46983 38539
rect 46983 38505 46992 38539
rect 46940 38496 46992 38505
rect 20812 38360 20864 38412
rect 21364 38360 21416 38412
rect 27620 38360 27672 38412
rect 39120 38360 39172 38412
rect 39948 38360 40000 38412
rect 43628 38292 43680 38344
rect 46572 38292 46624 38344
rect 18972 38156 19024 38208
rect 20536 38224 20588 38276
rect 22192 38267 22244 38276
rect 22192 38233 22201 38267
rect 22201 38233 22235 38267
rect 22235 38233 22244 38267
rect 22192 38224 22244 38233
rect 23480 38224 23532 38276
rect 24768 38224 24820 38276
rect 25688 38224 25740 38276
rect 26976 38224 27028 38276
rect 27896 38224 27948 38276
rect 45928 38267 45980 38276
rect 45928 38233 45937 38267
rect 45937 38233 45971 38267
rect 45971 38233 45980 38267
rect 45928 38224 45980 38233
rect 19984 38156 20036 38208
rect 21272 38199 21324 38208
rect 21272 38165 21281 38199
rect 21281 38165 21315 38199
rect 21315 38165 21324 38199
rect 21272 38156 21324 38165
rect 22836 38156 22888 38208
rect 23204 38156 23256 38208
rect 25964 38156 26016 38208
rect 28356 38199 28408 38208
rect 28356 38165 28365 38199
rect 28365 38165 28399 38199
rect 28399 38165 28408 38199
rect 28356 38156 28408 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 2320 37884 2372 37936
rect 17500 37952 17552 38004
rect 18512 37952 18564 38004
rect 18696 37995 18748 38004
rect 18696 37961 18705 37995
rect 18705 37961 18739 37995
rect 18739 37961 18748 37995
rect 18696 37952 18748 37961
rect 20536 37952 20588 38004
rect 24768 37995 24820 38004
rect 24768 37961 24777 37995
rect 24777 37961 24811 37995
rect 24811 37961 24820 37995
rect 24768 37952 24820 37961
rect 25688 37952 25740 38004
rect 26976 37995 27028 38004
rect 26976 37961 26985 37995
rect 26985 37961 27019 37995
rect 27019 37961 27028 37995
rect 26976 37952 27028 37961
rect 17684 37884 17736 37936
rect 19248 37884 19300 37936
rect 19800 37884 19852 37936
rect 20168 37884 20220 37936
rect 45928 37884 45980 37936
rect 17316 37816 17368 37868
rect 18144 37859 18196 37868
rect 14464 37748 14516 37800
rect 18144 37825 18153 37859
rect 18153 37825 18187 37859
rect 18187 37825 18196 37859
rect 18144 37816 18196 37825
rect 18420 37859 18472 37868
rect 18420 37825 18429 37859
rect 18429 37825 18463 37859
rect 18463 37825 18472 37859
rect 18420 37816 18472 37825
rect 19432 37816 19484 37868
rect 19294 37748 19346 37800
rect 9496 37680 9548 37732
rect 14372 37680 14424 37732
rect 16856 37612 16908 37664
rect 18512 37612 18564 37664
rect 19248 37612 19300 37664
rect 20444 37816 20496 37868
rect 22836 37859 22888 37868
rect 22836 37825 22845 37859
rect 22845 37825 22879 37859
rect 22879 37825 22888 37859
rect 22836 37816 22888 37825
rect 23020 37816 23072 37868
rect 23204 37816 23256 37868
rect 24952 37859 25004 37868
rect 24952 37825 24961 37859
rect 24961 37825 24995 37859
rect 24995 37825 25004 37859
rect 24952 37816 25004 37825
rect 26976 37816 27028 37868
rect 27160 37859 27212 37868
rect 27160 37825 27169 37859
rect 27169 37825 27203 37859
rect 27203 37825 27212 37859
rect 27160 37816 27212 37825
rect 27528 37859 27580 37868
rect 19616 37680 19668 37732
rect 20168 37748 20220 37800
rect 22744 37748 22796 37800
rect 25964 37748 26016 37800
rect 27068 37748 27120 37800
rect 27528 37825 27537 37859
rect 27537 37825 27571 37859
rect 27571 37825 27580 37859
rect 27528 37816 27580 37825
rect 43628 37816 43680 37868
rect 44272 37816 44324 37868
rect 27344 37748 27396 37800
rect 44916 37748 44968 37800
rect 19984 37723 20036 37732
rect 19984 37689 19993 37723
rect 19993 37689 20027 37723
rect 20027 37689 20036 37723
rect 19984 37680 20036 37689
rect 20904 37612 20956 37664
rect 21272 37612 21324 37664
rect 23204 37612 23256 37664
rect 23296 37655 23348 37664
rect 23296 37621 23305 37655
rect 23305 37621 23339 37655
rect 23339 37621 23348 37655
rect 23296 37612 23348 37621
rect 23572 37612 23624 37664
rect 27436 37655 27488 37664
rect 27436 37621 27445 37655
rect 27445 37621 27479 37655
rect 27479 37621 27488 37655
rect 27436 37612 27488 37621
rect 47768 37655 47820 37664
rect 47768 37621 47777 37655
rect 47777 37621 47811 37655
rect 47811 37621 47820 37655
rect 47768 37612 47820 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 15936 37451 15988 37460
rect 15936 37417 15945 37451
rect 15945 37417 15979 37451
rect 15979 37417 15988 37451
rect 15936 37408 15988 37417
rect 16488 37408 16540 37460
rect 1768 37204 1820 37256
rect 15568 37204 15620 37256
rect 15936 37204 15988 37256
rect 16028 37247 16080 37256
rect 16028 37213 16037 37247
rect 16037 37213 16071 37247
rect 16071 37213 16080 37247
rect 19340 37408 19392 37460
rect 19616 37408 19668 37460
rect 20904 37451 20956 37460
rect 20904 37417 20913 37451
rect 20913 37417 20947 37451
rect 20947 37417 20956 37451
rect 20904 37408 20956 37417
rect 24952 37451 25004 37460
rect 24952 37417 24961 37451
rect 24961 37417 24995 37451
rect 24995 37417 25004 37451
rect 24952 37408 25004 37417
rect 27160 37408 27212 37460
rect 44272 37451 44324 37460
rect 44272 37417 44281 37451
rect 44281 37417 44315 37451
rect 44315 37417 44324 37451
rect 44272 37408 44324 37417
rect 16856 37315 16908 37324
rect 16856 37281 16865 37315
rect 16865 37281 16899 37315
rect 16899 37281 16908 37315
rect 16856 37272 16908 37281
rect 18972 37272 19024 37324
rect 20168 37272 20220 37324
rect 21272 37272 21324 37324
rect 25504 37340 25556 37392
rect 26976 37340 27028 37392
rect 28816 37340 28868 37392
rect 25596 37272 25648 37324
rect 16028 37204 16080 37213
rect 19248 37247 19300 37256
rect 19248 37213 19257 37247
rect 19257 37213 19291 37247
rect 19291 37213 19300 37247
rect 19248 37204 19300 37213
rect 19708 37204 19760 37256
rect 20720 37247 20772 37256
rect 20720 37213 20729 37247
rect 20729 37213 20763 37247
rect 20763 37213 20772 37247
rect 20720 37204 20772 37213
rect 23204 37247 23256 37256
rect 16764 37136 16816 37188
rect 19800 37136 19852 37188
rect 23204 37213 23213 37247
rect 23213 37213 23247 37247
rect 23247 37213 23256 37247
rect 23204 37204 23256 37213
rect 23388 37247 23440 37256
rect 23388 37213 23397 37247
rect 23397 37213 23431 37247
rect 23431 37213 23440 37247
rect 23388 37204 23440 37213
rect 27344 37247 27396 37256
rect 27344 37213 27353 37247
rect 27353 37213 27387 37247
rect 27387 37213 27396 37247
rect 27344 37204 27396 37213
rect 27896 37204 27948 37256
rect 28356 37204 28408 37256
rect 31760 37272 31812 37324
rect 45468 37272 45520 37324
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 29460 37204 29512 37256
rect 44088 37247 44140 37256
rect 44088 37213 44097 37247
rect 44097 37213 44131 37247
rect 44131 37213 44140 37247
rect 44088 37204 44140 37213
rect 44272 37204 44324 37256
rect 15844 37068 15896 37120
rect 18420 37068 18472 37120
rect 22560 37068 22612 37120
rect 24124 37136 24176 37188
rect 24216 37068 24268 37120
rect 24952 37068 25004 37120
rect 27712 37111 27764 37120
rect 27712 37077 27721 37111
rect 27721 37077 27755 37111
rect 27755 37077 27764 37111
rect 27712 37068 27764 37077
rect 29184 37068 29236 37120
rect 47676 37136 47728 37188
rect 47768 37068 47820 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 18144 36907 18196 36916
rect 18144 36873 18153 36907
rect 18153 36873 18187 36907
rect 18187 36873 18196 36907
rect 18144 36864 18196 36873
rect 22192 36864 22244 36916
rect 24124 36907 24176 36916
rect 24124 36873 24133 36907
rect 24133 36873 24167 36907
rect 24167 36873 24176 36907
rect 24124 36864 24176 36873
rect 27068 36907 27120 36916
rect 27068 36873 27077 36907
rect 27077 36873 27111 36907
rect 27111 36873 27120 36907
rect 27068 36864 27120 36873
rect 27712 36864 27764 36916
rect 47676 36907 47728 36916
rect 47676 36873 47685 36907
rect 47685 36873 47719 36907
rect 47719 36873 47728 36907
rect 47676 36864 47728 36873
rect 19432 36796 19484 36848
rect 23204 36796 23256 36848
rect 23756 36839 23808 36848
rect 23756 36805 23765 36839
rect 23765 36805 23799 36839
rect 23799 36805 23808 36839
rect 23756 36796 23808 36805
rect 25044 36796 25096 36848
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 13912 36703 13964 36712
rect 13912 36669 13921 36703
rect 13921 36669 13955 36703
rect 13955 36669 13964 36703
rect 13912 36660 13964 36669
rect 15660 36660 15712 36712
rect 18420 36728 18472 36780
rect 22836 36771 22888 36780
rect 22836 36737 22845 36771
rect 22845 36737 22879 36771
rect 22879 36737 22888 36771
rect 22836 36728 22888 36737
rect 23020 36771 23072 36780
rect 23020 36737 23029 36771
rect 23029 36737 23063 36771
rect 23063 36737 23072 36771
rect 23020 36728 23072 36737
rect 24124 36728 24176 36780
rect 24952 36771 25004 36780
rect 24952 36737 24961 36771
rect 24961 36737 24995 36771
rect 24995 36737 25004 36771
rect 24952 36728 25004 36737
rect 18144 36660 18196 36712
rect 19340 36660 19392 36712
rect 24860 36660 24912 36712
rect 18052 36592 18104 36644
rect 19248 36592 19300 36644
rect 20720 36592 20772 36644
rect 29000 36796 29052 36848
rect 29184 36796 29236 36848
rect 44088 36796 44140 36848
rect 47032 36796 47084 36848
rect 26792 36728 26844 36780
rect 27620 36728 27672 36780
rect 47216 36728 47268 36780
rect 27896 36660 27948 36712
rect 29276 36660 29328 36712
rect 47492 36660 47544 36712
rect 47676 36660 47728 36712
rect 15936 36524 15988 36576
rect 16212 36524 16264 36576
rect 22560 36524 22612 36576
rect 23296 36524 23348 36576
rect 23388 36524 23440 36576
rect 25228 36524 25280 36576
rect 25688 36524 25740 36576
rect 28816 36524 28868 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 15660 36363 15712 36372
rect 15660 36329 15669 36363
rect 15669 36329 15703 36363
rect 15703 36329 15712 36363
rect 15660 36320 15712 36329
rect 22836 36363 22888 36372
rect 22836 36329 22845 36363
rect 22845 36329 22879 36363
rect 22879 36329 22888 36363
rect 22836 36320 22888 36329
rect 25044 36363 25096 36372
rect 25044 36329 25053 36363
rect 25053 36329 25087 36363
rect 25087 36329 25096 36363
rect 25044 36320 25096 36329
rect 25504 36363 25556 36372
rect 25504 36329 25513 36363
rect 25513 36329 25547 36363
rect 25547 36329 25556 36363
rect 25504 36320 25556 36329
rect 27988 36320 28040 36372
rect 14924 36227 14976 36236
rect 14924 36193 14933 36227
rect 14933 36193 14967 36227
rect 14967 36193 14976 36227
rect 14924 36184 14976 36193
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 16212 36184 16264 36236
rect 15844 36159 15896 36168
rect 15844 36125 15853 36159
rect 15853 36125 15887 36159
rect 15887 36125 15896 36159
rect 15844 36116 15896 36125
rect 16120 36159 16172 36168
rect 16120 36125 16129 36159
rect 16129 36125 16163 36159
rect 16163 36125 16172 36159
rect 16120 36116 16172 36125
rect 20168 36116 20220 36168
rect 22560 36116 22612 36168
rect 23572 36184 23624 36236
rect 26884 36252 26936 36304
rect 25964 36227 26016 36236
rect 23848 36116 23900 36168
rect 25504 36116 25556 36168
rect 25688 36159 25740 36168
rect 25688 36125 25697 36159
rect 25697 36125 25731 36159
rect 25731 36125 25740 36159
rect 25688 36116 25740 36125
rect 25964 36193 25973 36227
rect 25973 36193 26007 36227
rect 26007 36193 26016 36227
rect 25964 36184 26016 36193
rect 25872 36116 25924 36168
rect 26976 36159 27028 36168
rect 13912 36048 13964 36100
rect 16764 36048 16816 36100
rect 22192 36091 22244 36100
rect 22192 36057 22201 36091
rect 22201 36057 22235 36091
rect 22235 36057 22244 36091
rect 22192 36048 22244 36057
rect 23112 36091 23164 36100
rect 23112 36057 23121 36091
rect 23121 36057 23155 36091
rect 23155 36057 23164 36091
rect 23112 36048 23164 36057
rect 23296 36091 23348 36100
rect 23296 36057 23331 36091
rect 23331 36057 23348 36091
rect 23296 36048 23348 36057
rect 24768 36048 24820 36100
rect 26976 36125 26985 36159
rect 26985 36125 27019 36159
rect 27019 36125 27028 36159
rect 26976 36116 27028 36125
rect 27712 36116 27764 36168
rect 28816 36184 28868 36236
rect 26700 36048 26752 36100
rect 26884 36048 26936 36100
rect 28264 36159 28316 36168
rect 28264 36125 28273 36159
rect 28273 36125 28307 36159
rect 28307 36125 28316 36159
rect 28264 36116 28316 36125
rect 15200 35980 15252 36032
rect 16120 35980 16172 36032
rect 20904 35980 20956 36032
rect 22376 36023 22428 36032
rect 22376 35989 22385 36023
rect 22385 35989 22419 36023
rect 22419 35989 22428 36023
rect 22376 35980 22428 35989
rect 26240 35980 26292 36032
rect 28540 35980 28592 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 16764 35708 16816 35760
rect 20812 35776 20864 35828
rect 23388 35819 23440 35828
rect 23388 35785 23397 35819
rect 23397 35785 23431 35819
rect 23431 35785 23440 35819
rect 23388 35776 23440 35785
rect 24124 35819 24176 35828
rect 24124 35785 24133 35819
rect 24133 35785 24167 35819
rect 24167 35785 24176 35819
rect 24124 35776 24176 35785
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 14188 35504 14240 35556
rect 18512 35640 18564 35692
rect 22192 35708 22244 35760
rect 23572 35708 23624 35760
rect 26884 35776 26936 35828
rect 27344 35819 27396 35828
rect 27344 35785 27353 35819
rect 27353 35785 27387 35819
rect 27387 35785 27396 35819
rect 27344 35776 27396 35785
rect 29000 35776 29052 35828
rect 29276 35819 29328 35828
rect 29276 35785 29285 35819
rect 29285 35785 29319 35819
rect 29319 35785 29328 35819
rect 29276 35776 29328 35785
rect 29368 35776 29420 35828
rect 47860 35776 47912 35828
rect 20904 35640 20956 35692
rect 22284 35683 22336 35692
rect 22284 35649 22293 35683
rect 22293 35649 22327 35683
rect 22327 35649 22336 35683
rect 22284 35640 22336 35649
rect 22744 35640 22796 35692
rect 23480 35640 23532 35692
rect 29644 35708 29696 35760
rect 24768 35683 24820 35692
rect 18144 35615 18196 35624
rect 18144 35581 18153 35615
rect 18153 35581 18187 35615
rect 18187 35581 18196 35615
rect 18144 35572 18196 35581
rect 18420 35572 18472 35624
rect 19800 35615 19852 35624
rect 19800 35581 19809 35615
rect 19809 35581 19843 35615
rect 19843 35581 19852 35615
rect 19800 35572 19852 35581
rect 20260 35572 20312 35624
rect 18052 35504 18104 35556
rect 2044 35436 2096 35488
rect 17500 35436 17552 35488
rect 17684 35436 17736 35488
rect 24768 35649 24777 35683
rect 24777 35649 24811 35683
rect 24811 35649 24820 35683
rect 24768 35640 24820 35649
rect 25504 35683 25556 35692
rect 25504 35649 25513 35683
rect 25513 35649 25547 35683
rect 25547 35649 25556 35683
rect 25504 35640 25556 35649
rect 26240 35683 26292 35692
rect 26240 35649 26249 35683
rect 26249 35649 26283 35683
rect 26283 35649 26292 35683
rect 26240 35640 26292 35649
rect 26424 35683 26476 35692
rect 26424 35649 26433 35683
rect 26433 35649 26467 35683
rect 26467 35649 26476 35683
rect 26424 35640 26476 35649
rect 28540 35683 28592 35692
rect 28540 35649 28549 35683
rect 28549 35649 28583 35683
rect 28583 35649 28592 35683
rect 28540 35640 28592 35649
rect 29000 35640 29052 35692
rect 29184 35640 29236 35692
rect 29920 35640 29972 35692
rect 24676 35572 24728 35624
rect 27068 35615 27120 35624
rect 26056 35504 26108 35556
rect 27068 35581 27077 35615
rect 27077 35581 27111 35615
rect 27111 35581 27120 35615
rect 27068 35572 27120 35581
rect 28816 35615 28868 35624
rect 28816 35581 28825 35615
rect 28825 35581 28859 35615
rect 28859 35581 28868 35615
rect 28816 35572 28868 35581
rect 28908 35615 28960 35624
rect 28908 35581 28917 35615
rect 28917 35581 28951 35615
rect 28951 35581 28960 35615
rect 28908 35572 28960 35581
rect 30196 35683 30248 35692
rect 30196 35649 30205 35683
rect 30205 35649 30239 35683
rect 30239 35649 30248 35683
rect 30196 35640 30248 35649
rect 21088 35436 21140 35488
rect 21272 35479 21324 35488
rect 21272 35445 21281 35479
rect 21281 35445 21315 35479
rect 21315 35445 21324 35479
rect 21272 35436 21324 35445
rect 22468 35436 22520 35488
rect 23020 35479 23072 35488
rect 23020 35445 23029 35479
rect 23029 35445 23063 35479
rect 23063 35445 23072 35479
rect 23020 35436 23072 35445
rect 24860 35479 24912 35488
rect 24860 35445 24869 35479
rect 24869 35445 24903 35479
rect 24903 35445 24912 35479
rect 24860 35436 24912 35445
rect 26240 35436 26292 35488
rect 26700 35436 26752 35488
rect 30932 35436 30984 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19800 35232 19852 35284
rect 21088 35275 21140 35284
rect 21088 35241 21097 35275
rect 21097 35241 21131 35275
rect 21131 35241 21140 35275
rect 22376 35275 22428 35284
rect 21088 35232 21140 35241
rect 18604 35164 18656 35216
rect 22376 35241 22385 35275
rect 22385 35241 22419 35275
rect 22419 35241 22428 35275
rect 22376 35232 22428 35241
rect 30012 35232 30064 35284
rect 16764 35139 16816 35148
rect 16764 35105 16773 35139
rect 16773 35105 16807 35139
rect 16807 35105 16816 35139
rect 16764 35096 16816 35105
rect 19432 35028 19484 35080
rect 21180 35139 21232 35148
rect 21180 35105 21189 35139
rect 21189 35105 21223 35139
rect 21223 35105 21232 35139
rect 21180 35096 21232 35105
rect 21456 35096 21508 35148
rect 22468 35139 22520 35148
rect 22468 35105 22477 35139
rect 22477 35105 22511 35139
rect 22511 35105 22520 35139
rect 22468 35096 22520 35105
rect 25688 35096 25740 35148
rect 26424 35096 26476 35148
rect 26976 35139 27028 35148
rect 26976 35105 26985 35139
rect 26985 35105 27019 35139
rect 27019 35105 27028 35139
rect 26976 35096 27028 35105
rect 27344 35096 27396 35148
rect 17040 35003 17092 35012
rect 17040 34969 17049 35003
rect 17049 34969 17083 35003
rect 17083 34969 17092 35003
rect 17040 34960 17092 34969
rect 17500 34960 17552 35012
rect 15016 34892 15068 34944
rect 15568 34892 15620 34944
rect 18512 34935 18564 34944
rect 18512 34901 18521 34935
rect 18521 34901 18555 34935
rect 18555 34901 18564 34935
rect 18512 34892 18564 34901
rect 19984 34960 20036 35012
rect 20720 35028 20772 35080
rect 21272 35028 21324 35080
rect 23756 35028 23808 35080
rect 24400 35071 24452 35080
rect 24400 35037 24409 35071
rect 24409 35037 24443 35071
rect 24443 35037 24452 35071
rect 24400 35028 24452 35037
rect 25780 35071 25832 35080
rect 25780 35037 25789 35071
rect 25789 35037 25823 35071
rect 25823 35037 25832 35071
rect 25780 35028 25832 35037
rect 25872 35028 25924 35080
rect 26700 35071 26752 35080
rect 22376 34960 22428 35012
rect 24124 34960 24176 35012
rect 26700 35037 26709 35071
rect 26709 35037 26743 35071
rect 26743 35037 26752 35071
rect 26700 35028 26752 35037
rect 27712 35096 27764 35148
rect 32128 35096 32180 35148
rect 48136 35071 48188 35080
rect 48136 35037 48145 35071
rect 48145 35037 48179 35071
rect 48179 35037 48188 35071
rect 48136 35028 48188 35037
rect 30748 34960 30800 35012
rect 32220 34960 32272 35012
rect 20260 34892 20312 34944
rect 20444 34892 20496 34944
rect 21180 34892 21232 34944
rect 21732 34892 21784 34944
rect 23112 34892 23164 34944
rect 26884 34892 26936 34944
rect 29920 34892 29972 34944
rect 47124 34892 47176 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 10324 34688 10376 34740
rect 15476 34620 15528 34672
rect 17040 34688 17092 34740
rect 20812 34688 20864 34740
rect 25872 34731 25924 34740
rect 18420 34663 18472 34672
rect 14188 34595 14240 34604
rect 14188 34561 14197 34595
rect 14197 34561 14231 34595
rect 14231 34561 14240 34595
rect 14188 34552 14240 34561
rect 15016 34595 15068 34604
rect 15016 34561 15025 34595
rect 15025 34561 15059 34595
rect 15059 34561 15068 34595
rect 15016 34552 15068 34561
rect 15108 34595 15160 34604
rect 15108 34561 15117 34595
rect 15117 34561 15151 34595
rect 15151 34561 15160 34595
rect 15108 34552 15160 34561
rect 16028 34552 16080 34604
rect 17224 34595 17276 34604
rect 17224 34561 17233 34595
rect 17233 34561 17267 34595
rect 17267 34561 17276 34595
rect 17224 34552 17276 34561
rect 17316 34552 17368 34604
rect 18420 34629 18429 34663
rect 18429 34629 18463 34663
rect 18463 34629 18472 34663
rect 18420 34620 18472 34629
rect 19432 34620 19484 34672
rect 20720 34620 20772 34672
rect 20904 34620 20956 34672
rect 25872 34697 25881 34731
rect 25881 34697 25915 34731
rect 25915 34697 25924 34731
rect 25872 34688 25924 34697
rect 29368 34688 29420 34740
rect 30748 34731 30800 34740
rect 30748 34697 30757 34731
rect 30757 34697 30791 34731
rect 30791 34697 30800 34731
rect 30748 34688 30800 34697
rect 32220 34731 32272 34740
rect 32220 34697 32229 34731
rect 32229 34697 32263 34731
rect 32263 34697 32272 34731
rect 32220 34688 32272 34697
rect 17776 34595 17828 34604
rect 17776 34561 17785 34595
rect 17785 34561 17819 34595
rect 17819 34561 17828 34595
rect 17776 34552 17828 34561
rect 18512 34552 18564 34604
rect 15292 34527 15344 34536
rect 15292 34493 15301 34527
rect 15301 34493 15335 34527
rect 15335 34493 15344 34527
rect 15292 34484 15344 34493
rect 20260 34552 20312 34604
rect 20812 34552 20864 34604
rect 21180 34552 21232 34604
rect 17592 34416 17644 34468
rect 20996 34484 21048 34536
rect 21088 34484 21140 34536
rect 22284 34552 22336 34604
rect 26056 34595 26108 34604
rect 26056 34561 26065 34595
rect 26065 34561 26099 34595
rect 26099 34561 26108 34595
rect 26056 34552 26108 34561
rect 26976 34620 27028 34672
rect 30840 34620 30892 34672
rect 26240 34552 26292 34604
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 29920 34552 29972 34561
rect 30104 34552 30156 34604
rect 30932 34595 30984 34604
rect 30932 34561 30941 34595
rect 30941 34561 30975 34595
rect 30975 34561 30984 34595
rect 30932 34552 30984 34561
rect 23664 34484 23716 34536
rect 24768 34484 24820 34536
rect 29828 34527 29880 34536
rect 14556 34348 14608 34400
rect 18788 34391 18840 34400
rect 18788 34357 18797 34391
rect 18797 34357 18831 34391
rect 18831 34357 18840 34391
rect 18788 34348 18840 34357
rect 19432 34348 19484 34400
rect 19984 34348 20036 34400
rect 21456 34416 21508 34468
rect 20720 34348 20772 34400
rect 20996 34348 21048 34400
rect 21548 34348 21600 34400
rect 23480 34348 23532 34400
rect 29828 34493 29837 34527
rect 29837 34493 29871 34527
rect 29871 34493 29880 34527
rect 29828 34484 29880 34493
rect 25044 34416 25096 34468
rect 29184 34416 29236 34468
rect 32864 34552 32916 34604
rect 48136 34595 48188 34604
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 25136 34348 25188 34400
rect 26424 34348 26476 34400
rect 47860 34348 47912 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 15016 34144 15068 34196
rect 13912 34008 13964 34060
rect 14924 34008 14976 34060
rect 17040 34144 17092 34196
rect 17592 34187 17644 34196
rect 17592 34153 17601 34187
rect 17601 34153 17635 34187
rect 17635 34153 17644 34187
rect 17592 34144 17644 34153
rect 17776 34144 17828 34196
rect 25044 34144 25096 34196
rect 17224 34076 17276 34128
rect 26976 34144 27028 34196
rect 27344 34144 27396 34196
rect 28816 34076 28868 34128
rect 1584 33983 1636 33992
rect 1584 33949 1593 33983
rect 1593 33949 1627 33983
rect 1627 33949 1636 33983
rect 1584 33940 1636 33949
rect 15476 33940 15528 33992
rect 21732 34008 21784 34060
rect 17684 33983 17736 33992
rect 14372 33915 14424 33924
rect 14372 33881 14381 33915
rect 14381 33881 14415 33915
rect 14415 33881 14424 33915
rect 14372 33872 14424 33881
rect 17684 33949 17693 33983
rect 17693 33949 17727 33983
rect 17727 33949 17736 33983
rect 17684 33940 17736 33949
rect 20536 33940 20588 33992
rect 20720 33940 20772 33992
rect 1952 33804 2004 33856
rect 13912 33804 13964 33856
rect 18512 33872 18564 33924
rect 23480 33940 23532 33992
rect 25412 34008 25464 34060
rect 24400 33983 24452 33992
rect 24400 33949 24409 33983
rect 24409 33949 24443 33983
rect 24443 33949 24452 33983
rect 24400 33940 24452 33949
rect 27620 34008 27672 34060
rect 22192 33872 22244 33924
rect 27712 33940 27764 33992
rect 25780 33915 25832 33924
rect 25780 33881 25789 33915
rect 25789 33881 25823 33915
rect 25823 33881 25832 33915
rect 25780 33872 25832 33881
rect 26332 33872 26384 33924
rect 15844 33847 15896 33856
rect 15844 33813 15853 33847
rect 15853 33813 15887 33847
rect 15887 33813 15896 33847
rect 15844 33804 15896 33813
rect 16396 33847 16448 33856
rect 16396 33813 16405 33847
rect 16405 33813 16439 33847
rect 16439 33813 16448 33847
rect 16396 33804 16448 33813
rect 22468 33804 22520 33856
rect 23756 33847 23808 33856
rect 23756 33813 23765 33847
rect 23765 33813 23799 33847
rect 23799 33813 23808 33847
rect 23756 33804 23808 33813
rect 24584 33847 24636 33856
rect 24584 33813 24593 33847
rect 24593 33813 24627 33847
rect 24627 33813 24636 33847
rect 30104 33872 30156 33924
rect 31760 33940 31812 33992
rect 30840 33872 30892 33924
rect 47952 33915 48004 33924
rect 47952 33881 47961 33915
rect 47961 33881 47995 33915
rect 47995 33881 48004 33915
rect 47952 33872 48004 33881
rect 27988 33847 28040 33856
rect 24584 33804 24636 33813
rect 27988 33813 27997 33847
rect 27997 33813 28031 33847
rect 28031 33813 28040 33847
rect 27988 33804 28040 33813
rect 29368 33804 29420 33856
rect 31116 33847 31168 33856
rect 31116 33813 31125 33847
rect 31125 33813 31159 33847
rect 31159 33813 31168 33847
rect 31116 33804 31168 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 13912 33643 13964 33652
rect 13912 33609 13921 33643
rect 13921 33609 13955 33643
rect 13955 33609 13964 33643
rect 13912 33600 13964 33609
rect 14372 33643 14424 33652
rect 14372 33609 14381 33643
rect 14381 33609 14415 33643
rect 14415 33609 14424 33643
rect 14372 33600 14424 33609
rect 15844 33600 15896 33652
rect 14372 33464 14424 33516
rect 14556 33507 14608 33516
rect 14556 33473 14565 33507
rect 14565 33473 14599 33507
rect 14599 33473 14608 33507
rect 14556 33464 14608 33473
rect 16396 33532 16448 33584
rect 15200 33464 15252 33516
rect 16856 33507 16908 33516
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 17868 33507 17920 33516
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 1860 33396 1912 33448
rect 13912 33439 13964 33448
rect 13912 33405 13921 33439
rect 13921 33405 13955 33439
rect 13955 33405 13964 33439
rect 13912 33396 13964 33405
rect 14924 33396 14976 33448
rect 16212 33396 16264 33448
rect 16396 33396 16448 33448
rect 16488 33396 16540 33448
rect 17868 33473 17877 33507
rect 17877 33473 17911 33507
rect 17911 33473 17920 33507
rect 17868 33464 17920 33473
rect 20444 33600 20496 33652
rect 20536 33600 20588 33652
rect 24308 33600 24360 33652
rect 25412 33600 25464 33652
rect 26148 33600 26200 33652
rect 26332 33643 26384 33652
rect 26332 33609 26341 33643
rect 26341 33609 26375 33643
rect 26375 33609 26384 33643
rect 26332 33600 26384 33609
rect 27620 33643 27672 33652
rect 27620 33609 27629 33643
rect 27629 33609 27663 33643
rect 27663 33609 27672 33643
rect 27620 33600 27672 33609
rect 28816 33643 28868 33652
rect 28816 33609 28825 33643
rect 28825 33609 28859 33643
rect 28859 33609 28868 33643
rect 28816 33600 28868 33609
rect 22008 33532 22060 33584
rect 22468 33575 22520 33584
rect 22468 33541 22477 33575
rect 22477 33541 22511 33575
rect 22511 33541 22520 33575
rect 22468 33532 22520 33541
rect 23756 33532 23808 33584
rect 22192 33507 22244 33516
rect 22192 33473 22201 33507
rect 22201 33473 22235 33507
rect 22235 33473 22244 33507
rect 22192 33464 22244 33473
rect 27344 33532 27396 33584
rect 26148 33464 26200 33516
rect 26976 33464 27028 33516
rect 27804 33464 27856 33516
rect 29368 33507 29420 33516
rect 15016 33260 15068 33312
rect 17040 33303 17092 33312
rect 17040 33269 17049 33303
rect 17049 33269 17083 33303
rect 17083 33269 17092 33303
rect 17040 33260 17092 33269
rect 17132 33260 17184 33312
rect 18788 33396 18840 33448
rect 29368 33473 29377 33507
rect 29377 33473 29411 33507
rect 29411 33473 29420 33507
rect 29368 33464 29420 33473
rect 29828 33532 29880 33584
rect 30012 33532 30064 33584
rect 29736 33464 29788 33516
rect 25320 33328 25372 33380
rect 25596 33328 25648 33380
rect 29552 33328 29604 33380
rect 33140 33532 33192 33584
rect 31116 33464 31168 33516
rect 32128 33507 32180 33516
rect 32128 33473 32137 33507
rect 32137 33473 32171 33507
rect 32171 33473 32180 33507
rect 32128 33464 32180 33473
rect 30840 33439 30892 33448
rect 30840 33405 30849 33439
rect 30849 33405 30883 33439
rect 30883 33405 30892 33439
rect 30840 33396 30892 33405
rect 32404 33439 32456 33448
rect 32404 33405 32413 33439
rect 32413 33405 32447 33439
rect 32447 33405 32456 33439
rect 32404 33396 32456 33405
rect 48228 33464 48280 33516
rect 20904 33260 20956 33312
rect 23940 33303 23992 33312
rect 23940 33269 23949 33303
rect 23949 33269 23983 33303
rect 23983 33269 23992 33303
rect 23940 33260 23992 33269
rect 25412 33260 25464 33312
rect 29184 33260 29236 33312
rect 31484 33260 31536 33312
rect 31760 33260 31812 33312
rect 47216 33260 47268 33312
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1952 33099 2004 33108
rect 1952 33065 1961 33099
rect 1961 33065 1995 33099
rect 1995 33065 2004 33099
rect 1952 33056 2004 33065
rect 14372 33056 14424 33108
rect 14924 32988 14976 33040
rect 17868 33056 17920 33108
rect 17224 32988 17276 33040
rect 17316 32988 17368 33040
rect 20996 33056 21048 33108
rect 22100 33056 22152 33108
rect 23664 33031 23716 33040
rect 23664 32997 23673 33031
rect 23673 32997 23707 33031
rect 23707 32997 23716 33031
rect 23664 32988 23716 32997
rect 1952 32852 2004 32904
rect 13912 32920 13964 32972
rect 15108 32920 15160 32972
rect 14464 32895 14516 32904
rect 14464 32861 14473 32895
rect 14473 32861 14507 32895
rect 14507 32861 14516 32895
rect 14464 32852 14516 32861
rect 15016 32852 15068 32904
rect 15476 32895 15528 32904
rect 15476 32861 15485 32895
rect 15485 32861 15519 32895
rect 15519 32861 15528 32895
rect 15476 32852 15528 32861
rect 15844 32852 15896 32904
rect 16396 32895 16448 32904
rect 16396 32861 16405 32895
rect 16405 32861 16439 32895
rect 16439 32861 16448 32895
rect 16396 32852 16448 32861
rect 17132 32895 17184 32904
rect 17132 32861 17141 32895
rect 17141 32861 17175 32895
rect 17175 32861 17184 32895
rect 17132 32852 17184 32861
rect 17316 32895 17368 32904
rect 17316 32861 17325 32895
rect 17325 32861 17359 32895
rect 17359 32861 17368 32895
rect 17316 32852 17368 32861
rect 16212 32827 16264 32836
rect 16212 32793 16221 32827
rect 16221 32793 16255 32827
rect 16255 32793 16264 32827
rect 16212 32784 16264 32793
rect 2228 32716 2280 32768
rect 16856 32716 16908 32768
rect 17316 32716 17368 32768
rect 17500 32895 17552 32904
rect 17500 32861 17509 32895
rect 17509 32861 17543 32895
rect 17543 32861 17552 32895
rect 17500 32852 17552 32861
rect 17776 32852 17828 32904
rect 18512 32895 18564 32904
rect 18512 32861 18521 32895
rect 18521 32861 18555 32895
rect 18555 32861 18564 32895
rect 18512 32852 18564 32861
rect 19984 32895 20036 32904
rect 19984 32861 19993 32895
rect 19993 32861 20027 32895
rect 20027 32861 20036 32895
rect 19984 32852 20036 32861
rect 22192 32895 22244 32904
rect 22192 32861 22201 32895
rect 22201 32861 22235 32895
rect 22235 32861 22244 32895
rect 22192 32852 22244 32861
rect 23480 32920 23532 32972
rect 23940 32852 23992 32904
rect 29276 33056 29328 33108
rect 26424 32988 26476 33040
rect 31944 32988 31996 33040
rect 29828 32920 29880 32972
rect 31760 32963 31812 32972
rect 31760 32929 31769 32963
rect 31769 32929 31803 32963
rect 31803 32929 31812 32963
rect 31760 32920 31812 32929
rect 32404 33056 32456 33108
rect 33140 33056 33192 33108
rect 47124 32963 47176 32972
rect 47124 32929 47133 32963
rect 47133 32929 47167 32963
rect 47167 32929 47176 32963
rect 47124 32920 47176 32929
rect 47676 32963 47728 32972
rect 47676 32929 47685 32963
rect 47685 32929 47719 32963
rect 47719 32929 47728 32963
rect 47676 32920 47728 32929
rect 29736 32852 29788 32904
rect 31484 32895 31536 32904
rect 31484 32861 31493 32895
rect 31493 32861 31527 32895
rect 31527 32861 31536 32895
rect 31484 32852 31536 32861
rect 20260 32827 20312 32836
rect 20260 32793 20269 32827
rect 20269 32793 20303 32827
rect 20303 32793 20312 32827
rect 20260 32784 20312 32793
rect 24768 32827 24820 32836
rect 24768 32793 24777 32827
rect 24777 32793 24811 32827
rect 24811 32793 24820 32827
rect 24768 32784 24820 32793
rect 27804 32784 27856 32836
rect 31576 32784 31628 32836
rect 31852 32895 31904 32904
rect 31852 32861 31861 32895
rect 31861 32861 31895 32895
rect 31895 32861 31904 32895
rect 31852 32852 31904 32861
rect 32036 32895 32088 32904
rect 32036 32861 32045 32895
rect 32045 32861 32079 32895
rect 32079 32861 32088 32895
rect 32864 32895 32916 32904
rect 32036 32852 32088 32861
rect 32864 32861 32873 32895
rect 32873 32861 32907 32895
rect 32907 32861 32916 32895
rect 32864 32852 32916 32861
rect 46296 32852 46348 32904
rect 47216 32827 47268 32836
rect 47216 32793 47225 32827
rect 47225 32793 47259 32827
rect 47259 32793 47268 32827
rect 47216 32784 47268 32793
rect 17776 32716 17828 32768
rect 18512 32716 18564 32768
rect 21088 32716 21140 32768
rect 21824 32716 21876 32768
rect 27988 32716 28040 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 15476 32512 15528 32564
rect 2228 32487 2280 32496
rect 2228 32453 2237 32487
rect 2237 32453 2271 32487
rect 2271 32453 2280 32487
rect 2228 32444 2280 32453
rect 16396 32444 16448 32496
rect 17316 32512 17368 32564
rect 20260 32512 20312 32564
rect 24216 32555 24268 32564
rect 24216 32521 24241 32555
rect 24241 32521 24268 32555
rect 24400 32555 24452 32564
rect 24216 32512 24268 32521
rect 24400 32521 24409 32555
rect 24409 32521 24443 32555
rect 24443 32521 24452 32555
rect 24400 32512 24452 32521
rect 27620 32512 27672 32564
rect 29552 32555 29604 32564
rect 29552 32521 29561 32555
rect 29561 32521 29595 32555
rect 29595 32521 29604 32555
rect 29552 32512 29604 32521
rect 31944 32512 31996 32564
rect 17500 32444 17552 32496
rect 17776 32487 17828 32496
rect 17776 32453 17785 32487
rect 17785 32453 17819 32487
rect 17819 32453 17828 32487
rect 17776 32444 17828 32453
rect 18512 32444 18564 32496
rect 20812 32444 20864 32496
rect 20996 32444 21048 32496
rect 2044 32419 2096 32428
rect 2044 32385 2053 32419
rect 2053 32385 2087 32419
rect 2087 32385 2096 32419
rect 2044 32376 2096 32385
rect 16212 32376 16264 32428
rect 4712 32308 4764 32360
rect 16580 32308 16632 32360
rect 20352 32376 20404 32428
rect 21088 32419 21140 32428
rect 1400 32172 1452 32224
rect 19708 32308 19760 32360
rect 21088 32385 21097 32419
rect 21097 32385 21131 32419
rect 21131 32385 21140 32419
rect 21088 32376 21140 32385
rect 17868 32172 17920 32224
rect 21824 32444 21876 32496
rect 23112 32444 23164 32496
rect 25412 32444 25464 32496
rect 24952 32419 25004 32428
rect 24952 32385 24961 32419
rect 24961 32385 24995 32419
rect 24995 32385 25004 32419
rect 24952 32376 25004 32385
rect 26056 32376 26108 32428
rect 26700 32376 26752 32428
rect 28264 32444 28316 32496
rect 29920 32444 29972 32496
rect 29828 32376 29880 32428
rect 32864 32444 32916 32496
rect 32128 32419 32180 32428
rect 32128 32385 32137 32419
rect 32137 32385 32171 32419
rect 32171 32385 32180 32419
rect 32128 32376 32180 32385
rect 46664 32376 46716 32428
rect 47584 32376 47636 32428
rect 47952 32419 48004 32428
rect 47952 32385 47961 32419
rect 47961 32385 47995 32419
rect 47995 32385 48004 32419
rect 47952 32376 48004 32385
rect 25688 32351 25740 32360
rect 25688 32317 25697 32351
rect 25697 32317 25731 32351
rect 25731 32317 25740 32351
rect 25688 32308 25740 32317
rect 26792 32308 26844 32360
rect 28724 32351 28776 32360
rect 28724 32317 28733 32351
rect 28733 32317 28767 32351
rect 28767 32317 28776 32351
rect 28724 32308 28776 32317
rect 32404 32351 32456 32360
rect 32404 32317 32413 32351
rect 32413 32317 32447 32351
rect 32447 32317 32456 32351
rect 32404 32308 32456 32317
rect 20996 32240 21048 32292
rect 24124 32172 24176 32224
rect 24952 32240 25004 32292
rect 25136 32283 25188 32292
rect 25136 32249 25145 32283
rect 25145 32249 25179 32283
rect 25179 32249 25188 32283
rect 25136 32240 25188 32249
rect 28356 32240 28408 32292
rect 29184 32240 29236 32292
rect 25780 32172 25832 32224
rect 26240 32172 26292 32224
rect 27712 32172 27764 32224
rect 28540 32172 28592 32224
rect 30104 32215 30156 32224
rect 30104 32181 30113 32215
rect 30113 32181 30147 32215
rect 30147 32181 30156 32215
rect 30104 32172 30156 32181
rect 30380 32215 30432 32224
rect 30380 32181 30389 32215
rect 30389 32181 30423 32215
rect 30423 32181 30432 32215
rect 30380 32172 30432 32181
rect 31760 32172 31812 32224
rect 46480 32172 46532 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 15200 31968 15252 32020
rect 17500 31900 17552 31952
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 14464 31832 14516 31884
rect 14556 31832 14608 31884
rect 16856 31832 16908 31884
rect 15568 31764 15620 31816
rect 16488 31764 16540 31816
rect 16948 31764 17000 31816
rect 17224 31807 17276 31816
rect 17224 31773 17233 31807
rect 17233 31773 17267 31807
rect 17267 31773 17276 31807
rect 17224 31764 17276 31773
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 14372 31696 14424 31748
rect 17868 31968 17920 32020
rect 19984 31968 20036 32020
rect 17684 31900 17736 31952
rect 18420 31832 18472 31884
rect 17960 31764 18012 31816
rect 19708 31764 19760 31816
rect 20904 31900 20956 31952
rect 20996 31943 21048 31952
rect 20996 31909 21005 31943
rect 21005 31909 21039 31943
rect 21039 31909 21048 31943
rect 20996 31900 21048 31909
rect 20812 31764 20864 31816
rect 23480 32011 23532 32020
rect 23480 31977 23489 32011
rect 23489 31977 23523 32011
rect 23523 31977 23532 32011
rect 23480 31968 23532 31977
rect 24860 31968 24912 32020
rect 24952 31968 25004 32020
rect 26792 32011 26844 32020
rect 26792 31977 26801 32011
rect 26801 31977 26835 32011
rect 26835 31977 26844 32011
rect 26792 31968 26844 31977
rect 23572 31900 23624 31952
rect 24216 31900 24268 31952
rect 24400 31900 24452 31952
rect 25504 31832 25556 31884
rect 26148 31832 26200 31884
rect 27252 31875 27304 31884
rect 27252 31841 27261 31875
rect 27261 31841 27295 31875
rect 27295 31841 27304 31875
rect 27252 31832 27304 31841
rect 20904 31696 20956 31748
rect 23112 31739 23164 31748
rect 23112 31705 23121 31739
rect 23121 31705 23155 31739
rect 23155 31705 23164 31739
rect 23112 31696 23164 31705
rect 27344 31807 27396 31816
rect 24860 31696 24912 31748
rect 20168 31628 20220 31680
rect 22192 31628 22244 31680
rect 22560 31628 22612 31680
rect 24952 31628 25004 31680
rect 25136 31671 25188 31680
rect 25136 31637 25145 31671
rect 25145 31637 25179 31671
rect 25179 31637 25188 31671
rect 25136 31628 25188 31637
rect 25412 31628 25464 31680
rect 27344 31773 27353 31807
rect 27353 31773 27387 31807
rect 27387 31773 27396 31807
rect 27344 31764 27396 31773
rect 27528 31764 27580 31816
rect 27988 31807 28040 31816
rect 27988 31773 27997 31807
rect 27997 31773 28031 31807
rect 28031 31773 28040 31807
rect 27988 31764 28040 31773
rect 28356 31900 28408 31952
rect 29184 31968 29236 32020
rect 30288 32011 30340 32020
rect 30288 31977 30297 32011
rect 30297 31977 30331 32011
rect 30331 31977 30340 32011
rect 30288 31968 30340 31977
rect 32404 31968 32456 32020
rect 32864 32011 32916 32020
rect 32864 31977 32873 32011
rect 32873 31977 32907 32011
rect 32907 31977 32916 32011
rect 32864 31968 32916 31977
rect 28540 31832 28592 31884
rect 28724 31832 28776 31884
rect 28816 31807 28868 31816
rect 28816 31773 28825 31807
rect 28825 31773 28859 31807
rect 28859 31773 28868 31807
rect 28816 31764 28868 31773
rect 29828 31764 29880 31816
rect 30012 31807 30064 31816
rect 30012 31773 30021 31807
rect 30021 31773 30055 31807
rect 30055 31773 30064 31807
rect 30012 31764 30064 31773
rect 31760 31875 31812 31884
rect 31760 31841 31769 31875
rect 31769 31841 31803 31875
rect 31803 31841 31812 31875
rect 31760 31832 31812 31841
rect 40408 31900 40460 31952
rect 46296 31875 46348 31884
rect 46296 31841 46305 31875
rect 46305 31841 46339 31875
rect 46339 31841 46348 31875
rect 46296 31832 46348 31841
rect 46480 31875 46532 31884
rect 46480 31841 46489 31875
rect 46489 31841 46523 31875
rect 46523 31841 46532 31875
rect 46480 31832 46532 31841
rect 48136 31875 48188 31884
rect 48136 31841 48145 31875
rect 48145 31841 48179 31875
rect 48179 31841 48188 31875
rect 48136 31832 48188 31841
rect 31576 31764 31628 31816
rect 32036 31807 32088 31816
rect 32036 31773 32045 31807
rect 32045 31773 32079 31807
rect 32079 31773 32088 31807
rect 32036 31764 32088 31773
rect 32128 31764 32180 31816
rect 32772 31807 32824 31816
rect 32772 31773 32781 31807
rect 32781 31773 32815 31807
rect 32815 31773 32824 31807
rect 32772 31764 32824 31773
rect 28632 31696 28684 31748
rect 30380 31696 30432 31748
rect 27528 31628 27580 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 15568 31467 15620 31476
rect 15568 31433 15577 31467
rect 15577 31433 15611 31467
rect 15611 31433 15620 31467
rect 15568 31424 15620 31433
rect 24124 31424 24176 31476
rect 1952 31356 2004 31408
rect 4712 31399 4764 31408
rect 4712 31365 4721 31399
rect 4721 31365 4755 31399
rect 4755 31365 4764 31399
rect 4712 31356 4764 31365
rect 15660 31356 15712 31408
rect 20720 31399 20772 31408
rect 20720 31365 20729 31399
rect 20729 31365 20763 31399
rect 20763 31365 20772 31399
rect 20720 31356 20772 31365
rect 28632 31424 28684 31476
rect 2320 31288 2372 31340
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 18328 31288 18380 31340
rect 20168 31288 20220 31340
rect 20996 31288 21048 31340
rect 23572 31331 23624 31340
rect 23572 31297 23581 31331
rect 23581 31297 23615 31331
rect 23615 31297 23624 31331
rect 23572 31288 23624 31297
rect 24584 31331 24636 31340
rect 24584 31297 24593 31331
rect 24593 31297 24627 31331
rect 24627 31297 24636 31331
rect 24584 31288 24636 31297
rect 25780 31331 25832 31340
rect 25780 31297 25789 31331
rect 25789 31297 25823 31331
rect 25823 31297 25832 31331
rect 25780 31288 25832 31297
rect 27436 31288 27488 31340
rect 28632 31331 28684 31340
rect 28632 31297 28641 31331
rect 28641 31297 28675 31331
rect 28675 31297 28684 31331
rect 28632 31288 28684 31297
rect 28816 31288 28868 31340
rect 30104 31424 30156 31476
rect 30380 31424 30432 31476
rect 30012 31288 30064 31340
rect 32128 31331 32180 31340
rect 2872 31263 2924 31272
rect 2872 31229 2881 31263
rect 2881 31229 2915 31263
rect 2915 31229 2924 31263
rect 2872 31220 2924 31229
rect 15108 31220 15160 31272
rect 16856 31263 16908 31272
rect 16856 31229 16865 31263
rect 16865 31229 16899 31263
rect 16899 31229 16908 31263
rect 16856 31220 16908 31229
rect 23204 31220 23256 31272
rect 29920 31263 29972 31272
rect 29920 31229 29929 31263
rect 29929 31229 29963 31263
rect 29963 31229 29972 31263
rect 29920 31220 29972 31229
rect 17040 31152 17092 31204
rect 16396 31084 16448 31136
rect 17316 31084 17368 31136
rect 18052 31127 18104 31136
rect 18052 31093 18061 31127
rect 18061 31093 18095 31127
rect 18095 31093 18104 31127
rect 18052 31084 18104 31093
rect 20168 31127 20220 31136
rect 20168 31093 20177 31127
rect 20177 31093 20211 31127
rect 20211 31093 20220 31127
rect 20168 31084 20220 31093
rect 20444 31084 20496 31136
rect 20904 31084 20956 31136
rect 23756 31152 23808 31204
rect 27988 31152 28040 31204
rect 28724 31152 28776 31204
rect 32128 31297 32137 31331
rect 32137 31297 32171 31331
rect 32171 31297 32180 31331
rect 32128 31288 32180 31297
rect 24676 31084 24728 31136
rect 25412 31084 25464 31136
rect 25688 31084 25740 31136
rect 27712 31127 27764 31136
rect 27712 31093 27721 31127
rect 27721 31093 27755 31127
rect 27755 31093 27764 31127
rect 27712 31084 27764 31093
rect 30104 31084 30156 31136
rect 32220 31127 32272 31136
rect 32220 31093 32229 31127
rect 32229 31093 32263 31127
rect 32263 31093 32272 31127
rect 32220 31084 32272 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 15108 30923 15160 30932
rect 15108 30889 15117 30923
rect 15117 30889 15151 30923
rect 15151 30889 15160 30923
rect 15108 30880 15160 30889
rect 15660 30923 15712 30932
rect 15660 30889 15669 30923
rect 15669 30889 15703 30923
rect 15703 30889 15712 30923
rect 15660 30880 15712 30889
rect 16672 30880 16724 30932
rect 17132 30880 17184 30932
rect 17316 30923 17368 30932
rect 17316 30889 17325 30923
rect 17325 30889 17359 30923
rect 17359 30889 17368 30923
rect 17316 30880 17368 30889
rect 18420 30880 18472 30932
rect 20904 30880 20956 30932
rect 24860 30880 24912 30932
rect 25412 30880 25464 30932
rect 29920 30880 29972 30932
rect 14372 30744 14424 30796
rect 14464 30719 14516 30728
rect 14464 30685 14473 30719
rect 14473 30685 14507 30719
rect 14507 30685 14516 30719
rect 14464 30676 14516 30685
rect 15016 30676 15068 30728
rect 18052 30812 18104 30864
rect 17040 30744 17092 30796
rect 17868 30744 17920 30796
rect 20536 30744 20588 30796
rect 20812 30744 20864 30796
rect 21272 30744 21324 30796
rect 16396 30608 16448 30660
rect 16304 30540 16356 30592
rect 16580 30540 16632 30592
rect 17500 30676 17552 30728
rect 18328 30719 18380 30728
rect 18328 30685 18337 30719
rect 18337 30685 18371 30719
rect 18371 30685 18380 30719
rect 18328 30676 18380 30685
rect 18788 30676 18840 30728
rect 21640 30719 21692 30728
rect 21640 30685 21649 30719
rect 21649 30685 21683 30719
rect 21683 30685 21692 30719
rect 21640 30676 21692 30685
rect 22560 30719 22612 30728
rect 22560 30685 22569 30719
rect 22569 30685 22603 30719
rect 22603 30685 22612 30719
rect 22560 30676 22612 30685
rect 24584 30812 24636 30864
rect 29644 30812 29696 30864
rect 30012 30812 30064 30864
rect 23664 30744 23716 30796
rect 29552 30744 29604 30796
rect 43076 30744 43128 30796
rect 47676 30744 47728 30796
rect 20168 30608 20220 30660
rect 20812 30540 20864 30592
rect 20996 30583 21048 30592
rect 20996 30549 21005 30583
rect 21005 30549 21039 30583
rect 21039 30549 21048 30583
rect 20996 30540 21048 30549
rect 21456 30583 21508 30592
rect 21456 30549 21465 30583
rect 21465 30549 21499 30583
rect 21499 30549 21508 30583
rect 21456 30540 21508 30549
rect 22100 30540 22152 30592
rect 22744 30540 22796 30592
rect 23204 30608 23256 30660
rect 24860 30676 24912 30728
rect 25320 30676 25372 30728
rect 27804 30719 27856 30728
rect 27804 30685 27813 30719
rect 27813 30685 27847 30719
rect 27847 30685 27856 30719
rect 27804 30676 27856 30685
rect 28724 30719 28776 30728
rect 28724 30685 28733 30719
rect 28733 30685 28767 30719
rect 28767 30685 28776 30719
rect 28724 30676 28776 30685
rect 23756 30583 23808 30592
rect 23756 30549 23765 30583
rect 23765 30549 23799 30583
rect 23799 30549 23808 30583
rect 23756 30540 23808 30549
rect 27068 30608 27120 30660
rect 26332 30540 26384 30592
rect 26700 30540 26752 30592
rect 29644 30540 29696 30592
rect 29828 30719 29880 30728
rect 29828 30685 29837 30719
rect 29837 30685 29871 30719
rect 29871 30685 29880 30719
rect 30012 30719 30064 30728
rect 29828 30676 29880 30685
rect 30012 30685 30021 30719
rect 30021 30685 30055 30719
rect 30055 30685 30064 30719
rect 30012 30676 30064 30685
rect 30104 30719 30156 30728
rect 30104 30685 30113 30719
rect 30113 30685 30147 30719
rect 30147 30685 30156 30719
rect 30104 30676 30156 30685
rect 32220 30676 32272 30728
rect 31116 30651 31168 30660
rect 31116 30617 31125 30651
rect 31125 30617 31159 30651
rect 31159 30617 31168 30651
rect 31116 30608 31168 30617
rect 45744 30608 45796 30660
rect 43352 30540 43404 30592
rect 48228 30540 48280 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 14464 30336 14516 30388
rect 16856 30336 16908 30388
rect 17960 30268 18012 30320
rect 20444 30336 20496 30388
rect 20536 30336 20588 30388
rect 14556 30243 14608 30252
rect 14556 30209 14565 30243
rect 14565 30209 14599 30243
rect 14599 30209 14608 30243
rect 14556 30200 14608 30209
rect 14740 30243 14792 30252
rect 14740 30209 14749 30243
rect 14749 30209 14783 30243
rect 14783 30209 14792 30243
rect 14740 30200 14792 30209
rect 16948 30175 17000 30184
rect 16948 30141 16957 30175
rect 16957 30141 16991 30175
rect 16991 30141 17000 30175
rect 16948 30132 17000 30141
rect 17040 29996 17092 30048
rect 20720 30268 20772 30320
rect 20996 30268 21048 30320
rect 20536 30200 20588 30252
rect 20812 30200 20864 30252
rect 21180 30200 21232 30252
rect 22744 30268 22796 30320
rect 24584 30268 24636 30320
rect 24400 30200 24452 30252
rect 25688 30243 25740 30252
rect 25688 30209 25697 30243
rect 25697 30209 25731 30243
rect 25731 30209 25740 30243
rect 25688 30200 25740 30209
rect 26056 30336 26108 30388
rect 26332 30379 26384 30388
rect 26332 30345 26341 30379
rect 26341 30345 26375 30379
rect 26375 30345 26384 30379
rect 26332 30336 26384 30345
rect 27712 30336 27764 30388
rect 26700 30268 26752 30320
rect 27068 30311 27120 30320
rect 27068 30277 27077 30311
rect 27077 30277 27111 30311
rect 27111 30277 27120 30311
rect 27068 30268 27120 30277
rect 25964 30243 26016 30252
rect 25964 30209 25973 30243
rect 25973 30209 26007 30243
rect 26007 30209 26016 30243
rect 25964 30200 26016 30209
rect 26056 30243 26108 30252
rect 26056 30209 26065 30243
rect 26065 30209 26099 30243
rect 26099 30209 26108 30243
rect 26056 30200 26108 30209
rect 26976 30243 27028 30252
rect 20352 30064 20404 30116
rect 20444 30064 20496 30116
rect 22836 30132 22888 30184
rect 23388 30064 23440 30116
rect 23664 29996 23716 30048
rect 23756 30039 23808 30048
rect 23756 30005 23765 30039
rect 23765 30005 23799 30039
rect 23799 30005 23808 30039
rect 25504 30064 25556 30116
rect 26976 30209 26985 30243
rect 26985 30209 27019 30243
rect 27019 30209 27028 30243
rect 26976 30200 27028 30209
rect 32128 30336 32180 30388
rect 28264 30268 28316 30320
rect 31116 30268 31168 30320
rect 29644 30243 29696 30252
rect 29644 30209 29653 30243
rect 29653 30209 29687 30243
rect 29687 30209 29696 30243
rect 29644 30200 29696 30209
rect 29920 30243 29972 30252
rect 29920 30209 29929 30243
rect 29929 30209 29963 30243
rect 29963 30209 29972 30243
rect 29920 30200 29972 30209
rect 34520 30268 34572 30320
rect 29368 30132 29420 30184
rect 29828 30132 29880 30184
rect 33140 30175 33192 30184
rect 33140 30141 33149 30175
rect 33149 30141 33183 30175
rect 33183 30141 33192 30175
rect 33140 30132 33192 30141
rect 26332 30064 26384 30116
rect 23756 29996 23808 30005
rect 29000 29996 29052 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 16948 29792 17000 29844
rect 14740 29724 14792 29776
rect 20168 29792 20220 29844
rect 21272 29792 21324 29844
rect 21456 29835 21508 29844
rect 21456 29801 21465 29835
rect 21465 29801 21499 29835
rect 21499 29801 21508 29835
rect 21456 29792 21508 29801
rect 21548 29792 21600 29844
rect 22836 29835 22888 29844
rect 22836 29801 22845 29835
rect 22845 29801 22879 29835
rect 22879 29801 22888 29835
rect 22836 29792 22888 29801
rect 16580 29656 16632 29708
rect 16304 29631 16356 29640
rect 16304 29597 16313 29631
rect 16313 29597 16347 29631
rect 16347 29597 16356 29631
rect 16304 29588 16356 29597
rect 16488 29631 16540 29640
rect 16488 29597 16502 29631
rect 16502 29597 16536 29631
rect 16536 29597 16540 29631
rect 16488 29588 16540 29597
rect 16396 29563 16448 29572
rect 16396 29529 16405 29563
rect 16405 29529 16439 29563
rect 16439 29529 16448 29563
rect 16396 29520 16448 29529
rect 17408 29588 17460 29640
rect 20720 29656 20772 29708
rect 24400 29724 24452 29776
rect 21548 29656 21600 29708
rect 21640 29656 21692 29708
rect 23756 29656 23808 29708
rect 27344 29792 27396 29844
rect 21088 29631 21140 29640
rect 21088 29597 21097 29631
rect 21097 29597 21131 29631
rect 21131 29597 21140 29631
rect 21088 29588 21140 29597
rect 19984 29520 20036 29572
rect 16856 29452 16908 29504
rect 17316 29452 17368 29504
rect 21456 29452 21508 29504
rect 22468 29631 22520 29640
rect 21732 29520 21784 29572
rect 22468 29597 22477 29631
rect 22477 29597 22511 29631
rect 22511 29597 22520 29631
rect 22468 29588 22520 29597
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 24308 29588 24360 29640
rect 24952 29588 25004 29640
rect 29368 29724 29420 29776
rect 29736 29792 29788 29844
rect 33140 29835 33192 29844
rect 33140 29801 33149 29835
rect 33149 29801 33183 29835
rect 33183 29801 33192 29835
rect 33140 29792 33192 29801
rect 30380 29724 30432 29776
rect 25320 29656 25372 29708
rect 26332 29656 26384 29708
rect 28540 29656 28592 29708
rect 29828 29631 29880 29640
rect 23388 29520 23440 29572
rect 23940 29520 23992 29572
rect 28448 29520 28500 29572
rect 28724 29520 28776 29572
rect 28816 29520 28868 29572
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 29920 29588 29972 29640
rect 30840 29631 30892 29640
rect 30840 29597 30849 29631
rect 30849 29597 30883 29631
rect 30883 29597 30892 29631
rect 30840 29588 30892 29597
rect 30932 29631 30984 29640
rect 30932 29597 30941 29631
rect 30941 29597 30975 29631
rect 30975 29597 30984 29631
rect 30932 29588 30984 29597
rect 32956 29588 33008 29640
rect 46848 29588 46900 29640
rect 48136 29631 48188 29640
rect 48136 29597 48145 29631
rect 48145 29597 48179 29631
rect 48179 29597 48188 29631
rect 48136 29588 48188 29597
rect 32772 29520 32824 29572
rect 23296 29452 23348 29504
rect 26056 29452 26108 29504
rect 30472 29495 30524 29504
rect 30472 29461 30481 29495
rect 30481 29461 30515 29495
rect 30515 29461 30524 29495
rect 30472 29452 30524 29461
rect 47032 29452 47084 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 3332 29248 3384 29300
rect 25320 29248 25372 29300
rect 26056 29248 26108 29300
rect 26884 29248 26936 29300
rect 29920 29248 29972 29300
rect 30012 29248 30064 29300
rect 30288 29291 30340 29300
rect 30288 29257 30297 29291
rect 30297 29257 30331 29291
rect 30331 29257 30340 29291
rect 30288 29248 30340 29257
rect 1676 29180 1728 29232
rect 14464 29180 14516 29232
rect 17316 29155 17368 29164
rect 17316 29121 17325 29155
rect 17325 29121 17359 29155
rect 17359 29121 17368 29155
rect 17316 29112 17368 29121
rect 17408 29155 17460 29164
rect 17408 29121 17418 29155
rect 17418 29121 17452 29155
rect 17452 29121 17460 29155
rect 17408 29112 17460 29121
rect 18144 29180 18196 29232
rect 19984 29155 20036 29164
rect 17224 29044 17276 29096
rect 16304 28976 16356 29028
rect 19984 29121 19993 29155
rect 19993 29121 20027 29155
rect 20027 29121 20036 29155
rect 19984 29112 20036 29121
rect 20260 29112 20312 29164
rect 20352 29155 20404 29164
rect 20352 29121 20361 29155
rect 20361 29121 20395 29155
rect 20395 29121 20404 29155
rect 20352 29112 20404 29121
rect 21916 29112 21968 29164
rect 23940 29112 23992 29164
rect 20444 29044 20496 29096
rect 25780 29155 25832 29164
rect 25780 29121 25789 29155
rect 25789 29121 25823 29155
rect 25823 29121 25832 29155
rect 25780 29112 25832 29121
rect 28816 29180 28868 29232
rect 28540 29155 28592 29164
rect 28540 29121 28549 29155
rect 28549 29121 28583 29155
rect 28583 29121 28592 29155
rect 28540 29112 28592 29121
rect 29460 29155 29512 29164
rect 27436 29087 27488 29096
rect 20536 28976 20588 29028
rect 27436 29053 27445 29087
rect 27445 29053 27479 29087
rect 27479 29053 27488 29087
rect 27436 29044 27488 29053
rect 27620 29087 27672 29096
rect 27620 29053 27629 29087
rect 27629 29053 27663 29087
rect 27663 29053 27672 29087
rect 27620 29044 27672 29053
rect 24492 28976 24544 29028
rect 26976 29019 27028 29028
rect 26976 28985 26985 29019
rect 26985 28985 27019 29019
rect 27019 28985 27028 29019
rect 26976 28976 27028 28985
rect 17960 28951 18012 28960
rect 17960 28917 17969 28951
rect 17969 28917 18003 28951
rect 18003 28917 18012 28951
rect 17960 28908 18012 28917
rect 25596 28951 25648 28960
rect 25596 28917 25605 28951
rect 25605 28917 25639 28951
rect 25639 28917 25648 28951
rect 25596 28908 25648 28917
rect 27804 28908 27856 28960
rect 27988 28908 28040 28960
rect 28172 28908 28224 28960
rect 29460 29121 29469 29155
rect 29469 29121 29503 29155
rect 29503 29121 29512 29155
rect 29460 29112 29512 29121
rect 29368 29044 29420 29096
rect 30012 29112 30064 29164
rect 29828 29044 29880 29096
rect 31760 29112 31812 29164
rect 30288 28976 30340 29028
rect 30380 28908 30432 28960
rect 31300 29044 31352 29096
rect 32312 29087 32364 29096
rect 32312 29053 32321 29087
rect 32321 29053 32355 29087
rect 32355 29053 32364 29087
rect 32312 29044 32364 29053
rect 32496 29087 32548 29096
rect 32496 29053 32505 29087
rect 32505 29053 32539 29087
rect 32539 29053 32548 29087
rect 32496 29044 32548 29053
rect 32772 29087 32824 29096
rect 32772 29053 32781 29087
rect 32781 29053 32815 29087
rect 32815 29053 32824 29087
rect 32772 29044 32824 29053
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 17500 28747 17552 28756
rect 17500 28713 17509 28747
rect 17509 28713 17543 28747
rect 17543 28713 17552 28747
rect 17500 28704 17552 28713
rect 7472 28636 7524 28688
rect 19800 28704 19852 28756
rect 25964 28747 26016 28756
rect 25964 28713 25973 28747
rect 25973 28713 26007 28747
rect 26007 28713 26016 28747
rect 25964 28704 26016 28713
rect 29000 28747 29052 28756
rect 19432 28636 19484 28688
rect 19524 28636 19576 28688
rect 21732 28636 21784 28688
rect 28632 28636 28684 28688
rect 29000 28713 29009 28747
rect 29009 28713 29043 28747
rect 29043 28713 29052 28747
rect 29000 28704 29052 28713
rect 30288 28704 30340 28756
rect 31300 28747 31352 28756
rect 31300 28713 31309 28747
rect 31309 28713 31343 28747
rect 31343 28713 31352 28747
rect 31300 28704 31352 28713
rect 32496 28747 32548 28756
rect 32496 28713 32505 28747
rect 32505 28713 32539 28747
rect 32539 28713 32548 28747
rect 32496 28704 32548 28713
rect 29460 28636 29512 28688
rect 19156 28568 19208 28620
rect 17224 28543 17276 28552
rect 17224 28509 17233 28543
rect 17233 28509 17267 28543
rect 17267 28509 17276 28543
rect 17224 28500 17276 28509
rect 19800 28568 19852 28620
rect 20168 28568 20220 28620
rect 22100 28568 22152 28620
rect 27988 28568 28040 28620
rect 29552 28611 29604 28620
rect 29552 28577 29561 28611
rect 29561 28577 29595 28611
rect 29595 28577 29604 28611
rect 29552 28568 29604 28577
rect 30472 28568 30524 28620
rect 18236 28432 18288 28484
rect 22652 28500 22704 28552
rect 25044 28500 25096 28552
rect 26240 28500 26292 28552
rect 27436 28500 27488 28552
rect 27804 28500 27856 28552
rect 28172 28543 28224 28552
rect 28172 28509 28181 28543
rect 28181 28509 28215 28543
rect 28215 28509 28224 28543
rect 28172 28500 28224 28509
rect 28724 28500 28776 28552
rect 32220 28500 32272 28552
rect 46940 28500 46992 28552
rect 19984 28432 20036 28484
rect 28264 28432 28316 28484
rect 28540 28432 28592 28484
rect 30380 28432 30432 28484
rect 14464 28364 14516 28416
rect 15752 28407 15804 28416
rect 15752 28373 15761 28407
rect 15761 28373 15795 28407
rect 15795 28373 15804 28407
rect 15752 28364 15804 28373
rect 19340 28364 19392 28416
rect 24124 28364 24176 28416
rect 24308 28364 24360 28416
rect 29000 28364 29052 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 17224 28160 17276 28212
rect 14464 28135 14516 28144
rect 14464 28101 14473 28135
rect 14473 28101 14507 28135
rect 14507 28101 14516 28135
rect 14464 28092 14516 28101
rect 18604 28092 18656 28144
rect 12716 27956 12768 28008
rect 15844 27999 15896 28008
rect 15844 27965 15853 27999
rect 15853 27965 15887 27999
rect 15887 27965 15896 27999
rect 15844 27956 15896 27965
rect 17040 27999 17092 28008
rect 17040 27965 17049 27999
rect 17049 27965 17083 27999
rect 17083 27965 17092 27999
rect 17040 27956 17092 27965
rect 17960 27956 18012 28008
rect 21180 28160 21232 28212
rect 19984 28092 20036 28144
rect 21456 28092 21508 28144
rect 26240 28160 26292 28212
rect 30932 28160 30984 28212
rect 34520 28160 34572 28212
rect 22192 28092 22244 28144
rect 28632 28135 28684 28144
rect 20720 28024 20772 28076
rect 20996 28067 21048 28076
rect 20996 28033 21005 28067
rect 21005 28033 21039 28067
rect 21039 28033 21048 28067
rect 20996 28024 21048 28033
rect 21088 28024 21140 28076
rect 19156 27888 19208 27940
rect 23388 28024 23440 28076
rect 23664 28024 23716 28076
rect 28632 28101 28641 28135
rect 28641 28101 28675 28135
rect 28675 28101 28684 28135
rect 28632 28092 28684 28101
rect 34796 28092 34848 28144
rect 24676 28024 24728 28076
rect 22008 27888 22060 27940
rect 24400 27956 24452 28008
rect 25136 27956 25188 28008
rect 25320 27956 25372 28008
rect 27528 28024 27580 28076
rect 28448 28067 28500 28076
rect 28448 28033 28457 28067
rect 28457 28033 28491 28067
rect 28491 28033 28500 28067
rect 28448 28024 28500 28033
rect 31300 28024 31352 28076
rect 45468 28024 45520 28076
rect 47308 28024 47360 28076
rect 28540 27956 28592 28008
rect 30288 27999 30340 28008
rect 30288 27965 30297 27999
rect 30297 27965 30331 27999
rect 30331 27965 30340 27999
rect 30288 27956 30340 27965
rect 33140 27956 33192 28008
rect 34152 27999 34204 28008
rect 34152 27965 34161 27999
rect 34161 27965 34195 27999
rect 34195 27965 34204 27999
rect 34152 27956 34204 27965
rect 24124 27888 24176 27940
rect 19432 27820 19484 27872
rect 21088 27820 21140 27872
rect 23112 27863 23164 27872
rect 23112 27829 23121 27863
rect 23121 27829 23155 27863
rect 23155 27829 23164 27863
rect 23112 27820 23164 27829
rect 23388 27820 23440 27872
rect 24860 27888 24912 27940
rect 24308 27820 24360 27872
rect 28540 27820 28592 27872
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3332 27616 3384 27668
rect 19432 27659 19484 27668
rect 19432 27625 19441 27659
rect 19441 27625 19475 27659
rect 19475 27625 19484 27659
rect 19432 27616 19484 27625
rect 19524 27616 19576 27668
rect 20996 27616 21048 27668
rect 21456 27616 21508 27668
rect 23112 27616 23164 27668
rect 23664 27616 23716 27668
rect 25596 27616 25648 27668
rect 27620 27659 27672 27668
rect 27620 27625 27629 27659
rect 27629 27625 27663 27659
rect 27663 27625 27672 27659
rect 27620 27616 27672 27625
rect 28448 27616 28500 27668
rect 34152 27659 34204 27668
rect 34152 27625 34161 27659
rect 34161 27625 34195 27659
rect 34195 27625 34204 27659
rect 34152 27616 34204 27625
rect 43720 27616 43772 27668
rect 45560 27616 45612 27668
rect 18604 27591 18656 27600
rect 15752 27480 15804 27532
rect 18604 27557 18613 27591
rect 18613 27557 18647 27591
rect 18647 27557 18656 27591
rect 18604 27548 18656 27557
rect 18696 27412 18748 27464
rect 20168 27480 20220 27532
rect 21088 27548 21140 27600
rect 23388 27548 23440 27600
rect 25320 27548 25372 27600
rect 30380 27548 30432 27600
rect 33140 27548 33192 27600
rect 34796 27548 34848 27600
rect 20996 27480 21048 27532
rect 21824 27480 21876 27532
rect 23756 27480 23808 27532
rect 24032 27480 24084 27532
rect 27988 27480 28040 27532
rect 34152 27480 34204 27532
rect 46940 27548 46992 27600
rect 47676 27480 47728 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 21088 27455 21140 27464
rect 21088 27421 21097 27455
rect 21097 27421 21131 27455
rect 21131 27421 21140 27455
rect 21088 27412 21140 27421
rect 17592 27344 17644 27396
rect 21272 27412 21324 27464
rect 21916 27412 21968 27464
rect 23112 27455 23164 27464
rect 23112 27421 23121 27455
rect 23121 27421 23155 27455
rect 23155 27421 23164 27455
rect 23112 27412 23164 27421
rect 27252 27412 27304 27464
rect 28172 27455 28224 27464
rect 28172 27421 28181 27455
rect 28181 27421 28215 27455
rect 28215 27421 28224 27455
rect 28172 27412 28224 27421
rect 28816 27412 28868 27464
rect 29552 27412 29604 27464
rect 31208 27412 31260 27464
rect 34520 27412 34572 27464
rect 35532 27412 35584 27464
rect 23388 27387 23440 27396
rect 23388 27353 23397 27387
rect 23397 27353 23431 27387
rect 23431 27353 23440 27387
rect 23388 27344 23440 27353
rect 23940 27344 23992 27396
rect 24400 27387 24452 27396
rect 24400 27353 24409 27387
rect 24409 27353 24443 27387
rect 24443 27353 24452 27387
rect 24400 27344 24452 27353
rect 24584 27387 24636 27396
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 27436 27344 27488 27396
rect 28632 27344 28684 27396
rect 21364 27276 21416 27328
rect 23204 27276 23256 27328
rect 23756 27319 23808 27328
rect 23756 27285 23765 27319
rect 23765 27285 23799 27319
rect 23799 27285 23808 27319
rect 23756 27276 23808 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 20720 27115 20772 27124
rect 20720 27081 20729 27115
rect 20729 27081 20763 27115
rect 20763 27081 20772 27115
rect 20720 27072 20772 27081
rect 22192 27115 22244 27124
rect 22192 27081 22201 27115
rect 22201 27081 22235 27115
rect 22235 27081 22244 27115
rect 22192 27072 22244 27081
rect 17040 27004 17092 27056
rect 19340 27004 19392 27056
rect 19984 27004 20036 27056
rect 21824 27047 21876 27056
rect 21824 27013 21833 27047
rect 21833 27013 21867 27047
rect 21867 27013 21876 27047
rect 21824 27004 21876 27013
rect 22008 27047 22060 27056
rect 22008 27013 22017 27047
rect 22017 27013 22051 27047
rect 22051 27013 22060 27047
rect 22008 27004 22060 27013
rect 23940 27072 23992 27124
rect 24584 27072 24636 27124
rect 27252 27072 27304 27124
rect 28172 27072 28224 27124
rect 32312 27072 32364 27124
rect 24308 27004 24360 27056
rect 25320 27004 25372 27056
rect 29644 27004 29696 27056
rect 33140 27004 33192 27056
rect 34244 27004 34296 27056
rect 23296 26979 23348 26988
rect 23296 26945 23305 26979
rect 23305 26945 23339 26979
rect 23339 26945 23348 26979
rect 23296 26936 23348 26945
rect 24032 26979 24084 26988
rect 12348 26911 12400 26920
rect 12348 26877 12357 26911
rect 12357 26877 12391 26911
rect 12391 26877 12400 26911
rect 12348 26868 12400 26877
rect 13728 26868 13780 26920
rect 16856 26911 16908 26920
rect 16856 26877 16865 26911
rect 16865 26877 16899 26911
rect 16899 26877 16908 26911
rect 16856 26868 16908 26877
rect 17132 26911 17184 26920
rect 17132 26877 17141 26911
rect 17141 26877 17175 26911
rect 17175 26877 17184 26911
rect 17132 26868 17184 26877
rect 18972 26911 19024 26920
rect 18972 26877 18981 26911
rect 18981 26877 19015 26911
rect 19015 26877 19024 26911
rect 18972 26868 19024 26877
rect 22652 26868 22704 26920
rect 24032 26945 24041 26979
rect 24041 26945 24075 26979
rect 24075 26945 24084 26979
rect 24032 26936 24084 26945
rect 27620 26936 27672 26988
rect 27988 26979 28040 26988
rect 27988 26945 27997 26979
rect 27997 26945 28031 26979
rect 28031 26945 28040 26979
rect 27988 26936 28040 26945
rect 31208 26936 31260 26988
rect 34060 26936 34112 26988
rect 12624 26843 12676 26852
rect 12624 26809 12633 26843
rect 12633 26809 12667 26843
rect 12667 26809 12676 26843
rect 12624 26800 12676 26809
rect 28356 26868 28408 26920
rect 32404 26911 32456 26920
rect 32404 26877 32413 26911
rect 32413 26877 32447 26911
rect 32447 26877 32456 26911
rect 32404 26868 32456 26877
rect 33968 26868 34020 26920
rect 47124 26868 47176 26920
rect 48044 26868 48096 26920
rect 18788 26732 18840 26784
rect 26148 26732 26200 26784
rect 34796 26732 34848 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 12348 26528 12400 26580
rect 16856 26528 16908 26580
rect 19984 26528 20036 26580
rect 23112 26528 23164 26580
rect 23572 26528 23624 26580
rect 23940 26528 23992 26580
rect 25320 26571 25372 26580
rect 25320 26537 25329 26571
rect 25329 26537 25363 26571
rect 25363 26537 25372 26571
rect 25320 26528 25372 26537
rect 28356 26571 28408 26580
rect 28356 26537 28365 26571
rect 28365 26537 28399 26571
rect 28399 26537 28408 26571
rect 28356 26528 28408 26537
rect 29644 26571 29696 26580
rect 29644 26537 29653 26571
rect 29653 26537 29687 26571
rect 29687 26537 29696 26571
rect 29644 26528 29696 26537
rect 32404 26528 32456 26580
rect 34152 26571 34204 26580
rect 34152 26537 34161 26571
rect 34161 26537 34195 26571
rect 34195 26537 34204 26571
rect 34152 26528 34204 26537
rect 18788 26460 18840 26512
rect 8300 26392 8352 26444
rect 18972 26392 19024 26444
rect 23112 26392 23164 26444
rect 24584 26460 24636 26512
rect 27620 26460 27672 26512
rect 29552 26460 29604 26512
rect 31024 26435 31076 26444
rect 31024 26401 31033 26435
rect 31033 26401 31067 26435
rect 31067 26401 31076 26435
rect 31024 26392 31076 26401
rect 31484 26392 31536 26444
rect 34428 26392 34480 26444
rect 11888 26367 11940 26376
rect 11888 26333 11897 26367
rect 11897 26333 11931 26367
rect 11931 26333 11940 26367
rect 11888 26324 11940 26333
rect 12716 26367 12768 26376
rect 12440 26256 12492 26308
rect 12716 26333 12725 26367
rect 12725 26333 12759 26367
rect 12759 26333 12768 26367
rect 12716 26324 12768 26333
rect 13084 26324 13136 26376
rect 14832 26324 14884 26376
rect 13360 26256 13412 26308
rect 14188 26299 14240 26308
rect 14188 26265 14197 26299
rect 14197 26265 14231 26299
rect 14231 26265 14240 26299
rect 14188 26256 14240 26265
rect 13268 26231 13320 26240
rect 13268 26197 13277 26231
rect 13277 26197 13311 26231
rect 13311 26197 13320 26231
rect 13268 26188 13320 26197
rect 15292 26324 15344 26376
rect 18512 26367 18564 26376
rect 18512 26333 18521 26367
rect 18521 26333 18555 26367
rect 18555 26333 18564 26367
rect 19248 26367 19300 26376
rect 18512 26324 18564 26333
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 16948 26256 17000 26308
rect 18696 26256 18748 26308
rect 25044 26324 25096 26376
rect 16304 26188 16356 26240
rect 22192 26256 22244 26308
rect 22560 26256 22612 26308
rect 24492 26256 24544 26308
rect 26148 26324 26200 26376
rect 27344 26367 27396 26376
rect 27344 26333 27353 26367
rect 27353 26333 27387 26367
rect 27387 26333 27396 26367
rect 27344 26324 27396 26333
rect 28540 26367 28592 26376
rect 28540 26333 28549 26367
rect 28549 26333 28583 26367
rect 28583 26333 28592 26367
rect 28540 26324 28592 26333
rect 29552 26367 29604 26376
rect 29552 26333 29561 26367
rect 29561 26333 29595 26367
rect 29595 26333 29604 26367
rect 29552 26324 29604 26333
rect 30380 26324 30432 26376
rect 32312 26367 32364 26376
rect 32312 26333 32321 26367
rect 32321 26333 32355 26367
rect 32355 26333 32364 26367
rect 32312 26324 32364 26333
rect 33968 26367 34020 26376
rect 33968 26333 33977 26367
rect 33977 26333 34011 26367
rect 34011 26333 34020 26367
rect 33968 26324 34020 26333
rect 34244 26324 34296 26376
rect 43720 26392 43772 26444
rect 34704 26367 34756 26376
rect 34704 26333 34713 26367
rect 34713 26333 34747 26367
rect 34747 26333 34756 26367
rect 34704 26324 34756 26333
rect 36636 26324 36688 26376
rect 34980 26299 35032 26308
rect 34980 26265 34989 26299
rect 34989 26265 35023 26299
rect 35023 26265 35032 26299
rect 34980 26256 35032 26265
rect 35992 26256 36044 26308
rect 37648 26299 37700 26308
rect 37648 26265 37657 26299
rect 37657 26265 37691 26299
rect 37691 26265 37700 26299
rect 37648 26256 37700 26265
rect 33876 26231 33928 26240
rect 33876 26197 33885 26231
rect 33885 26197 33919 26231
rect 33919 26197 33928 26231
rect 33876 26188 33928 26197
rect 34060 26188 34112 26240
rect 42156 26188 42208 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 22560 26027 22612 26036
rect 22560 25993 22569 26027
rect 22569 25993 22603 26027
rect 22603 25993 22612 26027
rect 22560 25984 22612 25993
rect 23112 26027 23164 26036
rect 23112 25993 23121 26027
rect 23121 25993 23155 26027
rect 23155 25993 23164 26027
rect 23112 25984 23164 25993
rect 33140 25984 33192 26036
rect 34704 25984 34756 26036
rect 34980 26027 35032 26036
rect 34980 25993 34989 26027
rect 34989 25993 35023 26027
rect 35023 25993 35032 26027
rect 34980 25984 35032 25993
rect 35992 25984 36044 26036
rect 37648 26027 37700 26036
rect 37648 25993 37657 26027
rect 37657 25993 37691 26027
rect 37691 25993 37700 26027
rect 37648 25984 37700 25993
rect 12624 25916 12676 25968
rect 14188 25916 14240 25968
rect 14832 25916 14884 25968
rect 11888 25891 11940 25900
rect 11888 25857 11897 25891
rect 11897 25857 11931 25891
rect 11931 25857 11940 25891
rect 11888 25848 11940 25857
rect 15108 25848 15160 25900
rect 15844 25848 15896 25900
rect 17132 25848 17184 25900
rect 18512 25916 18564 25968
rect 18052 25891 18104 25900
rect 18052 25857 18061 25891
rect 18061 25857 18095 25891
rect 18095 25857 18104 25891
rect 18052 25848 18104 25857
rect 22192 25848 22244 25900
rect 12440 25823 12492 25832
rect 12440 25789 12449 25823
rect 12449 25789 12483 25823
rect 12483 25789 12492 25823
rect 12440 25780 12492 25789
rect 13728 25780 13780 25832
rect 15292 25780 15344 25832
rect 22928 25848 22980 25900
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23756 25916 23808 25968
rect 31208 25916 31260 25968
rect 34060 25959 34112 25968
rect 23388 25848 23440 25857
rect 23664 25891 23716 25900
rect 23664 25857 23673 25891
rect 23673 25857 23707 25891
rect 23707 25857 23716 25891
rect 25412 25891 25464 25900
rect 23664 25848 23716 25857
rect 25412 25857 25421 25891
rect 25421 25857 25455 25891
rect 25455 25857 25464 25891
rect 25412 25848 25464 25857
rect 32496 25891 32548 25900
rect 32496 25857 32505 25891
rect 32505 25857 32539 25891
rect 32539 25857 32548 25891
rect 32496 25848 32548 25857
rect 34060 25925 34069 25959
rect 34069 25925 34103 25959
rect 34103 25925 34112 25959
rect 34060 25916 34112 25925
rect 34428 25916 34480 25968
rect 33968 25848 34020 25900
rect 34152 25848 34204 25900
rect 34796 25848 34848 25900
rect 35164 25916 35216 25968
rect 41420 25916 41472 25968
rect 35532 25891 35584 25900
rect 35532 25857 35541 25891
rect 35541 25857 35575 25891
rect 35575 25857 35584 25891
rect 35532 25848 35584 25857
rect 37556 25891 37608 25900
rect 37556 25857 37565 25891
rect 37565 25857 37599 25891
rect 37599 25857 37608 25891
rect 37556 25848 37608 25857
rect 41512 25891 41564 25900
rect 41512 25857 41521 25891
rect 41521 25857 41555 25891
rect 41555 25857 41564 25891
rect 41512 25848 41564 25857
rect 46756 25848 46808 25900
rect 24492 25780 24544 25832
rect 13820 25712 13872 25764
rect 18236 25755 18288 25764
rect 18236 25721 18245 25755
rect 18245 25721 18279 25755
rect 18279 25721 18288 25755
rect 18236 25712 18288 25721
rect 25320 25712 25372 25764
rect 28632 25780 28684 25832
rect 29920 25823 29972 25832
rect 29920 25789 29929 25823
rect 29929 25789 29963 25823
rect 29963 25789 29972 25823
rect 29920 25780 29972 25789
rect 36268 25780 36320 25832
rect 36452 25780 36504 25832
rect 45468 25780 45520 25832
rect 35164 25712 35216 25764
rect 11704 25687 11756 25696
rect 11704 25653 11713 25687
rect 11713 25653 11747 25687
rect 11747 25653 11756 25687
rect 11704 25644 11756 25653
rect 14924 25644 14976 25696
rect 15936 25644 15988 25696
rect 17408 25687 17460 25696
rect 17408 25653 17417 25687
rect 17417 25653 17451 25687
rect 17451 25653 17460 25687
rect 17408 25644 17460 25653
rect 33876 25644 33928 25696
rect 34244 25687 34296 25696
rect 34244 25653 34253 25687
rect 34253 25653 34287 25687
rect 34287 25653 34296 25687
rect 34244 25644 34296 25653
rect 34428 25687 34480 25696
rect 34428 25653 34437 25687
rect 34437 25653 34471 25687
rect 34471 25653 34480 25687
rect 34428 25644 34480 25653
rect 34520 25644 34572 25696
rect 41512 25644 41564 25696
rect 42340 25644 42392 25696
rect 47584 25644 47636 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 12440 25440 12492 25492
rect 13084 25440 13136 25492
rect 15292 25440 15344 25492
rect 17132 25440 17184 25492
rect 17408 25440 17460 25492
rect 16304 25372 16356 25424
rect 25964 25440 26016 25492
rect 30104 25372 30156 25424
rect 32496 25440 32548 25492
rect 35532 25440 35584 25492
rect 40040 25440 40092 25492
rect 11704 25347 11756 25356
rect 11704 25313 11713 25347
rect 11713 25313 11747 25347
rect 11747 25313 11756 25347
rect 11704 25304 11756 25313
rect 12532 25304 12584 25356
rect 14924 25347 14976 25356
rect 14924 25313 14933 25347
rect 14933 25313 14967 25347
rect 14967 25313 14976 25347
rect 14924 25304 14976 25313
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 13268 25168 13320 25220
rect 13360 25168 13412 25220
rect 17224 25236 17276 25288
rect 17408 25236 17460 25288
rect 18052 25304 18104 25356
rect 2044 25100 2096 25152
rect 12716 25100 12768 25152
rect 15200 25168 15252 25220
rect 15936 25168 15988 25220
rect 20720 25236 20772 25288
rect 21180 25279 21232 25288
rect 21180 25245 21189 25279
rect 21189 25245 21223 25279
rect 21223 25245 21232 25279
rect 21180 25236 21232 25245
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 24492 25279 24544 25288
rect 24492 25245 24501 25279
rect 24501 25245 24535 25279
rect 24535 25245 24544 25279
rect 24492 25236 24544 25245
rect 25412 25304 25464 25356
rect 25780 25304 25832 25356
rect 25964 25347 26016 25356
rect 25964 25313 25973 25347
rect 25973 25313 26007 25347
rect 26007 25313 26016 25347
rect 25964 25304 26016 25313
rect 26240 25304 26292 25356
rect 29276 25236 29328 25288
rect 29644 25279 29696 25288
rect 29644 25245 29653 25279
rect 29653 25245 29687 25279
rect 29687 25245 29696 25279
rect 29644 25236 29696 25245
rect 30380 25279 30432 25288
rect 30380 25245 30389 25279
rect 30389 25245 30423 25279
rect 30423 25245 30432 25279
rect 30380 25236 30432 25245
rect 19432 25168 19484 25220
rect 24676 25168 24728 25220
rect 37556 25372 37608 25424
rect 39396 25372 39448 25424
rect 31392 25304 31444 25356
rect 46664 25440 46716 25492
rect 46388 25372 46440 25424
rect 41696 25347 41748 25356
rect 41696 25313 41705 25347
rect 41705 25313 41739 25347
rect 41739 25313 41748 25347
rect 41696 25304 41748 25313
rect 42156 25347 42208 25356
rect 42156 25313 42165 25347
rect 42165 25313 42199 25347
rect 42199 25313 42208 25347
rect 42156 25304 42208 25313
rect 42340 25347 42392 25356
rect 42340 25313 42349 25347
rect 42349 25313 42383 25347
rect 42383 25313 42392 25347
rect 42340 25304 42392 25313
rect 46848 25347 46900 25356
rect 46848 25313 46857 25347
rect 46857 25313 46891 25347
rect 46891 25313 46900 25347
rect 46848 25304 46900 25313
rect 39120 25279 39172 25288
rect 39120 25245 39129 25279
rect 39129 25245 39163 25279
rect 39163 25245 39172 25279
rect 39120 25236 39172 25245
rect 30840 25168 30892 25220
rect 34520 25168 34572 25220
rect 15568 25100 15620 25152
rect 21548 25100 21600 25152
rect 24952 25100 25004 25152
rect 30380 25100 30432 25152
rect 33968 25100 34020 25152
rect 45192 25236 45244 25288
rect 40040 25211 40092 25220
rect 40040 25177 40049 25211
rect 40049 25177 40083 25211
rect 40083 25177 40092 25211
rect 40040 25168 40092 25177
rect 43996 25211 44048 25220
rect 43996 25177 44005 25211
rect 44005 25177 44039 25211
rect 44039 25177 44048 25211
rect 43996 25168 44048 25177
rect 45652 25211 45704 25220
rect 45652 25177 45661 25211
rect 45661 25177 45695 25211
rect 45695 25177 45704 25211
rect 45652 25168 45704 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 12440 24896 12492 24948
rect 12624 24896 12676 24948
rect 13728 24896 13780 24948
rect 19432 24939 19484 24948
rect 19432 24905 19441 24939
rect 19441 24905 19475 24939
rect 19475 24905 19484 24939
rect 19432 24896 19484 24905
rect 20536 24896 20588 24948
rect 29920 24896 29972 24948
rect 34244 24896 34296 24948
rect 12072 24803 12124 24812
rect 12072 24769 12081 24803
rect 12081 24769 12115 24803
rect 12115 24769 12124 24803
rect 12072 24760 12124 24769
rect 12624 24692 12676 24744
rect 13084 24760 13136 24812
rect 13360 24760 13412 24812
rect 13820 24760 13872 24812
rect 13544 24692 13596 24744
rect 15568 24828 15620 24880
rect 20720 24828 20772 24880
rect 15108 24692 15160 24744
rect 12716 24624 12768 24676
rect 15292 24624 15344 24676
rect 16948 24803 17000 24812
rect 16948 24769 16957 24803
rect 16957 24769 16991 24803
rect 16991 24769 17000 24803
rect 16948 24760 17000 24769
rect 17132 24760 17184 24812
rect 19524 24803 19576 24812
rect 19524 24769 19533 24803
rect 19533 24769 19567 24803
rect 19567 24769 19576 24803
rect 19524 24760 19576 24769
rect 20168 24760 20220 24812
rect 20904 24803 20956 24812
rect 20904 24769 20913 24803
rect 20913 24769 20947 24803
rect 20947 24769 20956 24803
rect 21824 24803 21876 24812
rect 20904 24760 20956 24769
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 26148 24803 26200 24812
rect 26148 24769 26157 24803
rect 26157 24769 26191 24803
rect 26191 24769 26200 24803
rect 26148 24760 26200 24769
rect 26516 24760 26568 24812
rect 27620 24760 27672 24812
rect 30380 24803 30432 24812
rect 30380 24769 30389 24803
rect 30389 24769 30423 24803
rect 30423 24769 30432 24803
rect 30380 24760 30432 24769
rect 31300 24760 31352 24812
rect 32128 24803 32180 24812
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 12440 24599 12492 24608
rect 12440 24565 12449 24599
rect 12449 24565 12483 24599
rect 12483 24565 12492 24599
rect 12440 24556 12492 24565
rect 17684 24599 17736 24608
rect 17684 24565 17693 24599
rect 17693 24565 17727 24599
rect 17727 24565 17736 24599
rect 17684 24556 17736 24565
rect 19248 24667 19300 24676
rect 19248 24633 19257 24667
rect 19257 24633 19291 24667
rect 19291 24633 19300 24667
rect 19248 24624 19300 24633
rect 21180 24624 21232 24676
rect 19524 24556 19576 24608
rect 19984 24556 20036 24608
rect 21272 24556 21324 24608
rect 23388 24692 23440 24744
rect 28724 24692 28776 24744
rect 31116 24735 31168 24744
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 31668 24692 31720 24744
rect 33876 24760 33928 24812
rect 34244 24760 34296 24812
rect 36268 24760 36320 24812
rect 38752 24803 38804 24812
rect 32404 24692 32456 24744
rect 33968 24692 34020 24744
rect 34152 24735 34204 24744
rect 34152 24701 34161 24735
rect 34161 24701 34195 24735
rect 34195 24701 34204 24735
rect 34152 24692 34204 24701
rect 35256 24692 35308 24744
rect 36636 24735 36688 24744
rect 36636 24701 36645 24735
rect 36645 24701 36679 24735
rect 36679 24701 36688 24735
rect 36636 24692 36688 24701
rect 38752 24769 38761 24803
rect 38761 24769 38795 24803
rect 38795 24769 38804 24803
rect 38752 24760 38804 24769
rect 39396 24803 39448 24812
rect 39396 24769 39405 24803
rect 39405 24769 39439 24803
rect 39439 24769 39448 24803
rect 39396 24760 39448 24769
rect 44916 24803 44968 24812
rect 44916 24769 44925 24803
rect 44925 24769 44959 24803
rect 44959 24769 44968 24803
rect 44916 24760 44968 24769
rect 45652 24760 45704 24812
rect 47216 24760 47268 24812
rect 47952 24760 48004 24812
rect 41236 24735 41288 24744
rect 41236 24701 41245 24735
rect 41245 24701 41279 24735
rect 41279 24701 41288 24735
rect 41236 24692 41288 24701
rect 24768 24624 24820 24676
rect 26240 24556 26292 24608
rect 26424 24556 26476 24608
rect 26976 24599 27028 24608
rect 26976 24565 26985 24599
rect 26985 24565 27019 24599
rect 27019 24565 27028 24599
rect 26976 24556 27028 24565
rect 27896 24599 27948 24608
rect 27896 24565 27905 24599
rect 27905 24565 27939 24599
rect 27939 24565 27948 24599
rect 27896 24556 27948 24565
rect 28540 24599 28592 24608
rect 28540 24565 28549 24599
rect 28549 24565 28583 24599
rect 28583 24565 28592 24599
rect 28540 24556 28592 24565
rect 31944 24556 31996 24608
rect 32772 24556 32824 24608
rect 34796 24556 34848 24608
rect 45560 24624 45612 24676
rect 39028 24556 39080 24608
rect 46296 24556 46348 24608
rect 47676 24599 47728 24608
rect 47676 24565 47685 24599
rect 47685 24565 47719 24599
rect 47719 24565 47728 24599
rect 47676 24556 47728 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 12532 24352 12584 24404
rect 15200 24395 15252 24404
rect 15200 24361 15209 24395
rect 15209 24361 15243 24395
rect 15243 24361 15252 24395
rect 15200 24352 15252 24361
rect 20720 24395 20772 24404
rect 20720 24361 20729 24395
rect 20729 24361 20763 24395
rect 20763 24361 20772 24395
rect 20720 24352 20772 24361
rect 12072 24284 12124 24336
rect 32312 24352 32364 24404
rect 32496 24352 32548 24404
rect 34244 24352 34296 24404
rect 36268 24352 36320 24404
rect 38752 24352 38804 24404
rect 44916 24352 44968 24404
rect 20904 24216 20956 24268
rect 21272 24259 21324 24268
rect 21272 24225 21281 24259
rect 21281 24225 21315 24259
rect 21315 24225 21324 24259
rect 21272 24216 21324 24225
rect 21548 24259 21600 24268
rect 21548 24225 21557 24259
rect 21557 24225 21591 24259
rect 21591 24225 21600 24259
rect 21548 24216 21600 24225
rect 25688 24259 25740 24268
rect 25688 24225 25697 24259
rect 25697 24225 25731 24259
rect 25731 24225 25740 24259
rect 25688 24216 25740 24225
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 13820 24148 13872 24200
rect 15936 24191 15988 24200
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 16948 24191 17000 24200
rect 16948 24157 16957 24191
rect 16957 24157 16991 24191
rect 16991 24157 17000 24191
rect 16948 24148 17000 24157
rect 19248 24148 19300 24200
rect 13360 24123 13412 24132
rect 13360 24089 13369 24123
rect 13369 24089 13403 24123
rect 13403 24089 13412 24123
rect 13360 24080 13412 24089
rect 14464 24080 14516 24132
rect 16764 24080 16816 24132
rect 16672 24012 16724 24064
rect 17684 24080 17736 24132
rect 19340 24123 19392 24132
rect 19340 24089 19349 24123
rect 19349 24089 19383 24123
rect 19383 24089 19392 24123
rect 19340 24080 19392 24089
rect 19524 24148 19576 24200
rect 20444 24191 20496 24200
rect 20444 24157 20453 24191
rect 20453 24157 20487 24191
rect 20487 24157 20496 24191
rect 20444 24148 20496 24157
rect 26056 24216 26108 24268
rect 30564 24284 30616 24336
rect 31668 24284 31720 24336
rect 33232 24284 33284 24336
rect 34152 24284 34204 24336
rect 35256 24327 35308 24336
rect 35256 24293 35265 24327
rect 35265 24293 35299 24327
rect 35299 24293 35308 24327
rect 35256 24284 35308 24293
rect 28724 24216 28776 24268
rect 40776 24284 40828 24336
rect 38568 24259 38620 24268
rect 38568 24225 38577 24259
rect 38577 24225 38611 24259
rect 38611 24225 38620 24259
rect 38568 24216 38620 24225
rect 20352 24080 20404 24132
rect 22836 24080 22888 24132
rect 26332 24148 26384 24200
rect 29552 24148 29604 24200
rect 30472 24191 30524 24200
rect 30472 24157 30481 24191
rect 30481 24157 30515 24191
rect 30515 24157 30524 24191
rect 30472 24148 30524 24157
rect 26516 24080 26568 24132
rect 18604 24012 18656 24064
rect 19432 24012 19484 24064
rect 20536 24012 20588 24064
rect 21916 24012 21968 24064
rect 23940 24012 23992 24064
rect 27896 24080 27948 24132
rect 30380 24080 30432 24132
rect 31300 24148 31352 24200
rect 29736 24055 29788 24064
rect 29736 24021 29745 24055
rect 29745 24021 29779 24055
rect 29779 24021 29788 24055
rect 29736 24012 29788 24021
rect 29828 24012 29880 24064
rect 32036 24080 32088 24132
rect 32772 24148 32824 24200
rect 33140 24191 33192 24200
rect 33140 24157 33149 24191
rect 33149 24157 33183 24191
rect 33183 24157 33192 24191
rect 33140 24148 33192 24157
rect 34244 24148 34296 24200
rect 35532 24148 35584 24200
rect 36084 24148 36136 24200
rect 31576 24012 31628 24064
rect 33600 24080 33652 24132
rect 37372 24080 37424 24132
rect 38568 24080 38620 24132
rect 47492 24284 47544 24336
rect 46296 24259 46348 24268
rect 46296 24225 46305 24259
rect 46305 24225 46339 24259
rect 46339 24225 46348 24259
rect 46296 24216 46348 24225
rect 47676 24216 47728 24268
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 42984 24191 43036 24200
rect 42984 24157 42993 24191
rect 42993 24157 43027 24191
rect 43027 24157 43036 24191
rect 42984 24148 43036 24157
rect 43168 24191 43220 24200
rect 43168 24157 43177 24191
rect 43177 24157 43211 24191
rect 43211 24157 43220 24191
rect 43168 24148 43220 24157
rect 33232 24012 33284 24064
rect 33876 24012 33928 24064
rect 45008 24080 45060 24132
rect 41236 24012 41288 24064
rect 43536 24012 43588 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 14832 23672 14884 23724
rect 19248 23808 19300 23860
rect 20444 23808 20496 23860
rect 20536 23851 20588 23860
rect 20536 23817 20545 23851
rect 20545 23817 20579 23851
rect 20579 23817 20588 23851
rect 20536 23808 20588 23817
rect 21088 23808 21140 23860
rect 22836 23851 22888 23860
rect 22836 23817 22845 23851
rect 22845 23817 22879 23851
rect 22879 23817 22888 23851
rect 22836 23808 22888 23817
rect 26332 23851 26384 23860
rect 26332 23817 26341 23851
rect 26341 23817 26375 23851
rect 26375 23817 26384 23851
rect 26332 23808 26384 23817
rect 20168 23783 20220 23792
rect 15844 23672 15896 23724
rect 16672 23715 16724 23724
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 14464 23536 14516 23588
rect 15108 23536 15160 23588
rect 17592 23604 17644 23656
rect 20168 23749 20177 23783
rect 20177 23749 20211 23783
rect 20211 23749 20220 23783
rect 20168 23740 20220 23749
rect 21916 23740 21968 23792
rect 23940 23783 23992 23792
rect 23940 23749 23949 23783
rect 23949 23749 23983 23783
rect 23983 23749 23992 23783
rect 23940 23740 23992 23749
rect 24952 23740 25004 23792
rect 29828 23808 29880 23860
rect 32128 23808 32180 23860
rect 32864 23808 32916 23860
rect 33140 23851 33192 23860
rect 33140 23817 33149 23851
rect 33149 23817 33183 23851
rect 33183 23817 33192 23851
rect 33140 23808 33192 23817
rect 33232 23808 33284 23860
rect 36084 23851 36136 23860
rect 19432 23672 19484 23724
rect 21824 23715 21876 23724
rect 19984 23604 20036 23656
rect 20168 23604 20220 23656
rect 20352 23604 20404 23656
rect 21824 23681 21833 23715
rect 21833 23681 21867 23715
rect 21867 23681 21876 23715
rect 21824 23672 21876 23681
rect 22744 23715 22796 23724
rect 22744 23681 22753 23715
rect 22753 23681 22787 23715
rect 22787 23681 22796 23715
rect 22744 23672 22796 23681
rect 18604 23536 18656 23588
rect 28540 23740 28592 23792
rect 26240 23672 26292 23724
rect 26516 23672 26568 23724
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 29644 23715 29696 23724
rect 29644 23681 29653 23715
rect 29653 23681 29687 23715
rect 29687 23681 29696 23715
rect 29644 23672 29696 23681
rect 30656 23715 30708 23724
rect 30656 23681 30665 23715
rect 30665 23681 30699 23715
rect 30699 23681 30708 23715
rect 30656 23672 30708 23681
rect 30932 23672 30984 23724
rect 27252 23647 27304 23656
rect 11796 23511 11848 23520
rect 11796 23477 11805 23511
rect 11805 23477 11839 23511
rect 11839 23477 11848 23511
rect 11796 23468 11848 23477
rect 17316 23468 17368 23520
rect 25596 23536 25648 23588
rect 27252 23613 27261 23647
rect 27261 23613 27295 23647
rect 27295 23613 27304 23647
rect 27252 23604 27304 23613
rect 27988 23604 28040 23656
rect 28632 23604 28684 23656
rect 31576 23715 31628 23724
rect 31576 23681 31585 23715
rect 31585 23681 31619 23715
rect 31619 23681 31628 23715
rect 31576 23672 31628 23681
rect 32772 23672 32824 23724
rect 33600 23715 33652 23724
rect 32496 23604 32548 23656
rect 33600 23681 33609 23715
rect 33609 23681 33643 23715
rect 33643 23681 33652 23715
rect 33600 23672 33652 23681
rect 21824 23511 21876 23520
rect 21824 23477 21833 23511
rect 21833 23477 21867 23511
rect 21867 23477 21876 23511
rect 21824 23468 21876 23477
rect 26608 23468 26660 23520
rect 29644 23468 29696 23520
rect 30748 23511 30800 23520
rect 30748 23477 30757 23511
rect 30757 23477 30791 23511
rect 30791 23477 30800 23511
rect 30748 23468 30800 23477
rect 35256 23740 35308 23792
rect 36084 23817 36093 23851
rect 36093 23817 36127 23851
rect 36127 23817 36136 23851
rect 36084 23808 36136 23817
rect 37372 23851 37424 23860
rect 37372 23817 37381 23851
rect 37381 23817 37415 23851
rect 37415 23817 37424 23851
rect 37372 23808 37424 23817
rect 39028 23783 39080 23792
rect 39028 23749 39037 23783
rect 39037 23749 39071 23783
rect 39071 23749 39080 23783
rect 39028 23740 39080 23749
rect 40776 23808 40828 23860
rect 45836 23808 45888 23860
rect 37280 23715 37332 23724
rect 37280 23681 37289 23715
rect 37289 23681 37323 23715
rect 37323 23681 37332 23715
rect 37280 23672 37332 23681
rect 34612 23647 34664 23656
rect 33876 23468 33928 23520
rect 34612 23613 34621 23647
rect 34621 23613 34655 23647
rect 34655 23613 34664 23647
rect 34612 23604 34664 23613
rect 42524 23672 42576 23724
rect 42800 23672 42852 23724
rect 43536 23715 43588 23724
rect 43536 23681 43545 23715
rect 43545 23681 43579 23715
rect 43579 23681 43588 23715
rect 43536 23672 43588 23681
rect 40500 23604 40552 23656
rect 41236 23647 41288 23656
rect 41236 23613 41245 23647
rect 41245 23613 41279 23647
rect 41279 23613 41288 23647
rect 41236 23604 41288 23613
rect 44640 23647 44692 23656
rect 44640 23613 44649 23647
rect 44649 23613 44683 23647
rect 44683 23613 44692 23647
rect 44640 23604 44692 23613
rect 46940 23672 46992 23724
rect 47216 23672 47268 23724
rect 46848 23604 46900 23656
rect 47860 23604 47912 23656
rect 34704 23468 34756 23520
rect 40500 23468 40552 23520
rect 47492 23536 47544 23588
rect 46572 23468 46624 23520
rect 46848 23511 46900 23520
rect 46848 23477 46857 23511
rect 46857 23477 46891 23511
rect 46891 23477 46900 23511
rect 46848 23468 46900 23477
rect 47032 23511 47084 23520
rect 47032 23477 47041 23511
rect 47041 23477 47075 23511
rect 47075 23477 47084 23511
rect 47032 23468 47084 23477
rect 47676 23511 47728 23520
rect 47676 23477 47685 23511
rect 47685 23477 47719 23511
rect 47719 23477 47728 23511
rect 47676 23468 47728 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 16948 23264 17000 23316
rect 19340 23264 19392 23316
rect 19524 23264 19576 23316
rect 23388 23264 23440 23316
rect 15936 23196 15988 23248
rect 17316 23196 17368 23248
rect 22744 23196 22796 23248
rect 25688 23196 25740 23248
rect 27252 23264 27304 23316
rect 11796 23128 11848 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 21824 23128 21876 23180
rect 29552 23196 29604 23248
rect 32036 23264 32088 23316
rect 32772 23307 32824 23316
rect 32772 23273 32781 23307
rect 32781 23273 32815 23307
rect 32815 23273 32824 23307
rect 32772 23264 32824 23273
rect 34704 23307 34756 23316
rect 34704 23273 34713 23307
rect 34713 23273 34747 23307
rect 34747 23273 34756 23307
rect 34704 23264 34756 23273
rect 43168 23307 43220 23316
rect 43168 23273 43177 23307
rect 43177 23273 43211 23307
rect 43211 23273 43220 23307
rect 43168 23264 43220 23273
rect 28448 23171 28500 23180
rect 28448 23137 28457 23171
rect 28457 23137 28491 23171
rect 28491 23137 28500 23171
rect 28448 23128 28500 23137
rect 29000 23128 29052 23180
rect 30748 23128 30800 23180
rect 31944 23128 31996 23180
rect 34612 23128 34664 23180
rect 40500 23171 40552 23180
rect 40500 23137 40509 23171
rect 40509 23137 40543 23171
rect 40543 23137 40552 23171
rect 40500 23128 40552 23137
rect 17316 23103 17368 23112
rect 12072 22992 12124 23044
rect 13084 22992 13136 23044
rect 14924 22992 14976 23044
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 19524 23103 19576 23112
rect 19524 23069 19533 23103
rect 19533 23069 19567 23103
rect 19567 23069 19576 23103
rect 19524 23060 19576 23069
rect 19984 23060 20036 23112
rect 20536 23060 20588 23112
rect 20904 23060 20956 23112
rect 22836 23060 22888 23112
rect 19432 22924 19484 22976
rect 24952 23060 25004 23112
rect 25228 22992 25280 23044
rect 28264 23060 28316 23112
rect 30104 23103 30156 23112
rect 30104 23069 30113 23103
rect 30113 23069 30147 23103
rect 30147 23069 30156 23103
rect 30104 23060 30156 23069
rect 33876 23103 33928 23112
rect 33876 23069 33885 23103
rect 33885 23069 33919 23103
rect 33919 23069 33928 23103
rect 33876 23060 33928 23069
rect 34152 23060 34204 23112
rect 34244 23060 34296 23112
rect 34704 23103 34756 23112
rect 34704 23069 34713 23103
rect 34713 23069 34747 23103
rect 34747 23069 34756 23103
rect 34704 23060 34756 23069
rect 40040 23103 40092 23112
rect 40040 23069 40049 23103
rect 40049 23069 40083 23103
rect 40083 23069 40092 23103
rect 40040 23060 40092 23069
rect 43444 23128 43496 23180
rect 47768 23264 47820 23316
rect 43536 23060 43588 23112
rect 47032 23196 47084 23248
rect 46296 23171 46348 23180
rect 46296 23137 46305 23171
rect 46305 23137 46339 23171
rect 46339 23137 46348 23171
rect 46296 23128 46348 23137
rect 47676 23128 47728 23180
rect 48228 23128 48280 23180
rect 28448 22992 28500 23044
rect 31576 22992 31628 23044
rect 32312 22992 32364 23044
rect 25596 22924 25648 22976
rect 27344 22924 27396 22976
rect 31944 22924 31996 22976
rect 32220 22924 32272 22976
rect 45744 22992 45796 23044
rect 43720 22967 43772 22976
rect 43720 22933 43729 22967
rect 43729 22933 43763 22967
rect 43763 22933 43772 22967
rect 43720 22924 43772 22933
rect 45376 22924 45428 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 13084 22763 13136 22772
rect 13084 22729 13093 22763
rect 13093 22729 13127 22763
rect 13127 22729 13136 22763
rect 13084 22720 13136 22729
rect 22836 22763 22888 22772
rect 22836 22729 22845 22763
rect 22845 22729 22879 22763
rect 22879 22729 22888 22763
rect 22836 22720 22888 22729
rect 28264 22720 28316 22772
rect 30932 22720 30984 22772
rect 32312 22720 32364 22772
rect 40040 22720 40092 22772
rect 13544 22652 13596 22704
rect 21364 22652 21416 22704
rect 28448 22652 28500 22704
rect 29000 22695 29052 22704
rect 29000 22661 29009 22695
rect 29009 22661 29043 22695
rect 29043 22661 29052 22695
rect 29000 22652 29052 22661
rect 29736 22652 29788 22704
rect 11980 22584 12032 22636
rect 12348 22584 12400 22636
rect 12992 22627 13044 22636
rect 12992 22593 13001 22627
rect 13001 22593 13035 22627
rect 13035 22593 13044 22627
rect 12992 22584 13044 22593
rect 18236 22584 18288 22636
rect 22744 22627 22796 22636
rect 22744 22593 22753 22627
rect 22753 22593 22787 22627
rect 22787 22593 22796 22627
rect 22744 22584 22796 22593
rect 25596 22627 25648 22636
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 27344 22584 27396 22636
rect 12072 22559 12124 22568
rect 12072 22525 12081 22559
rect 12081 22525 12115 22559
rect 12115 22525 12124 22559
rect 12072 22516 12124 22525
rect 29552 22516 29604 22568
rect 15200 22423 15252 22432
rect 15200 22389 15209 22423
rect 15209 22389 15243 22423
rect 15243 22389 15252 22423
rect 15200 22380 15252 22389
rect 25688 22380 25740 22432
rect 30196 22380 30248 22432
rect 30656 22584 30708 22636
rect 34704 22652 34756 22704
rect 42984 22720 43036 22772
rect 43720 22720 43772 22772
rect 45376 22695 45428 22704
rect 45376 22661 45385 22695
rect 45385 22661 45419 22695
rect 45419 22661 45428 22695
rect 45376 22652 45428 22661
rect 32036 22584 32088 22636
rect 40316 22584 40368 22636
rect 42800 22627 42852 22636
rect 42800 22593 42809 22627
rect 42809 22593 42843 22627
rect 42843 22593 42852 22627
rect 42800 22584 42852 22593
rect 43444 22627 43496 22636
rect 43444 22593 43453 22627
rect 43453 22593 43487 22627
rect 43487 22593 43496 22627
rect 43444 22584 43496 22593
rect 45192 22627 45244 22636
rect 43536 22516 43588 22568
rect 42524 22491 42576 22500
rect 42524 22457 42533 22491
rect 42533 22457 42567 22491
rect 42567 22457 42576 22491
rect 42524 22448 42576 22457
rect 45192 22593 45201 22627
rect 45201 22593 45235 22627
rect 45235 22593 45244 22627
rect 45192 22584 45244 22593
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 47952 22584 48004 22636
rect 45744 22559 45796 22568
rect 45744 22525 45753 22559
rect 45753 22525 45787 22559
rect 45787 22525 45796 22559
rect 45744 22516 45796 22525
rect 47676 22516 47728 22568
rect 31300 22423 31352 22432
rect 31300 22389 31309 22423
rect 31309 22389 31343 22423
rect 31343 22389 31352 22423
rect 31300 22380 31352 22389
rect 40132 22380 40184 22432
rect 45376 22380 45428 22432
rect 47492 22380 47544 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 25596 22176 25648 22228
rect 29552 22219 29604 22228
rect 29552 22185 29561 22219
rect 29561 22185 29595 22219
rect 29595 22185 29604 22219
rect 29552 22176 29604 22185
rect 35440 22176 35492 22228
rect 25964 22151 26016 22160
rect 20 22040 72 22092
rect 25964 22117 25973 22151
rect 25973 22117 26007 22151
rect 26007 22117 26016 22151
rect 25964 22108 26016 22117
rect 26700 22151 26752 22160
rect 26700 22117 26709 22151
rect 26709 22117 26743 22151
rect 26743 22117 26752 22151
rect 26700 22108 26752 22117
rect 14832 22083 14884 22092
rect 14832 22049 14841 22083
rect 14841 22049 14875 22083
rect 14875 22049 14884 22083
rect 14832 22040 14884 22049
rect 15200 22040 15252 22092
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 11888 21972 11940 22024
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 12440 21972 12492 22024
rect 14740 21972 14792 22024
rect 16304 21972 16356 22024
rect 19984 22040 20036 22092
rect 23388 22040 23440 22092
rect 27988 22040 28040 22092
rect 30564 22083 30616 22092
rect 30564 22049 30573 22083
rect 30573 22049 30607 22083
rect 30607 22049 30616 22083
rect 30564 22040 30616 22049
rect 31300 22083 31352 22092
rect 31300 22049 31309 22083
rect 31309 22049 31343 22083
rect 31343 22049 31352 22083
rect 31300 22040 31352 22049
rect 31668 22040 31720 22092
rect 31944 22040 31996 22092
rect 37280 22040 37332 22092
rect 40132 22040 40184 22092
rect 16580 21904 16632 21956
rect 11520 21836 11572 21888
rect 11888 21836 11940 21888
rect 16396 21836 16448 21888
rect 18236 21904 18288 21956
rect 22192 21972 22244 22024
rect 20628 21904 20680 21956
rect 20904 21947 20956 21956
rect 20904 21913 20913 21947
rect 20913 21913 20947 21947
rect 20947 21913 20956 21947
rect 20904 21904 20956 21913
rect 22744 21904 22796 21956
rect 16856 21836 16908 21888
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 19340 21879 19392 21888
rect 19340 21845 19349 21879
rect 19349 21845 19383 21879
rect 19383 21845 19392 21879
rect 19340 21836 19392 21845
rect 24952 21972 25004 22024
rect 26424 21972 26476 22024
rect 25136 21904 25188 21956
rect 29644 21972 29696 22024
rect 30196 21972 30248 22024
rect 30472 22015 30524 22024
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 35900 21972 35952 22024
rect 40316 22015 40368 22024
rect 40316 21981 40325 22015
rect 40325 21981 40359 22015
rect 40359 21981 40368 22015
rect 40316 21972 40368 21981
rect 44640 22040 44692 22092
rect 45376 22083 45428 22092
rect 45376 22049 45385 22083
rect 45385 22049 45419 22083
rect 45419 22049 45428 22083
rect 45376 22040 45428 22049
rect 45744 22083 45796 22092
rect 45744 22049 45753 22083
rect 45753 22049 45787 22083
rect 45787 22049 45796 22083
rect 45744 22040 45796 22049
rect 47860 22040 47912 22092
rect 40500 21972 40552 22024
rect 28540 21904 28592 21956
rect 31668 21904 31720 21956
rect 32220 21904 32272 21956
rect 43260 21972 43312 22024
rect 43444 21972 43496 22024
rect 45100 21972 45152 22024
rect 47768 21972 47820 22024
rect 47952 21972 48004 22024
rect 30472 21836 30524 21888
rect 32864 21836 32916 21888
rect 34612 21836 34664 21888
rect 40408 21836 40460 21888
rect 43444 21879 43496 21888
rect 43444 21845 43453 21879
rect 43453 21845 43487 21879
rect 43487 21845 43496 21879
rect 43444 21836 43496 21845
rect 44364 21879 44416 21888
rect 44364 21845 44373 21879
rect 44373 21845 44407 21879
rect 44407 21845 44416 21879
rect 44364 21836 44416 21845
rect 47676 21836 47728 21888
rect 47860 21879 47912 21888
rect 47860 21845 47869 21879
rect 47869 21845 47903 21879
rect 47903 21845 47912 21879
rect 47860 21836 47912 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3700 21632 3752 21684
rect 3516 21564 3568 21616
rect 11796 21564 11848 21616
rect 16396 21564 16448 21616
rect 18052 21632 18104 21684
rect 19984 21632 20036 21684
rect 20536 21632 20588 21684
rect 25228 21632 25280 21684
rect 25596 21632 25648 21684
rect 25964 21632 26016 21684
rect 26976 21632 27028 21684
rect 31208 21632 31260 21684
rect 32220 21675 32272 21684
rect 32220 21641 32229 21675
rect 32229 21641 32263 21675
rect 32263 21641 32272 21675
rect 32220 21632 32272 21641
rect 16856 21607 16908 21616
rect 16856 21573 16865 21607
rect 16865 21573 16899 21607
rect 16899 21573 16908 21607
rect 16856 21564 16908 21573
rect 19340 21564 19392 21616
rect 46112 21632 46164 21684
rect 46940 21632 46992 21684
rect 47860 21632 47912 21684
rect 35256 21607 35308 21616
rect 35256 21573 35265 21607
rect 35265 21573 35299 21607
rect 35299 21573 35308 21607
rect 35256 21564 35308 21573
rect 43076 21564 43128 21616
rect 45192 21607 45244 21616
rect 45192 21573 45201 21607
rect 45201 21573 45235 21607
rect 45235 21573 45244 21607
rect 45192 21564 45244 21573
rect 47584 21607 47636 21616
rect 47584 21573 47593 21607
rect 47593 21573 47627 21607
rect 47627 21573 47636 21607
rect 47584 21564 47636 21573
rect 47768 21607 47820 21616
rect 47768 21573 47777 21607
rect 47777 21573 47811 21607
rect 47811 21573 47820 21607
rect 47768 21564 47820 21573
rect 22192 21496 22244 21548
rect 23204 21539 23256 21548
rect 23204 21505 23213 21539
rect 23213 21505 23247 21539
rect 23247 21505 23256 21539
rect 23204 21496 23256 21505
rect 11704 21428 11756 21480
rect 14280 21471 14332 21480
rect 14280 21437 14289 21471
rect 14289 21437 14323 21471
rect 14323 21437 14332 21471
rect 14280 21428 14332 21437
rect 14464 21471 14516 21480
rect 14464 21437 14473 21471
rect 14473 21437 14507 21471
rect 14507 21437 14516 21471
rect 14464 21428 14516 21437
rect 16580 21360 16632 21412
rect 19984 21428 20036 21480
rect 21640 21428 21692 21480
rect 24676 21496 24728 21548
rect 24860 21539 24912 21548
rect 24860 21505 24869 21539
rect 24869 21505 24903 21539
rect 24903 21505 24912 21539
rect 24860 21496 24912 21505
rect 24952 21539 25004 21548
rect 24952 21505 24961 21539
rect 24961 21505 24995 21539
rect 24995 21505 25004 21539
rect 24952 21496 25004 21505
rect 25136 21496 25188 21548
rect 25596 21496 25648 21548
rect 27344 21539 27396 21548
rect 26056 21471 26108 21480
rect 26056 21437 26065 21471
rect 26065 21437 26099 21471
rect 26099 21437 26108 21471
rect 26056 21428 26108 21437
rect 22744 21360 22796 21412
rect 24400 21360 24452 21412
rect 24584 21292 24636 21344
rect 24860 21360 24912 21412
rect 27344 21505 27353 21539
rect 27353 21505 27387 21539
rect 27387 21505 27396 21539
rect 27344 21496 27396 21505
rect 28264 21539 28316 21548
rect 28264 21505 28273 21539
rect 28273 21505 28307 21539
rect 28307 21505 28316 21539
rect 28264 21496 28316 21505
rect 29644 21496 29696 21548
rect 32036 21496 32088 21548
rect 34612 21539 34664 21548
rect 34612 21505 34621 21539
rect 34621 21505 34655 21539
rect 34655 21505 34664 21539
rect 34612 21496 34664 21505
rect 42892 21496 42944 21548
rect 28632 21428 28684 21480
rect 29000 21471 29052 21480
rect 29000 21437 29009 21471
rect 29009 21437 29043 21471
rect 29043 21437 29052 21471
rect 29000 21428 29052 21437
rect 32956 21428 33008 21480
rect 27160 21292 27212 21344
rect 27712 21292 27764 21344
rect 36176 21471 36228 21480
rect 36176 21437 36185 21471
rect 36185 21437 36219 21471
rect 36219 21437 36228 21471
rect 36176 21428 36228 21437
rect 35256 21360 35308 21412
rect 44364 21496 44416 21548
rect 46204 21539 46256 21548
rect 46204 21505 46213 21539
rect 46213 21505 46247 21539
rect 46247 21505 46256 21539
rect 46204 21496 46256 21505
rect 44640 21471 44692 21480
rect 44640 21437 44649 21471
rect 44649 21437 44683 21471
rect 44683 21437 44692 21471
rect 44640 21428 44692 21437
rect 45652 21428 45704 21480
rect 43168 21335 43220 21344
rect 43168 21301 43177 21335
rect 43177 21301 43211 21335
rect 43211 21301 43220 21335
rect 43168 21292 43220 21301
rect 44272 21292 44324 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 12348 21088 12400 21140
rect 14464 21088 14516 21140
rect 20168 21088 20220 21140
rect 16580 21020 16632 21072
rect 17316 21020 17368 21072
rect 18328 21020 18380 21072
rect 23112 21088 23164 21140
rect 27160 21131 27212 21140
rect 3424 20952 3476 21004
rect 11520 20927 11572 20936
rect 11520 20893 11529 20927
rect 11529 20893 11563 20927
rect 11563 20893 11572 20927
rect 11520 20884 11572 20893
rect 12900 20884 12952 20936
rect 14372 20927 14424 20936
rect 14372 20893 14381 20927
rect 14381 20893 14415 20927
rect 14415 20893 14424 20927
rect 14372 20884 14424 20893
rect 14832 20927 14884 20936
rect 14832 20893 14841 20927
rect 14841 20893 14875 20927
rect 14875 20893 14884 20927
rect 14832 20884 14884 20893
rect 15936 20884 15988 20936
rect 16304 20884 16356 20936
rect 17132 20884 17184 20936
rect 11888 20816 11940 20868
rect 11704 20748 11756 20800
rect 17040 20816 17092 20868
rect 17316 20927 17368 20936
rect 17316 20893 17325 20927
rect 17325 20893 17359 20927
rect 17359 20893 17368 20927
rect 17316 20884 17368 20893
rect 18236 20884 18288 20936
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 19248 20884 19300 20893
rect 17592 20816 17644 20868
rect 18604 20816 18656 20868
rect 21640 20927 21692 20936
rect 21640 20893 21649 20927
rect 21649 20893 21683 20927
rect 21683 20893 21692 20927
rect 21640 20884 21692 20893
rect 23848 21020 23900 21072
rect 24400 20995 24452 21004
rect 23112 20816 23164 20868
rect 24400 20961 24409 20995
rect 24409 20961 24443 20995
rect 24443 20961 24452 20995
rect 24400 20952 24452 20961
rect 24584 20952 24636 21004
rect 25688 20995 25740 21004
rect 24676 20927 24728 20936
rect 24676 20893 24685 20927
rect 24685 20893 24719 20927
rect 24719 20893 24728 20927
rect 24676 20884 24728 20893
rect 24952 20884 25004 20936
rect 23572 20859 23624 20868
rect 14464 20748 14516 20800
rect 16580 20748 16632 20800
rect 16764 20791 16816 20800
rect 16764 20757 16773 20791
rect 16773 20757 16807 20791
rect 16807 20757 16816 20791
rect 16764 20748 16816 20757
rect 16948 20748 17000 20800
rect 18144 20791 18196 20800
rect 18144 20757 18153 20791
rect 18153 20757 18187 20791
rect 18187 20757 18196 20791
rect 18144 20748 18196 20757
rect 20720 20748 20772 20800
rect 22836 20748 22888 20800
rect 23572 20825 23581 20859
rect 23581 20825 23615 20859
rect 23615 20825 23624 20859
rect 23572 20816 23624 20825
rect 25688 20961 25697 20995
rect 25697 20961 25731 20995
rect 25731 20961 25740 20995
rect 25688 20952 25740 20961
rect 27160 21097 27169 21131
rect 27169 21097 27203 21131
rect 27203 21097 27212 21131
rect 27160 21088 27212 21097
rect 28632 21131 28684 21140
rect 28632 21097 28641 21131
rect 28641 21097 28675 21131
rect 28675 21097 28684 21131
rect 28632 21088 28684 21097
rect 25412 20927 25464 20936
rect 25412 20893 25421 20927
rect 25421 20893 25455 20927
rect 25455 20893 25464 20927
rect 25412 20884 25464 20893
rect 28540 20927 28592 20936
rect 28540 20893 28549 20927
rect 28549 20893 28583 20927
rect 28583 20893 28592 20927
rect 28540 20884 28592 20893
rect 29552 20927 29604 20936
rect 29552 20893 29561 20927
rect 29561 20893 29595 20927
rect 29595 20893 29604 20927
rect 29552 20884 29604 20893
rect 23388 20791 23440 20800
rect 23388 20757 23397 20791
rect 23397 20757 23431 20791
rect 23431 20757 23440 20791
rect 23388 20748 23440 20757
rect 23480 20791 23532 20800
rect 23480 20757 23489 20791
rect 23489 20757 23523 20791
rect 23523 20757 23532 20791
rect 23480 20748 23532 20757
rect 24768 20791 24820 20800
rect 24768 20757 24777 20791
rect 24777 20757 24811 20791
rect 24811 20757 24820 20791
rect 24768 20748 24820 20757
rect 25320 20748 25372 20800
rect 25688 20748 25740 20800
rect 26700 20816 26752 20868
rect 29736 20859 29788 20868
rect 27620 20748 27672 20800
rect 29736 20825 29745 20859
rect 29745 20825 29779 20859
rect 29779 20825 29788 20859
rect 29736 20816 29788 20825
rect 43076 21020 43128 21072
rect 45100 21088 45152 21140
rect 47216 21020 47268 21072
rect 36176 20952 36228 21004
rect 48136 20995 48188 21004
rect 35532 20859 35584 20868
rect 35532 20825 35541 20859
rect 35541 20825 35575 20859
rect 35575 20825 35584 20859
rect 35532 20816 35584 20825
rect 35900 20816 35952 20868
rect 36360 20816 36412 20868
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 42892 20884 42944 20936
rect 43076 20927 43128 20936
rect 43076 20893 43085 20927
rect 43085 20893 43119 20927
rect 43119 20893 43128 20927
rect 43076 20884 43128 20893
rect 43444 20927 43496 20936
rect 43444 20893 43453 20927
rect 43453 20893 43487 20927
rect 43487 20893 43496 20927
rect 43444 20884 43496 20893
rect 44732 20884 44784 20936
rect 46296 20927 46348 20936
rect 46296 20893 46305 20927
rect 46305 20893 46339 20927
rect 46339 20893 46348 20927
rect 46296 20884 46348 20893
rect 44364 20816 44416 20868
rect 47676 20816 47728 20868
rect 42616 20748 42668 20800
rect 44088 20791 44140 20800
rect 44088 20757 44097 20791
rect 44097 20757 44131 20791
rect 44131 20757 44140 20791
rect 44088 20748 44140 20757
rect 47216 20748 47268 20800
rect 47768 20748 47820 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3056 20544 3108 20596
rect 13636 20476 13688 20528
rect 11980 20451 12032 20460
rect 11980 20417 11989 20451
rect 11989 20417 12023 20451
rect 12023 20417 12032 20451
rect 11980 20408 12032 20417
rect 14096 20340 14148 20392
rect 14280 20340 14332 20392
rect 17040 20476 17092 20528
rect 19800 20476 19852 20528
rect 19892 20476 19944 20528
rect 20168 20519 20220 20528
rect 20168 20485 20193 20519
rect 20193 20485 20220 20519
rect 20168 20476 20220 20485
rect 14924 20340 14976 20392
rect 16304 20340 16356 20392
rect 16856 20408 16908 20460
rect 17868 20451 17920 20460
rect 17868 20417 17877 20451
rect 17877 20417 17911 20451
rect 17911 20417 17920 20451
rect 17868 20408 17920 20417
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 21824 20451 21876 20460
rect 21824 20417 21833 20451
rect 21833 20417 21867 20451
rect 21867 20417 21876 20451
rect 21824 20408 21876 20417
rect 23480 20544 23532 20596
rect 24768 20544 24820 20596
rect 25412 20544 25464 20596
rect 26240 20544 26292 20596
rect 29736 20544 29788 20596
rect 43076 20544 43128 20596
rect 43352 20587 43404 20596
rect 43352 20553 43361 20587
rect 43361 20553 43395 20587
rect 43395 20553 43404 20587
rect 43352 20544 43404 20553
rect 23572 20476 23624 20528
rect 24860 20476 24912 20528
rect 29000 20476 29052 20528
rect 26240 20408 26292 20460
rect 26976 20451 27028 20460
rect 26976 20417 26985 20451
rect 26985 20417 27019 20451
rect 27019 20417 27028 20451
rect 26976 20408 27028 20417
rect 29736 20408 29788 20460
rect 30380 20408 30432 20460
rect 30840 20408 30892 20460
rect 33416 20451 33468 20460
rect 33416 20417 33425 20451
rect 33425 20417 33459 20451
rect 33459 20417 33468 20451
rect 33416 20408 33468 20417
rect 42616 20451 42668 20460
rect 42616 20417 42625 20451
rect 42625 20417 42659 20451
rect 42659 20417 42668 20451
rect 42616 20408 42668 20417
rect 42800 20408 42852 20460
rect 43260 20451 43312 20460
rect 43260 20417 43269 20451
rect 43269 20417 43303 20451
rect 43303 20417 43312 20451
rect 43260 20408 43312 20417
rect 43628 20451 43680 20460
rect 43628 20417 43637 20451
rect 43637 20417 43671 20451
rect 43671 20417 43680 20451
rect 43628 20408 43680 20417
rect 14464 20272 14516 20324
rect 15108 20247 15160 20256
rect 15108 20213 15117 20247
rect 15117 20213 15151 20247
rect 15151 20213 15160 20247
rect 15108 20204 15160 20213
rect 16856 20247 16908 20256
rect 16856 20213 16865 20247
rect 16865 20213 16899 20247
rect 16899 20213 16908 20247
rect 16856 20204 16908 20213
rect 17224 20204 17276 20256
rect 20444 20272 20496 20324
rect 19800 20204 19852 20256
rect 43168 20340 43220 20392
rect 43812 20340 43864 20392
rect 28816 20272 28868 20324
rect 44272 20476 44324 20528
rect 47952 20519 48004 20528
rect 47952 20485 47961 20519
rect 47961 20485 47995 20519
rect 47995 20485 48004 20519
rect 47952 20476 48004 20485
rect 44364 20451 44416 20460
rect 44364 20417 44373 20451
rect 44373 20417 44407 20451
rect 44407 20417 44416 20451
rect 44364 20408 44416 20417
rect 44732 20408 44784 20460
rect 44456 20340 44508 20392
rect 45744 20383 45796 20392
rect 45744 20349 45753 20383
rect 45753 20349 45787 20383
rect 45787 20349 45796 20383
rect 45744 20340 45796 20349
rect 21732 20204 21784 20256
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 25320 20204 25372 20256
rect 30656 20204 30708 20256
rect 33232 20247 33284 20256
rect 33232 20213 33241 20247
rect 33241 20213 33275 20247
rect 33275 20213 33284 20247
rect 33232 20204 33284 20213
rect 43260 20204 43312 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 12900 20043 12952 20052
rect 12900 20009 12909 20043
rect 12909 20009 12943 20043
rect 12943 20009 12952 20043
rect 12900 20000 12952 20009
rect 14096 20043 14148 20052
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 14280 20000 14332 20052
rect 14924 20000 14976 20052
rect 17868 20000 17920 20052
rect 19800 20043 19852 20052
rect 15200 19932 15252 19984
rect 19800 20009 19809 20043
rect 19809 20009 19843 20043
rect 19843 20009 19852 20043
rect 19800 20000 19852 20009
rect 20168 20000 20220 20052
rect 1768 19796 1820 19848
rect 12992 19796 13044 19848
rect 14464 19796 14516 19848
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 17592 19864 17644 19916
rect 21824 19864 21876 19916
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19984 19796 20036 19848
rect 20720 19796 20772 19848
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 15108 19728 15160 19780
rect 16304 19771 16356 19780
rect 16304 19737 16329 19771
rect 16329 19737 16356 19771
rect 16304 19728 16356 19737
rect 19156 19728 19208 19780
rect 14280 19703 14332 19712
rect 14280 19669 14289 19703
rect 14289 19669 14323 19703
rect 14323 19669 14332 19703
rect 14280 19660 14332 19669
rect 15476 19660 15528 19712
rect 18052 19660 18104 19712
rect 20352 19728 20404 19780
rect 43628 20000 43680 20052
rect 43812 20000 43864 20052
rect 44180 20000 44232 20052
rect 44640 20000 44692 20052
rect 46296 20000 46348 20052
rect 23480 19932 23532 19984
rect 29184 19932 29236 19984
rect 32220 19932 32272 19984
rect 43352 19932 43404 19984
rect 45008 19932 45060 19984
rect 47400 19932 47452 19984
rect 25136 19864 25188 19916
rect 25412 19907 25464 19916
rect 25412 19873 25421 19907
rect 25421 19873 25455 19907
rect 25455 19873 25464 19907
rect 25412 19864 25464 19873
rect 30472 19907 30524 19916
rect 30472 19873 30481 19907
rect 30481 19873 30515 19907
rect 30515 19873 30524 19907
rect 30472 19864 30524 19873
rect 30656 19907 30708 19916
rect 30656 19873 30665 19907
rect 30665 19873 30699 19907
rect 30699 19873 30708 19907
rect 30656 19864 30708 19873
rect 23572 19771 23624 19780
rect 23572 19737 23581 19771
rect 23581 19737 23615 19771
rect 23615 19737 23624 19771
rect 23572 19728 23624 19737
rect 24124 19728 24176 19780
rect 24768 19728 24820 19780
rect 26976 19796 27028 19848
rect 29644 19796 29696 19848
rect 32312 19771 32364 19780
rect 32312 19737 32321 19771
rect 32321 19737 32355 19771
rect 32355 19737 32364 19771
rect 32312 19728 32364 19737
rect 33232 19771 33284 19780
rect 33232 19737 33241 19771
rect 33241 19737 33275 19771
rect 33275 19737 33284 19771
rect 34152 19771 34204 19780
rect 33232 19728 33284 19737
rect 34152 19737 34161 19771
rect 34161 19737 34195 19771
rect 34195 19737 34204 19771
rect 34152 19728 34204 19737
rect 42892 19864 42944 19916
rect 42984 19796 43036 19848
rect 43260 19839 43312 19848
rect 43260 19805 43269 19839
rect 43269 19805 43303 19839
rect 43303 19805 43312 19839
rect 43260 19796 43312 19805
rect 44548 19864 44600 19916
rect 44640 19796 44692 19848
rect 45652 19728 45704 19780
rect 47216 19728 47268 19780
rect 48136 19771 48188 19780
rect 48136 19737 48145 19771
rect 48145 19737 48179 19771
rect 48179 19737 48188 19771
rect 48136 19728 48188 19737
rect 20536 19703 20588 19712
rect 20536 19669 20545 19703
rect 20545 19669 20579 19703
rect 20579 19669 20588 19703
rect 20536 19660 20588 19669
rect 20628 19660 20680 19712
rect 21824 19703 21876 19712
rect 21824 19669 21833 19703
rect 21833 19669 21867 19703
rect 21867 19669 21876 19703
rect 21824 19660 21876 19669
rect 24676 19660 24728 19712
rect 29552 19703 29604 19712
rect 29552 19669 29561 19703
rect 29561 19669 29595 19703
rect 29595 19669 29604 19703
rect 29552 19660 29604 19669
rect 29920 19660 29972 19712
rect 31116 19660 31168 19712
rect 36544 19660 36596 19712
rect 45928 19660 45980 19712
rect 47400 19660 47452 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 13636 19456 13688 19508
rect 14924 19456 14976 19508
rect 19156 19456 19208 19508
rect 15108 19388 15160 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 12808 19363 12860 19372
rect 12808 19329 12817 19363
rect 12817 19329 12851 19363
rect 12851 19329 12860 19363
rect 12808 19320 12860 19329
rect 12992 19320 13044 19372
rect 13728 19320 13780 19372
rect 16948 19388 17000 19440
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 14280 19252 14332 19304
rect 15200 19252 15252 19304
rect 16856 19320 16908 19372
rect 18144 19388 18196 19440
rect 19064 19363 19116 19372
rect 19064 19329 19073 19363
rect 19073 19329 19107 19363
rect 19107 19329 19116 19363
rect 19064 19320 19116 19329
rect 19156 19320 19208 19372
rect 20628 19388 20680 19440
rect 20536 19320 20588 19372
rect 21824 19388 21876 19440
rect 23572 19456 23624 19508
rect 28080 19499 28132 19508
rect 28080 19465 28089 19499
rect 28089 19465 28123 19499
rect 28123 19465 28132 19499
rect 29644 19499 29696 19508
rect 28080 19456 28132 19465
rect 29644 19465 29653 19499
rect 29653 19465 29687 19499
rect 29687 19465 29696 19499
rect 29644 19456 29696 19465
rect 24860 19388 24912 19440
rect 28632 19431 28684 19440
rect 28632 19397 28641 19431
rect 28641 19397 28675 19431
rect 28675 19397 28684 19431
rect 28632 19388 28684 19397
rect 24032 19320 24084 19372
rect 26424 19320 26476 19372
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 21824 19295 21876 19304
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 24308 19295 24360 19304
rect 24308 19261 24317 19295
rect 24317 19261 24351 19295
rect 24351 19261 24360 19295
rect 24308 19252 24360 19261
rect 24584 19295 24636 19304
rect 24584 19261 24593 19295
rect 24593 19261 24627 19295
rect 24627 19261 24636 19295
rect 24584 19252 24636 19261
rect 29276 19295 29328 19304
rect 29276 19261 29285 19295
rect 29285 19261 29319 19295
rect 29319 19261 29328 19295
rect 33600 19456 33652 19508
rect 47492 19456 47544 19508
rect 47676 19499 47728 19508
rect 47676 19465 47685 19499
rect 47685 19465 47719 19499
rect 47719 19465 47728 19499
rect 47676 19456 47728 19465
rect 32220 19388 32272 19440
rect 46296 19431 46348 19440
rect 46296 19397 46305 19431
rect 46305 19397 46339 19431
rect 46339 19397 46348 19431
rect 46296 19388 46348 19397
rect 47124 19388 47176 19440
rect 36544 19320 36596 19372
rect 45008 19320 45060 19372
rect 45652 19363 45704 19372
rect 45652 19329 45661 19363
rect 45661 19329 45695 19363
rect 45695 19329 45704 19363
rect 45652 19320 45704 19329
rect 46204 19320 46256 19372
rect 47400 19320 47452 19372
rect 29276 19252 29328 19261
rect 13636 19116 13688 19168
rect 24400 19116 24452 19168
rect 27068 19159 27120 19168
rect 27068 19125 27077 19159
rect 27077 19125 27111 19159
rect 27111 19125 27120 19159
rect 27068 19116 27120 19125
rect 28448 19184 28500 19236
rect 34152 19252 34204 19304
rect 35532 19252 35584 19304
rect 37556 19252 37608 19304
rect 46940 19252 46992 19304
rect 33600 19227 33652 19236
rect 33600 19193 33609 19227
rect 33609 19193 33643 19227
rect 33643 19193 33652 19227
rect 33600 19184 33652 19193
rect 41328 19184 41380 19236
rect 47032 19184 47084 19236
rect 31392 19116 31444 19168
rect 42800 19116 42852 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 16948 18955 17000 18964
rect 12716 18844 12768 18896
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 11888 18683 11940 18692
rect 11888 18649 11897 18683
rect 11897 18649 11931 18683
rect 11931 18649 11940 18683
rect 11888 18640 11940 18649
rect 13544 18572 13596 18624
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 21824 18912 21876 18964
rect 24584 18912 24636 18964
rect 24860 18955 24912 18964
rect 24860 18921 24869 18955
rect 24869 18921 24903 18955
rect 24903 18921 24912 18955
rect 24860 18912 24912 18921
rect 24400 18844 24452 18896
rect 24768 18844 24820 18896
rect 33140 18955 33192 18964
rect 33140 18921 33149 18955
rect 33149 18921 33183 18955
rect 33183 18921 33192 18955
rect 33140 18912 33192 18921
rect 33416 18955 33468 18964
rect 33416 18921 33425 18955
rect 33425 18921 33459 18955
rect 33459 18921 33468 18955
rect 33416 18912 33468 18921
rect 41144 18912 41196 18964
rect 25412 18844 25464 18896
rect 47216 18912 47268 18964
rect 15476 18776 15528 18828
rect 24308 18776 24360 18828
rect 28540 18776 28592 18828
rect 30380 18776 30432 18828
rect 42800 18819 42852 18828
rect 42800 18785 42809 18819
rect 42809 18785 42843 18819
rect 42843 18785 42852 18819
rect 42800 18776 42852 18785
rect 15200 18751 15252 18760
rect 15200 18717 15209 18751
rect 15209 18717 15243 18751
rect 15243 18717 15252 18751
rect 15200 18708 15252 18717
rect 22008 18708 22060 18760
rect 23480 18751 23532 18760
rect 16764 18640 16816 18692
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 23480 18708 23532 18717
rect 23848 18708 23900 18760
rect 24676 18640 24728 18692
rect 25320 18708 25372 18760
rect 28448 18751 28500 18760
rect 28448 18717 28457 18751
rect 28457 18717 28491 18751
rect 28491 18717 28500 18751
rect 28448 18708 28500 18717
rect 28632 18751 28684 18760
rect 28632 18717 28641 18751
rect 28641 18717 28675 18751
rect 28675 18717 28684 18751
rect 28632 18708 28684 18717
rect 27068 18640 27120 18692
rect 29276 18640 29328 18692
rect 29920 18708 29972 18760
rect 32220 18708 32272 18760
rect 45192 18751 45244 18760
rect 32036 18640 32088 18692
rect 32128 18640 32180 18692
rect 32864 18640 32916 18692
rect 45192 18717 45201 18751
rect 45201 18717 45235 18751
rect 45235 18717 45244 18751
rect 45192 18708 45244 18717
rect 45376 18751 45428 18760
rect 45376 18717 45385 18751
rect 45385 18717 45419 18751
rect 45419 18717 45428 18751
rect 45376 18708 45428 18717
rect 47124 18776 47176 18828
rect 46204 18751 46256 18760
rect 46204 18717 46213 18751
rect 46213 18717 46247 18751
rect 46247 18717 46256 18751
rect 46204 18708 46256 18717
rect 46388 18708 46440 18760
rect 47032 18708 47084 18760
rect 47308 18751 47360 18760
rect 47308 18717 47317 18751
rect 47317 18717 47351 18751
rect 47351 18717 47360 18751
rect 47308 18708 47360 18717
rect 48044 18708 48096 18760
rect 44088 18640 44140 18692
rect 44456 18683 44508 18692
rect 44456 18649 44465 18683
rect 44465 18649 44499 18683
rect 44499 18649 44508 18683
rect 44456 18640 44508 18649
rect 46112 18683 46164 18692
rect 46112 18649 46121 18683
rect 46121 18649 46155 18683
rect 46155 18649 46164 18683
rect 46112 18640 46164 18649
rect 26424 18572 26476 18624
rect 44364 18572 44416 18624
rect 46480 18572 46532 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3424 18368 3476 18420
rect 11888 18343 11940 18352
rect 11888 18309 11897 18343
rect 11897 18309 11931 18343
rect 11931 18309 11940 18343
rect 11888 18300 11940 18309
rect 13636 18343 13688 18352
rect 13636 18309 13645 18343
rect 13645 18309 13679 18343
rect 13679 18309 13688 18343
rect 13636 18300 13688 18309
rect 14372 18300 14424 18352
rect 15200 18300 15252 18352
rect 16764 18343 16816 18352
rect 16764 18309 16773 18343
rect 16773 18309 16807 18343
rect 16807 18309 16816 18343
rect 16764 18300 16816 18309
rect 18604 18300 18656 18352
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 15660 18275 15712 18284
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 16672 18275 16724 18284
rect 16672 18241 16681 18275
rect 16681 18241 16715 18275
rect 16715 18241 16724 18275
rect 16672 18232 16724 18241
rect 14004 18164 14056 18216
rect 17684 18207 17736 18216
rect 17684 18173 17693 18207
rect 17693 18173 17727 18207
rect 17727 18173 17736 18207
rect 17684 18164 17736 18173
rect 19800 18164 19852 18216
rect 15384 18096 15436 18148
rect 19432 18139 19484 18148
rect 19432 18105 19441 18139
rect 19441 18105 19475 18139
rect 19475 18105 19484 18139
rect 19432 18096 19484 18105
rect 27712 18232 27764 18284
rect 27988 18300 28040 18352
rect 28080 18343 28132 18352
rect 28080 18309 28089 18343
rect 28089 18309 28123 18343
rect 28123 18309 28132 18343
rect 28080 18300 28132 18309
rect 24768 18164 24820 18216
rect 25320 18164 25372 18216
rect 23020 18096 23072 18148
rect 28172 18164 28224 18216
rect 29920 18207 29972 18216
rect 14924 18028 14976 18080
rect 15108 18071 15160 18080
rect 15108 18037 15117 18071
rect 15117 18037 15151 18071
rect 15151 18037 15160 18071
rect 15108 18028 15160 18037
rect 27804 18028 27856 18080
rect 28448 18096 28500 18148
rect 29920 18173 29929 18207
rect 29929 18173 29963 18207
rect 29963 18173 29972 18207
rect 29920 18164 29972 18173
rect 29184 18028 29236 18080
rect 30380 18096 30432 18148
rect 31024 18096 31076 18148
rect 44824 18368 44876 18420
rect 45192 18368 45244 18420
rect 32220 18300 32272 18352
rect 41328 18300 41380 18352
rect 32036 18232 32088 18284
rect 41144 18232 41196 18284
rect 46112 18300 46164 18352
rect 47492 18300 47544 18352
rect 43720 18275 43772 18284
rect 43720 18241 43729 18275
rect 43729 18241 43763 18275
rect 43763 18241 43772 18275
rect 43720 18232 43772 18241
rect 44364 18232 44416 18284
rect 46756 18232 46808 18284
rect 41604 18139 41656 18148
rect 41604 18105 41613 18139
rect 41613 18105 41647 18139
rect 41647 18105 41656 18139
rect 41604 18096 41656 18105
rect 32220 18071 32272 18080
rect 32220 18037 32229 18071
rect 32229 18037 32263 18071
rect 32263 18037 32272 18071
rect 32220 18028 32272 18037
rect 32404 18028 32456 18080
rect 45652 18207 45704 18216
rect 44364 18096 44416 18148
rect 45652 18173 45661 18207
rect 45661 18173 45695 18207
rect 45695 18173 45704 18207
rect 45652 18164 45704 18173
rect 46388 18028 46440 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3056 17824 3108 17876
rect 12440 17824 12492 17876
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 17684 17824 17736 17876
rect 18604 17867 18656 17876
rect 18604 17833 18613 17867
rect 18613 17833 18647 17867
rect 18647 17833 18656 17867
rect 18604 17824 18656 17833
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 23112 17824 23164 17876
rect 29920 17824 29972 17876
rect 12808 17756 12860 17808
rect 15108 17756 15160 17808
rect 24032 17756 24084 17808
rect 42616 17824 42668 17876
rect 44180 17824 44232 17876
rect 36544 17756 36596 17808
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 13728 17620 13780 17672
rect 16672 17688 16724 17740
rect 18696 17688 18748 17740
rect 15660 17620 15712 17672
rect 16580 17620 16632 17672
rect 17500 17620 17552 17672
rect 19156 17620 19208 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 20444 17620 20496 17672
rect 27804 17620 27856 17672
rect 38752 17688 38804 17740
rect 41420 17731 41472 17740
rect 41420 17697 41429 17731
rect 41429 17697 41463 17731
rect 41463 17697 41472 17731
rect 41604 17731 41656 17740
rect 41420 17688 41472 17697
rect 41604 17697 41613 17731
rect 41613 17697 41647 17731
rect 41647 17697 41656 17731
rect 41604 17688 41656 17697
rect 41880 17731 41932 17740
rect 41880 17697 41889 17731
rect 41889 17697 41923 17731
rect 41923 17697 41932 17731
rect 41880 17688 41932 17697
rect 11888 17595 11940 17604
rect 11888 17561 11897 17595
rect 11897 17561 11931 17595
rect 11931 17561 11940 17595
rect 11888 17552 11940 17561
rect 23204 17552 23256 17604
rect 23848 17552 23900 17604
rect 27344 17552 27396 17604
rect 27712 17552 27764 17604
rect 28080 17595 28132 17604
rect 28080 17561 28089 17595
rect 28089 17561 28123 17595
rect 28123 17561 28132 17595
rect 28080 17552 28132 17561
rect 28448 17595 28500 17604
rect 28448 17561 28457 17595
rect 28457 17561 28491 17595
rect 28491 17561 28500 17595
rect 28448 17552 28500 17561
rect 17316 17484 17368 17536
rect 20168 17484 20220 17536
rect 20812 17484 20864 17536
rect 23480 17527 23532 17536
rect 23480 17493 23489 17527
rect 23489 17493 23523 17527
rect 23523 17493 23532 17527
rect 23480 17484 23532 17493
rect 27896 17484 27948 17536
rect 28172 17527 28224 17536
rect 28172 17493 28181 17527
rect 28181 17493 28215 17527
rect 28215 17493 28224 17527
rect 28172 17484 28224 17493
rect 28264 17527 28316 17536
rect 28264 17493 28273 17527
rect 28273 17493 28307 17527
rect 28307 17493 28316 17527
rect 31024 17663 31076 17672
rect 31024 17629 31033 17663
rect 31033 17629 31067 17663
rect 31067 17629 31076 17663
rect 31024 17620 31076 17629
rect 45192 17688 45244 17740
rect 47492 17688 47544 17740
rect 45376 17663 45428 17672
rect 45376 17629 45385 17663
rect 45385 17629 45419 17663
rect 45419 17629 45428 17663
rect 45376 17620 45428 17629
rect 32404 17552 32456 17604
rect 32864 17595 32916 17604
rect 32864 17561 32873 17595
rect 32873 17561 32907 17595
rect 32907 17561 32916 17595
rect 32864 17552 32916 17561
rect 47676 17552 47728 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 28264 17484 28316 17493
rect 43720 17484 43772 17536
rect 44272 17484 44324 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4712 17280 4764 17332
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 14004 17255 14056 17264
rect 14004 17221 14013 17255
rect 14013 17221 14047 17255
rect 14047 17221 14056 17255
rect 14004 17212 14056 17221
rect 19432 17212 19484 17264
rect 20352 17255 20404 17264
rect 20352 17221 20361 17255
rect 20361 17221 20395 17255
rect 20395 17221 20404 17255
rect 20352 17212 20404 17221
rect 20720 17212 20772 17264
rect 20996 17212 21048 17264
rect 22560 17212 22612 17264
rect 28264 17280 28316 17332
rect 29736 17280 29788 17332
rect 36544 17280 36596 17332
rect 28448 17212 28500 17264
rect 32864 17212 32916 17264
rect 41880 17212 41932 17264
rect 44272 17255 44324 17264
rect 44272 17221 44281 17255
rect 44281 17221 44315 17255
rect 44315 17221 44324 17255
rect 44272 17212 44324 17221
rect 45376 17280 45428 17332
rect 47676 17323 47728 17332
rect 47676 17289 47685 17323
rect 47685 17289 47719 17323
rect 47719 17289 47728 17323
rect 47676 17280 47728 17289
rect 45652 17212 45704 17264
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 15660 17144 15712 17196
rect 15936 17144 15988 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 24676 17144 24728 17196
rect 26424 17144 26476 17196
rect 27068 17187 27120 17196
rect 27068 17153 27077 17187
rect 27077 17153 27111 17187
rect 27111 17153 27120 17187
rect 27068 17144 27120 17153
rect 27160 17144 27212 17196
rect 27988 17187 28040 17196
rect 27988 17153 27997 17187
rect 27997 17153 28031 17187
rect 28031 17153 28040 17187
rect 27988 17144 28040 17153
rect 28080 17187 28132 17196
rect 28080 17153 28089 17187
rect 28089 17153 28123 17187
rect 28123 17153 28132 17187
rect 28080 17144 28132 17153
rect 29184 17187 29236 17196
rect 29184 17153 29193 17187
rect 29193 17153 29227 17187
rect 29227 17153 29236 17187
rect 29184 17144 29236 17153
rect 46756 17187 46808 17196
rect 46756 17153 46765 17187
rect 46765 17153 46799 17187
rect 46799 17153 46808 17187
rect 46756 17144 46808 17153
rect 47400 17144 47452 17196
rect 47676 17144 47728 17196
rect 18512 17076 18564 17128
rect 18788 17076 18840 17128
rect 21824 17119 21876 17128
rect 19524 17008 19576 17060
rect 20352 17008 20404 17060
rect 21824 17085 21833 17119
rect 21833 17085 21867 17119
rect 21867 17085 21876 17119
rect 21824 17076 21876 17085
rect 22100 17119 22152 17128
rect 22100 17085 22109 17119
rect 22109 17085 22143 17119
rect 22143 17085 22152 17119
rect 22100 17076 22152 17085
rect 44364 17076 44416 17128
rect 44548 17119 44600 17128
rect 44548 17085 44557 17119
rect 44557 17085 44591 17119
rect 44591 17085 44600 17119
rect 44548 17076 44600 17085
rect 1400 16940 1452 16992
rect 15844 16940 15896 16992
rect 19708 16940 19760 16992
rect 20536 16983 20588 16992
rect 20536 16949 20545 16983
rect 20545 16949 20579 16983
rect 20579 16949 20588 16983
rect 20536 16940 20588 16949
rect 23572 16983 23624 16992
rect 23572 16949 23581 16983
rect 23581 16949 23615 16983
rect 23615 16949 23624 16983
rect 23572 16940 23624 16949
rect 24400 16940 24452 16992
rect 25228 16983 25280 16992
rect 25228 16949 25237 16983
rect 25237 16949 25271 16983
rect 25271 16949 25280 16983
rect 25228 16940 25280 16949
rect 26056 16983 26108 16992
rect 26056 16949 26065 16983
rect 26065 16949 26099 16983
rect 26099 16949 26108 16983
rect 26056 16940 26108 16949
rect 41420 16940 41472 16992
rect 42248 16940 42300 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 18512 16779 18564 16788
rect 18512 16745 18521 16779
rect 18521 16745 18555 16779
rect 18555 16745 18564 16779
rect 18512 16736 18564 16745
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 17316 16668 17368 16720
rect 17408 16668 17460 16720
rect 22100 16736 22152 16788
rect 44548 16736 44600 16788
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 27344 16668 27396 16720
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 20996 16600 21048 16652
rect 24400 16643 24452 16652
rect 20352 16532 20404 16584
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 25412 16600 25464 16652
rect 26148 16643 26200 16652
rect 26148 16609 26157 16643
rect 26157 16609 26191 16643
rect 26191 16609 26200 16643
rect 26148 16600 26200 16609
rect 26424 16600 26476 16652
rect 27988 16668 28040 16720
rect 23480 16532 23532 16584
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 23572 16532 23624 16541
rect 27804 16575 27856 16584
rect 27804 16541 27813 16575
rect 27813 16541 27847 16575
rect 27847 16541 27856 16575
rect 28264 16600 28316 16652
rect 38660 16668 38712 16720
rect 39120 16668 39172 16720
rect 45008 16668 45060 16720
rect 46940 16668 46992 16720
rect 42616 16643 42668 16652
rect 42616 16609 42625 16643
rect 42625 16609 42659 16643
rect 42659 16609 42668 16643
rect 42616 16600 42668 16609
rect 47768 16600 47820 16652
rect 27804 16532 27856 16541
rect 2136 16464 2188 16516
rect 17500 16507 17552 16516
rect 17500 16473 17509 16507
rect 17509 16473 17543 16507
rect 17543 16473 17552 16507
rect 17500 16464 17552 16473
rect 19524 16507 19576 16516
rect 19524 16473 19533 16507
rect 19533 16473 19567 16507
rect 19567 16473 19576 16507
rect 19524 16464 19576 16473
rect 20812 16507 20864 16516
rect 20812 16473 20821 16507
rect 20821 16473 20855 16507
rect 20855 16473 20864 16507
rect 20812 16464 20864 16473
rect 26056 16464 26108 16516
rect 26700 16439 26752 16448
rect 26700 16405 26709 16439
rect 26709 16405 26743 16439
rect 26743 16405 26752 16439
rect 26700 16396 26752 16405
rect 28172 16396 28224 16448
rect 30564 16396 30616 16448
rect 42892 16464 42944 16516
rect 46020 16464 46072 16516
rect 46480 16507 46532 16516
rect 46480 16473 46489 16507
rect 46489 16473 46523 16507
rect 46523 16473 46532 16507
rect 46480 16464 46532 16473
rect 48136 16507 48188 16516
rect 48136 16473 48145 16507
rect 48145 16473 48179 16507
rect 48179 16473 48188 16507
rect 48136 16464 48188 16473
rect 43720 16396 43772 16448
rect 44088 16396 44140 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 1952 16056 2004 16108
rect 19432 16192 19484 16244
rect 21824 16192 21876 16244
rect 25412 16192 25464 16244
rect 28080 16192 28132 16244
rect 28540 16235 28592 16244
rect 28540 16201 28549 16235
rect 28549 16201 28583 16235
rect 28583 16201 28592 16235
rect 28540 16192 28592 16201
rect 42892 16235 42944 16244
rect 42892 16201 42901 16235
rect 42901 16201 42935 16235
rect 42935 16201 42944 16235
rect 42892 16192 42944 16201
rect 43720 16192 43772 16244
rect 45652 16192 45704 16244
rect 20904 16124 20956 16176
rect 28172 16124 28224 16176
rect 44088 16167 44140 16176
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 19156 16056 19208 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 16672 16031 16724 16040
rect 16672 15997 16681 16031
rect 16681 15997 16715 16031
rect 16715 15997 16724 16031
rect 16672 15988 16724 15997
rect 3240 15920 3292 15972
rect 23388 15988 23440 16040
rect 24308 16031 24360 16040
rect 24308 15997 24317 16031
rect 24317 15997 24351 16031
rect 24351 15997 24360 16031
rect 24308 15988 24360 15997
rect 25136 16031 25188 16040
rect 25136 15997 25145 16031
rect 25145 15997 25179 16031
rect 25179 15997 25188 16031
rect 25136 15988 25188 15997
rect 23204 15920 23256 15972
rect 26148 16056 26200 16108
rect 27068 16099 27120 16108
rect 27068 16065 27077 16099
rect 27077 16065 27111 16099
rect 27111 16065 27120 16099
rect 27068 16056 27120 16065
rect 27160 16056 27212 16108
rect 27896 16056 27948 16108
rect 44088 16133 44097 16167
rect 44097 16133 44131 16167
rect 44131 16133 44140 16167
rect 44088 16124 44140 16133
rect 38660 16056 38712 16108
rect 47768 16099 47820 16108
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 42248 15988 42300 16040
rect 45100 16031 45152 16040
rect 45100 15997 45109 16031
rect 45109 15997 45143 16031
rect 45143 15997 45152 16031
rect 45100 15988 45152 15997
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 22560 15648 22612 15700
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 23296 15648 23348 15700
rect 25136 15648 25188 15700
rect 47492 15648 47544 15700
rect 25228 15512 25280 15564
rect 30564 15555 30616 15564
rect 30564 15521 30573 15555
rect 30573 15521 30607 15555
rect 30607 15521 30616 15555
rect 30564 15512 30616 15521
rect 1768 15444 1820 15496
rect 19156 15444 19208 15496
rect 23848 15444 23900 15496
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 26700 15444 26752 15496
rect 16672 15376 16724 15428
rect 23572 15376 23624 15428
rect 25596 15419 25648 15428
rect 25596 15385 25605 15419
rect 25605 15385 25639 15419
rect 25639 15385 25648 15419
rect 25596 15376 25648 15385
rect 32220 15419 32272 15428
rect 32220 15385 32229 15419
rect 32229 15385 32263 15419
rect 32263 15385 32272 15419
rect 32220 15376 32272 15385
rect 23112 15308 23164 15360
rect 24584 15308 24636 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 23388 15147 23440 15156
rect 23388 15113 23397 15147
rect 23397 15113 23431 15147
rect 23431 15113 23440 15147
rect 23388 15104 23440 15113
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 23020 14968 23072 15020
rect 24584 14968 24636 15020
rect 2320 14900 2372 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 23848 14900 23900 14952
rect 25596 14900 25648 14952
rect 22744 14832 22796 14884
rect 23020 14832 23072 14884
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 2688 14356 2740 14408
rect 25780 14356 25832 14408
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 3424 13744 3476 13796
rect 15292 13744 15344 13796
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 22836 13336 22888 13388
rect 23664 13379 23716 13388
rect 23664 13345 23673 13379
rect 23673 13345 23707 13379
rect 23707 13345 23716 13379
rect 23664 13336 23716 13345
rect 47676 13311 47728 13320
rect 47676 13277 47685 13311
rect 47685 13277 47719 13311
rect 47719 13277 47728 13311
rect 47676 13268 47728 13277
rect 22468 13200 22520 13252
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 22468 12971 22520 12980
rect 22468 12937 22477 12971
rect 22477 12937 22511 12971
rect 22511 12937 22520 12971
rect 22468 12928 22520 12937
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 22376 12835 22428 12844
rect 22376 12801 22385 12835
rect 22385 12801 22419 12835
rect 22419 12801 22428 12835
rect 22376 12792 22428 12801
rect 47308 12792 47360 12844
rect 30012 12656 30064 12708
rect 47768 12631 47820 12640
rect 47768 12597 47777 12631
rect 47777 12597 47811 12631
rect 47811 12597 47820 12631
rect 47768 12588 47820 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 47676 12248 47728 12300
rect 48136 12291 48188 12300
rect 48136 12257 48145 12291
rect 48145 12257 48179 12291
rect 48179 12257 48188 12291
rect 48136 12248 48188 12257
rect 47676 12112 47728 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 47676 11883 47728 11892
rect 47676 11849 47685 11883
rect 47685 11849 47719 11883
rect 47719 11849 47728 11883
rect 47676 11840 47728 11849
rect 41512 11704 41564 11756
rect 46940 11704 46992 11756
rect 46480 11500 46532 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 47768 11228 47820 11280
rect 46480 11203 46532 11212
rect 46480 11169 46489 11203
rect 46489 11169 46523 11203
rect 46523 11169 46532 11203
rect 46480 11160 46532 11169
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 4068 10956 4120 11008
rect 12440 10956 12492 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 47492 10616 47544 10668
rect 46296 10412 46348 10464
rect 47676 10455 47728 10464
rect 47676 10421 47685 10455
rect 47685 10421 47719 10455
rect 47719 10421 47728 10455
rect 47676 10412 47728 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 47676 10072 47728 10124
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 48228 9392 48280 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47768 8891 47820 8900
rect 47768 8857 47777 8891
rect 47777 8857 47811 8891
rect 47811 8857 47820 8891
rect 47768 8848 47820 8857
rect 27528 8780 27580 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 48136 8483 48188 8492
rect 48136 8449 48145 8483
rect 48145 8449 48179 8483
rect 48179 8449 48188 8483
rect 48136 8440 48188 8449
rect 47124 8236 47176 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 45560 7939 45612 7948
rect 45560 7905 45569 7939
rect 45569 7905 45603 7939
rect 45603 7905 45612 7939
rect 45560 7896 45612 7905
rect 46756 7896 46808 7948
rect 47124 7939 47176 7948
rect 47124 7905 47133 7939
rect 47133 7905 47167 7939
rect 47167 7905 47176 7939
rect 47124 7896 47176 7905
rect 47584 7760 47636 7812
rect 46296 7692 46348 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 47584 7531 47636 7540
rect 47584 7497 47593 7531
rect 47593 7497 47627 7531
rect 47627 7497 47636 7531
rect 47584 7488 47636 7497
rect 46296 7395 46348 7404
rect 46296 7361 46305 7395
rect 46305 7361 46339 7395
rect 46339 7361 46348 7395
rect 46296 7352 46348 7361
rect 2044 7216 2096 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4068 6808 4120 6860
rect 17500 6808 17552 6860
rect 43536 6808 43588 6860
rect 47308 6851 47360 6860
rect 47308 6817 47317 6851
rect 47317 6817 47351 6851
rect 47351 6817 47360 6851
rect 47308 6808 47360 6817
rect 47400 6808 47452 6860
rect 3976 6672 4028 6724
rect 40868 6715 40920 6724
rect 40868 6681 40877 6715
rect 40877 6681 40911 6715
rect 40911 6681 40920 6715
rect 40868 6672 40920 6681
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 40868 6400 40920 6452
rect 44640 6400 44692 6452
rect 40868 6307 40920 6316
rect 40868 6273 40877 6307
rect 40877 6273 40911 6307
rect 40911 6273 40920 6307
rect 40868 6264 40920 6273
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 45560 5788 45612 5840
rect 41880 5763 41932 5772
rect 41880 5729 41889 5763
rect 41889 5729 41923 5763
rect 41923 5729 41932 5763
rect 41880 5720 41932 5729
rect 43536 5720 43588 5772
rect 41972 5627 42024 5636
rect 41972 5593 41981 5627
rect 41981 5593 42015 5627
rect 42015 5593 42024 5627
rect 41972 5584 42024 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 40868 5312 40920 5364
rect 22100 5176 22152 5228
rect 23848 5176 23900 5228
rect 41972 5176 42024 5228
rect 47768 5219 47820 5228
rect 47768 5185 47777 5219
rect 47777 5185 47811 5219
rect 47811 5185 47820 5219
rect 47768 5176 47820 5185
rect 19064 5108 19116 5160
rect 32036 5108 32088 5160
rect 23112 5040 23164 5092
rect 22284 4972 22336 5024
rect 22928 4972 22980 5024
rect 40316 5015 40368 5024
rect 40316 4981 40325 5015
rect 40325 4981 40359 5015
rect 40359 4981 40368 5015
rect 40316 4972 40368 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19340 4768 19392 4820
rect 32312 4768 32364 4820
rect 22376 4700 22428 4752
rect 31760 4700 31812 4752
rect 40316 4700 40368 4752
rect 22100 4675 22152 4684
rect 22100 4641 22109 4675
rect 22109 4641 22143 4675
rect 22143 4641 22152 4675
rect 22100 4632 22152 4641
rect 23756 4632 23808 4684
rect 38568 4632 38620 4684
rect 46296 4632 46348 4684
rect 21088 4564 21140 4616
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 22376 4564 22428 4616
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23480 4607 23532 4616
rect 23480 4573 23489 4607
rect 23489 4573 23523 4607
rect 23523 4573 23532 4607
rect 23480 4564 23532 4573
rect 40500 4564 40552 4616
rect 6644 4496 6696 4548
rect 37004 4539 37056 4548
rect 37004 4505 37013 4539
rect 37013 4505 37047 4539
rect 37047 4505 37056 4539
rect 37004 4496 37056 4505
rect 38660 4496 38712 4548
rect 46848 4564 46900 4616
rect 47492 4496 47544 4548
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 20812 4471 20864 4480
rect 20812 4437 20821 4471
rect 20821 4437 20855 4471
rect 20855 4437 20864 4471
rect 20812 4428 20864 4437
rect 22468 4428 22520 4480
rect 25320 4428 25372 4480
rect 40040 4471 40092 4480
rect 40040 4437 40049 4471
rect 40049 4437 40083 4471
rect 40083 4437 40092 4471
rect 40040 4428 40092 4437
rect 40132 4428 40184 4480
rect 46756 4471 46808 4480
rect 46756 4437 46765 4471
rect 46765 4437 46799 4471
rect 46799 4437 46808 4471
rect 46756 4428 46808 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 13452 4088 13504 4140
rect 13544 4088 13596 4140
rect 17224 4088 17276 4140
rect 17592 4088 17644 4140
rect 18328 4131 18380 4140
rect 18328 4097 18337 4131
rect 18337 4097 18371 4131
rect 18371 4097 18380 4131
rect 18328 4088 18380 4097
rect 8300 4020 8352 4072
rect 1584 3884 1636 3936
rect 2780 3884 2832 3936
rect 7104 3884 7156 3936
rect 9128 4020 9180 4072
rect 17316 4020 17368 4072
rect 20904 4224 20956 4276
rect 21364 4224 21416 4276
rect 22652 4224 22704 4276
rect 20168 4156 20220 4208
rect 19340 4088 19392 4140
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 20352 4088 20404 4140
rect 20168 4020 20220 4072
rect 20812 4088 20864 4140
rect 22100 4088 22152 4140
rect 22468 4131 22520 4140
rect 22468 4097 22477 4131
rect 22477 4097 22511 4131
rect 22511 4097 22520 4131
rect 22468 4088 22520 4097
rect 22744 4156 22796 4208
rect 23112 4131 23164 4140
rect 21272 4020 21324 4072
rect 21364 4020 21416 4072
rect 9220 3884 9272 3936
rect 9956 3884 10008 3936
rect 18236 3952 18288 4004
rect 18788 3952 18840 4004
rect 22008 3952 22060 4004
rect 22376 4020 22428 4072
rect 23112 4097 23121 4131
rect 23121 4097 23155 4131
rect 23155 4097 23164 4131
rect 23112 4088 23164 4097
rect 23204 4088 23256 4140
rect 23756 4131 23808 4140
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 23756 4088 23808 4097
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 24860 4088 24912 4140
rect 25688 4224 25740 4276
rect 37004 4224 37056 4276
rect 25596 4156 25648 4208
rect 37648 4199 37700 4208
rect 37648 4165 37657 4199
rect 37657 4165 37691 4199
rect 37691 4165 37700 4199
rect 37648 4156 37700 4165
rect 38568 4199 38620 4208
rect 38568 4165 38577 4199
rect 38577 4165 38611 4199
rect 38611 4165 38620 4199
rect 38568 4156 38620 4165
rect 36728 4131 36780 4140
rect 25228 4020 25280 4072
rect 25412 4063 25464 4072
rect 25412 4029 25421 4063
rect 25421 4029 25455 4063
rect 25455 4029 25464 4063
rect 25412 4020 25464 4029
rect 27804 4020 27856 4072
rect 36728 4097 36737 4131
rect 36737 4097 36771 4131
rect 36771 4097 36780 4131
rect 36728 4088 36780 4097
rect 37556 4063 37608 4072
rect 37556 4029 37565 4063
rect 37565 4029 37599 4063
rect 37599 4029 37608 4063
rect 37556 4020 37608 4029
rect 40040 4156 40092 4208
rect 40040 4063 40092 4072
rect 11704 3884 11756 3936
rect 14004 3884 14056 3936
rect 17684 3884 17736 3936
rect 17868 3884 17920 3936
rect 20720 3884 20772 3936
rect 21824 3884 21876 3936
rect 21916 3884 21968 3936
rect 24308 3884 24360 3936
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 25504 3952 25556 4004
rect 40040 4029 40049 4063
rect 40049 4029 40083 4063
rect 40083 4029 40092 4063
rect 40040 4020 40092 4029
rect 40316 4020 40368 4072
rect 40500 4063 40552 4072
rect 40500 4029 40509 4063
rect 40509 4029 40543 4063
rect 40543 4029 40552 4063
rect 40500 4020 40552 4029
rect 46388 4156 46440 4208
rect 46664 4156 46716 4208
rect 44916 4088 44968 4140
rect 27436 3884 27488 3936
rect 27712 3884 27764 3936
rect 39580 3952 39632 4004
rect 39764 3952 39816 4004
rect 38476 3884 38528 3936
rect 42800 3884 42852 3936
rect 43812 3927 43864 3936
rect 43812 3893 43821 3927
rect 43821 3893 43855 3927
rect 43855 3893 43864 3927
rect 43812 3884 43864 3893
rect 46296 3884 46348 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 17316 3680 17368 3732
rect 22744 3680 22796 3732
rect 1860 3544 1912 3596
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 7288 3476 7340 3528
rect 22928 3612 22980 3664
rect 23204 3680 23256 3732
rect 24860 3612 24912 3664
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9220 3544 9272 3553
rect 9404 3544 9456 3596
rect 12348 3544 12400 3596
rect 9128 3476 9180 3528
rect 11520 3476 11572 3528
rect 13820 3476 13872 3528
rect 16396 3544 16448 3596
rect 20996 3544 21048 3596
rect 21088 3544 21140 3596
rect 22008 3544 22060 3596
rect 32864 3680 32916 3732
rect 1308 3408 1360 3460
rect 2044 3340 2096 3392
rect 6920 3340 6972 3392
rect 10140 3408 10192 3460
rect 16764 3476 16816 3528
rect 17684 3476 17736 3528
rect 17960 3476 18012 3528
rect 18604 3476 18656 3528
rect 19432 3476 19484 3528
rect 18788 3408 18840 3460
rect 20720 3476 20772 3528
rect 21456 3476 21508 3528
rect 21824 3519 21876 3528
rect 21824 3485 21833 3519
rect 21833 3485 21867 3519
rect 21867 3485 21876 3519
rect 21824 3476 21876 3485
rect 23848 3519 23900 3528
rect 23848 3485 23857 3519
rect 23857 3485 23891 3519
rect 23891 3485 23900 3519
rect 23848 3476 23900 3485
rect 25228 3544 25280 3596
rect 29736 3544 29788 3596
rect 27252 3519 27304 3528
rect 27252 3485 27261 3519
rect 27261 3485 27295 3519
rect 27295 3485 27304 3519
rect 27252 3476 27304 3485
rect 30932 3612 30984 3664
rect 32220 3612 32272 3664
rect 31484 3519 31536 3528
rect 31484 3485 31493 3519
rect 31493 3485 31527 3519
rect 31527 3485 31536 3519
rect 31484 3476 31536 3485
rect 32220 3476 32272 3528
rect 24492 3408 24544 3460
rect 25320 3408 25372 3460
rect 16396 3340 16448 3392
rect 16672 3340 16724 3392
rect 17776 3340 17828 3392
rect 18512 3340 18564 3392
rect 19984 3340 20036 3392
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 20720 3340 20772 3392
rect 22836 3340 22888 3392
rect 27804 3408 27856 3460
rect 38660 3680 38712 3732
rect 39396 3680 39448 3732
rect 40316 3612 40368 3664
rect 40592 3612 40644 3664
rect 37556 3544 37608 3596
rect 38476 3519 38528 3528
rect 38476 3485 38485 3519
rect 38485 3485 38519 3519
rect 38519 3485 38528 3519
rect 38476 3476 38528 3485
rect 39304 3519 39356 3528
rect 39304 3485 39313 3519
rect 39313 3485 39347 3519
rect 39347 3485 39356 3519
rect 39304 3476 39356 3485
rect 41880 3544 41932 3596
rect 43812 3612 43864 3664
rect 42800 3587 42852 3596
rect 42800 3553 42809 3587
rect 42809 3553 42843 3587
rect 42843 3553 42852 3587
rect 42800 3544 42852 3553
rect 43168 3587 43220 3596
rect 43168 3553 43177 3587
rect 43177 3553 43211 3587
rect 43211 3553 43220 3587
rect 43168 3544 43220 3553
rect 39948 3476 40000 3528
rect 41788 3476 41840 3528
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 40500 3408 40552 3460
rect 42524 3408 42576 3460
rect 43996 3408 44048 3460
rect 48964 3408 49016 3460
rect 27436 3340 27488 3392
rect 31116 3340 31168 3392
rect 32404 3340 32456 3392
rect 37648 3340 37700 3392
rect 41420 3340 41472 3392
rect 42432 3340 42484 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4068 3136 4120 3188
rect 9956 3136 10008 3188
rect 16764 3179 16816 3188
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 7472 3111 7524 3120
rect 7472 3077 7481 3111
rect 7481 3077 7515 3111
rect 7515 3077 7524 3111
rect 7472 3068 7524 3077
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 10140 3111 10192 3120
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 11704 3111 11756 3120
rect 10140 3068 10192 3077
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 14004 3111 14056 3120
rect 14004 3077 14013 3111
rect 14013 3077 14047 3111
rect 14047 3077 14056 3111
rect 14004 3068 14056 3077
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 17960 3179 18012 3188
rect 17960 3145 17969 3179
rect 17969 3145 18003 3179
rect 18003 3145 18012 3179
rect 17960 3136 18012 3145
rect 18604 3179 18656 3188
rect 18604 3145 18613 3179
rect 18613 3145 18647 3179
rect 18647 3145 18656 3179
rect 18604 3136 18656 3145
rect 20720 3136 20772 3188
rect 20812 3136 20864 3188
rect 20628 3068 20680 3120
rect 22192 3136 22244 3188
rect 22560 3068 22612 3120
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 17868 3043 17920 3052
rect 17868 3009 17877 3043
rect 17877 3009 17911 3043
rect 17911 3009 17920 3043
rect 17868 3000 17920 3009
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 21916 3000 21968 3052
rect 664 2932 716 2984
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 10968 2864 11020 2916
rect 14188 2932 14240 2984
rect 14832 2932 14884 2984
rect 19708 2932 19760 2984
rect 19892 2975 19944 2984
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 19984 2932 20036 2984
rect 20168 2932 20220 2984
rect 20352 2932 20404 2984
rect 25596 3068 25648 3120
rect 27252 3136 27304 3188
rect 27344 3136 27396 3188
rect 36728 3179 36780 3188
rect 36728 3145 36737 3179
rect 36737 3145 36771 3179
rect 36771 3145 36780 3179
rect 36728 3136 36780 3145
rect 39304 3136 39356 3188
rect 40408 3136 40460 3188
rect 22836 3043 22888 3052
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 27712 3068 27764 3120
rect 25780 3000 25832 3052
rect 26240 3000 26292 3052
rect 27068 3000 27120 3052
rect 23572 2975 23624 2984
rect 3884 2796 3936 2848
rect 22192 2864 22244 2916
rect 22376 2907 22428 2916
rect 22376 2873 22385 2907
rect 22385 2873 22419 2907
rect 22419 2873 22428 2907
rect 22376 2864 22428 2873
rect 23572 2941 23581 2975
rect 23581 2941 23615 2975
rect 23615 2941 23624 2975
rect 23572 2932 23624 2941
rect 27620 2932 27672 2984
rect 26240 2864 26292 2916
rect 32128 3068 32180 3120
rect 32404 3111 32456 3120
rect 32404 3077 32413 3111
rect 32413 3077 32447 3111
rect 32447 3077 32456 3111
rect 32404 3068 32456 3077
rect 47032 3136 47084 3188
rect 41696 3068 41748 3120
rect 44456 3068 44508 3120
rect 46756 3068 46808 3120
rect 32220 3043 32272 3052
rect 32220 3009 32229 3043
rect 32229 3009 32263 3043
rect 32263 3009 32272 3043
rect 32220 3000 32272 3009
rect 37648 3000 37700 3052
rect 39120 3000 39172 3052
rect 39948 3000 40000 3052
rect 41512 3000 41564 3052
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 48320 3000 48372 3052
rect 33508 2864 33560 2916
rect 13452 2796 13504 2848
rect 20812 2796 20864 2848
rect 20904 2796 20956 2848
rect 22100 2796 22152 2848
rect 25780 2839 25832 2848
rect 25780 2805 25789 2839
rect 25789 2805 25823 2839
rect 25823 2805 25832 2839
rect 25780 2796 25832 2805
rect 26148 2796 26200 2848
rect 41788 2932 41840 2984
rect 36176 2796 36228 2848
rect 40408 2796 40460 2848
rect 40592 2796 40644 2848
rect 47676 2932 47728 2984
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2780 2524 2832 2576
rect 6644 2524 6696 2576
rect 9588 2592 9640 2644
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 6460 2456 6512 2508
rect 6920 2456 6972 2508
rect 12348 2524 12400 2576
rect 16488 2524 16540 2576
rect 17592 2592 17644 2644
rect 18328 2592 18380 2644
rect 19708 2592 19760 2644
rect 20076 2592 20128 2644
rect 20260 2592 20312 2644
rect 23664 2592 23716 2644
rect 26056 2592 26108 2644
rect 31760 2592 31812 2644
rect 32128 2592 32180 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 39120 2635 39172 2644
rect 39120 2601 39129 2635
rect 39129 2601 39163 2635
rect 39163 2601 39172 2635
rect 39120 2592 39172 2601
rect 41788 2592 41840 2644
rect 11704 2456 11756 2508
rect 25412 2524 25464 2576
rect 28908 2524 28960 2576
rect 22284 2456 22336 2508
rect 2596 2320 2648 2372
rect 5172 2388 5224 2440
rect 15016 2388 15068 2440
rect 15476 2388 15528 2440
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 17776 2431 17828 2440
rect 15568 2388 15620 2397
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 18236 2388 18288 2440
rect 19800 2388 19852 2440
rect 20076 2388 20128 2440
rect 22376 2431 22428 2440
rect 22376 2397 22385 2431
rect 22385 2397 22419 2431
rect 22419 2397 22428 2431
rect 22376 2388 22428 2397
rect 23848 2456 23900 2508
rect 24676 2499 24728 2508
rect 24676 2465 24685 2499
rect 24685 2465 24719 2499
rect 24719 2465 24728 2499
rect 24676 2456 24728 2465
rect 25136 2499 25188 2508
rect 25136 2465 25145 2499
rect 25145 2465 25179 2499
rect 25179 2465 25188 2499
rect 25136 2456 25188 2465
rect 27160 2456 27212 2508
rect 33140 2456 33192 2508
rect 41972 2456 42024 2508
rect 46572 2456 46624 2508
rect 26424 2388 26476 2440
rect 28356 2388 28408 2440
rect 29644 2388 29696 2440
rect 35440 2388 35492 2440
rect 38016 2388 38068 2440
rect 39948 2388 40000 2440
rect 41236 2388 41288 2440
rect 43812 2388 43864 2440
rect 8392 2320 8444 2372
rect 16120 2320 16172 2372
rect 20628 2320 20680 2372
rect 36084 2320 36136 2372
rect 39396 2320 39448 2372
rect 40592 2320 40644 2372
rect 41420 2320 41472 2372
rect 47032 2388 47084 2440
rect 48044 2388 48096 2440
rect 46756 2320 46808 2372
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 31852 2252 31904 2304
rect 43260 2252 43312 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3516 2048 3568 2100
rect 9588 2048 9640 2100
rect 9680 2048 9732 2100
rect 23940 2048 23992 2100
rect 2964 1980 3016 2032
rect 11704 1980 11756 2032
rect 15568 1980 15620 2032
rect 36176 1980 36228 2032
rect 22560 1368 22612 1420
rect 23572 1368 23624 1420
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4844 49314
rect 4498 49200 4610 49286
rect 32 22098 60 49200
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 46578 1440 47631
rect 1964 47054 1992 49200
rect 2044 47456 2096 47462
rect 2044 47398 2096 47404
rect 2056 47122 2084 47398
rect 2044 47116 2096 47122
rect 2044 47058 2096 47064
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2608 46918 2636 49200
rect 3056 47524 3108 47530
rect 3056 47466 3108 47472
rect 3068 47258 3096 47466
rect 3056 47252 3108 47258
rect 3056 47194 3108 47200
rect 3252 47054 3280 49200
rect 3332 47252 3384 47258
rect 3332 47194 3384 47200
rect 3240 47048 3292 47054
rect 3344 47025 3372 47194
rect 3240 46990 3292 46996
rect 3330 47016 3386 47025
rect 3330 46951 3386 46960
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 3896 46646 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4816 47054 4844 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7420 49314
rect 7074 49200 7186 49286
rect 5828 47054 5856 49200
rect 7392 47054 7420 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7380 47048 7432 47054
rect 7380 46990 7432 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 6644 46980 6696 46986
rect 6644 46922 6696 46928
rect 7472 46980 7524 46986
rect 7472 46922 7524 46928
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 1676 46368 1728 46374
rect 1676 46310 1728 46316
rect 2778 46336 2834 46345
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35465 1624 35634
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1584 33992 1636 33998
rect 1584 33934 1636 33940
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1596 32745 1624 33934
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1688 29238 1716 46310
rect 2778 46271 2834 46280
rect 1768 45960 1820 45966
rect 1768 45902 1820 45908
rect 1780 45490 1808 45902
rect 1768 45484 1820 45490
rect 1768 45426 1820 45432
rect 2792 45422 2820 46271
rect 3988 46170 4016 46446
rect 3976 46164 4028 46170
rect 3976 46106 4028 46112
rect 2228 45416 2280 45422
rect 2228 45358 2280 45364
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 2240 45082 2268 45358
rect 2228 45076 2280 45082
rect 2228 45018 2280 45024
rect 3422 44976 3478 44985
rect 3422 44911 3478 44920
rect 2320 44872 2372 44878
rect 2320 44814 2372 44820
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 2332 37942 2360 44814
rect 2320 37936 2372 37942
rect 2320 37878 2372 37884
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2136 36168 2188 36174
rect 2136 36110 2188 36116
rect 2044 35488 2096 35494
rect 2044 35430 2096 35436
rect 1952 33856 2004 33862
rect 1952 33798 2004 33804
rect 1860 33448 1912 33454
rect 1860 33390 1912 33396
rect 1872 32994 1900 33390
rect 1964 33114 1992 33798
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 1872 32966 1992 32994
rect 1964 32910 1992 32966
rect 1952 32904 2004 32910
rect 1952 32846 2004 32852
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1964 31414 1992 32846
rect 2056 32434 2084 35430
rect 2044 32428 2096 32434
rect 2044 32370 2096 32376
rect 1952 31408 2004 31414
rect 1952 31350 2004 31356
rect 1676 29232 1728 29238
rect 1676 29174 1728 29180
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 20 22092 72 22098
rect 20 22034 72 22040
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1872 17785 1900 18226
rect 1858 17776 1914 17785
rect 1858 17711 1914 17720
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1964 6914 1992 16050
rect 2056 7274 2084 25094
rect 2148 18766 2176 36110
rect 2228 32768 2280 32774
rect 2228 32710 2280 32716
rect 2240 32502 2268 32710
rect 2228 32496 2280 32502
rect 2228 32438 2280 32444
rect 2332 31346 2360 37878
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 3330 31376 3386 31385
rect 2320 31340 2372 31346
rect 3330 31311 3386 31320
rect 2320 31282 2372 31288
rect 2872 31272 2924 31278
rect 2872 31214 2924 31220
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2884 16574 2912 31214
rect 3344 29306 3372 31311
rect 3332 29300 3384 29306
rect 3332 29242 3384 29248
rect 3330 28656 3386 28665
rect 3330 28591 3386 28600
rect 3344 27674 3372 28591
rect 3332 27668 3384 27674
rect 3332 27610 3384 27616
rect 3436 21010 3464 44911
rect 3514 43616 3570 43625
rect 3514 43551 3570 43560
rect 3528 21622 3556 43551
rect 3698 39536 3754 39545
rect 3698 39471 3754 39480
rect 3712 21690 3740 39471
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3516 21616 3568 21622
rect 3516 21558 3568 21564
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 3068 19825 3096 20538
rect 3054 19816 3110 19825
rect 3054 19751 3110 19760
rect 3422 18456 3478 18465
rect 3422 18391 3424 18400
rect 3476 18391 3478 18400
rect 3424 18362 3476 18368
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3068 17105 3096 17818
rect 3054 17096 3110 17105
rect 3054 17031 3110 17040
rect 2884 16546 3004 16574
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2332 14618 2360 14894
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1964 6886 2084 6914
rect 2056 4146 2084 6886
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3402
rect 1596 2514 1624 3878
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3058 1900 3538
rect 2700 3534 2728 14350
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 3126 2084 3334
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 2792 2582 2820 3878
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2608 800 2636 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2884 785 2912 2450
rect 2976 2038 3004 16546
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 3252 7585 3280 15914
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 13705 3464 13738
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 4080 12434 4108 46922
rect 5080 46504 5132 46510
rect 5080 46446 5132 46452
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 5092 46170 5120 46446
rect 5080 46164 5132 46170
rect 5080 46106 5132 46112
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4712 32360 4764 32366
rect 4712 32302 4764 32308
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4724 31414 4752 32302
rect 4712 31408 4764 31414
rect 4712 31350 4764 31356
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4724 17338 4752 31350
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3988 12406 4108 12434
rect 3238 7576 3294 7585
rect 3238 7511 3294 7520
rect 3988 6730 4016 12406
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10305 4108 10950
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4066 10296 4122 10305
rect 4214 10288 4522 10308
rect 4066 10231 4122 10240
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 6656 4554 6684 46922
rect 7484 28694 7512 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 7472 28688 7524 28694
rect 7472 28630 7524 28636
rect 8312 26450 8340 45526
rect 9508 37738 9536 46922
rect 10980 46374 11008 49200
rect 11624 47122 11652 49200
rect 11612 47116 11664 47122
rect 11612 47058 11664 47064
rect 12072 46504 12124 46510
rect 12072 46446 12124 46452
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 12084 45626 12112 46446
rect 12268 45966 12296 49200
rect 12912 47054 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49200 16202 50000
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49314 27150 50000
rect 26712 49286 27150 49314
rect 13740 47122 13860 47138
rect 13740 47116 13872 47122
rect 13740 47110 13820 47116
rect 13820 47058 13872 47064
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 14200 46594 14228 49200
rect 14464 47048 14516 47054
rect 14464 46990 14516 46996
rect 14200 46566 14320 46594
rect 14292 46510 14320 46566
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 13556 46170 13584 46446
rect 14200 46170 14228 46446
rect 13544 46164 13596 46170
rect 13544 46106 13596 46112
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 12256 45960 12308 45966
rect 12256 45902 12308 45908
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 12348 45824 12400 45830
rect 12348 45766 12400 45772
rect 12072 45620 12124 45626
rect 12072 45562 12124 45568
rect 11980 45484 12032 45490
rect 11980 45426 12032 45432
rect 10324 40384 10376 40390
rect 10324 40326 10376 40332
rect 9496 37732 9548 37738
rect 9496 37674 9548 37680
rect 10336 34746 10364 40326
rect 11992 38282 12020 45426
rect 12360 38350 12388 45766
rect 14108 41138 14136 45902
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 12348 38344 12400 38350
rect 12348 38286 12400 38292
rect 11980 38276 12032 38282
rect 11980 38218 12032 38224
rect 14476 37806 14504 46990
rect 15488 45554 15516 49200
rect 15936 47592 15988 47598
rect 15936 47534 15988 47540
rect 15488 45526 15792 45554
rect 14464 37800 14516 37806
rect 14370 37768 14426 37777
rect 14464 37742 14516 37748
rect 14370 37703 14372 37712
rect 14424 37703 14426 37712
rect 14372 37674 14424 37680
rect 15568 37256 15620 37262
rect 15568 37198 15620 37204
rect 13912 36712 13964 36718
rect 13912 36654 13964 36660
rect 13924 36106 13952 36654
rect 14924 36236 14976 36242
rect 14924 36178 14976 36184
rect 13912 36100 13964 36106
rect 13912 36042 13964 36048
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 13924 34066 13952 36042
rect 14188 35556 14240 35562
rect 14188 35498 14240 35504
rect 14200 34610 14228 35498
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 13912 33856 13964 33862
rect 13912 33798 13964 33804
rect 13924 33658 13952 33798
rect 14384 33658 14412 33866
rect 13912 33652 13964 33658
rect 13912 33594 13964 33600
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 14568 33522 14596 34342
rect 14936 34066 14964 36178
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15016 34944 15068 34950
rect 15016 34886 15068 34892
rect 15028 34610 15056 34886
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 15108 34604 15160 34610
rect 15108 34546 15160 34552
rect 15016 34196 15068 34202
rect 15016 34138 15068 34144
rect 14924 34060 14976 34066
rect 14924 34002 14976 34008
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 13912 33448 13964 33454
rect 13912 33390 13964 33396
rect 13924 32978 13952 33390
rect 14384 33114 14412 33458
rect 14936 33454 14964 34002
rect 14924 33448 14976 33454
rect 14924 33390 14976 33396
rect 14372 33108 14424 33114
rect 14372 33050 14424 33056
rect 13912 32972 13964 32978
rect 13912 32914 13964 32920
rect 14384 31754 14412 33050
rect 14936 33046 14964 33390
rect 15028 33318 15056 34138
rect 15016 33312 15068 33318
rect 15016 33254 15068 33260
rect 14924 33040 14976 33046
rect 14924 32982 14976 32988
rect 15028 32910 15056 33254
rect 15120 32978 15148 34546
rect 15212 33522 15240 35974
rect 15580 34950 15608 37198
rect 15660 36712 15712 36718
rect 15660 36654 15712 36660
rect 15672 36378 15700 36654
rect 15660 36372 15712 36378
rect 15660 36314 15712 36320
rect 15568 34944 15620 34950
rect 15568 34886 15620 34892
rect 15476 34672 15528 34678
rect 15476 34614 15528 34620
rect 15292 34536 15344 34542
rect 15292 34478 15344 34484
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 14464 32904 14516 32910
rect 14464 32846 14516 32852
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 14476 31890 14504 32846
rect 15212 32026 15240 33458
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 14464 31884 14516 31890
rect 14464 31826 14516 31832
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14372 31748 14424 31754
rect 14372 31690 14424 31696
rect 14384 30802 14412 31690
rect 14372 30796 14424 30802
rect 14372 30738 14424 30744
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14476 30394 14504 30670
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 14568 30258 14596 31826
rect 15304 31754 15332 34478
rect 15488 33998 15516 34614
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 15488 32570 15516 32846
rect 15476 32564 15528 32570
rect 15476 32506 15528 32512
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15304 31726 15424 31754
rect 15108 31272 15160 31278
rect 15108 31214 15160 31220
rect 15120 30938 15148 31214
rect 15108 30932 15160 30938
rect 15108 30874 15160 30880
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 14556 30252 14608 30258
rect 14556 30194 14608 30200
rect 14740 30252 14792 30258
rect 14740 30194 14792 30200
rect 14752 29782 14780 30194
rect 14740 29776 14792 29782
rect 14740 29718 14792 29724
rect 14464 29232 14516 29238
rect 14462 29200 14464 29209
rect 14516 29200 14518 29209
rect 14462 29135 14518 29144
rect 14464 28416 14516 28422
rect 14464 28358 14516 28364
rect 14476 28150 14504 28358
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 12716 28008 12768 28014
rect 12716 27950 12768 27956
rect 12348 26920 12400 26926
rect 12348 26862 12400 26868
rect 12360 26586 12388 26862
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11900 25906 11928 26318
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 11716 25362 11744 25638
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 11900 23730 11928 25842
rect 12452 25838 12480 26250
rect 12636 25974 12664 26794
rect 12728 26382 12756 27950
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 12624 25968 12676 25974
rect 12624 25910 12676 25916
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 13096 25498 13124 26318
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 12452 24954 12480 25434
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 12084 24342 12112 24754
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12072 24336 12124 24342
rect 12072 24278 12124 24284
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11808 23186 11836 23462
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11900 22030 11928 23666
rect 12084 23202 12112 24278
rect 12452 24206 12480 24550
rect 12544 24410 12572 25298
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12636 24750 12664 24890
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12728 24682 12756 25094
rect 13096 24818 13124 25434
rect 13280 25226 13308 26182
rect 13372 25226 13400 26250
rect 13740 25838 13768 26862
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 14188 26308 14240 26314
rect 14188 26250 14240 26256
rect 14200 25974 14228 26250
rect 14844 25974 14872 26318
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 14832 25968 14884 25974
rect 14832 25910 14884 25916
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13268 25220 13320 25226
rect 13268 25162 13320 25168
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 13372 24818 13400 25162
rect 13740 24954 13768 25774
rect 13820 25764 13872 25770
rect 13820 25706 13872 25712
rect 13728 24948 13780 24954
rect 13728 24890 13780 24896
rect 13832 24818 13860 25706
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14936 25362 14964 25638
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 12716 24676 12768 24682
rect 12716 24618 12768 24624
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 11992 23174 12112 23202
rect 11992 22642 12020 23174
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 12084 22574 12112 22986
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 12360 22114 12388 22578
rect 12360 22086 12480 22114
rect 12452 22030 12480 22086
rect 11888 22024 11940 22030
rect 12348 22024 12400 22030
rect 11940 21972 12020 21978
rect 11888 21966 12020 21972
rect 12348 21966 12400 21972
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 11900 21950 12020 21966
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11532 20942 11560 21830
rect 11796 21616 11848 21622
rect 11796 21558 11848 21564
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11716 20806 11744 21422
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11808 18290 11836 21558
rect 11900 20874 11928 21830
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11992 20466 12020 21950
rect 12360 21146 12388 21966
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 12728 18902 12756 24618
rect 13372 24138 13400 24754
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13360 24132 13412 24138
rect 13360 24074 13412 24080
rect 13556 23186 13584 24686
rect 13832 24206 13860 24754
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14476 23594 14504 24074
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14464 23588 14516 23594
rect 14464 23530 14516 23536
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13084 23044 13136 23050
rect 13084 22986 13136 22992
rect 13096 22778 13124 22986
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 13556 22710 13584 23122
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12912 20058 12940 20878
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13004 19854 13032 22578
rect 14844 22098 14872 23666
rect 14924 23044 14976 23050
rect 14924 22986 14976 22992
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14740 22024 14792 22030
rect 14936 21978 14964 22986
rect 14792 21972 14964 21978
rect 14740 21966 14964 21972
rect 14752 21950 14964 21966
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 13636 20528 13688 20534
rect 13636 20470 13688 20476
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19378 13032 19790
rect 13648 19514 13676 20470
rect 14292 20398 14320 21422
rect 14476 21146 14504 21422
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14844 20942 14872 21950
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14108 20058 14136 20334
rect 14292 20058 14320 20334
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14384 19938 14412 20878
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14476 20330 14504 20742
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 14292 19910 14412 19938
rect 14292 19718 14320 19910
rect 14476 19854 14504 20266
rect 14936 20058 14964 20334
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 11888 18692 11940 18698
rect 11888 18634 11940 18640
rect 11900 18358 11928 18634
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11808 17202 11836 18226
rect 12452 17882 12480 18770
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12820 17814 12848 19314
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11900 17338 11928 17546
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 12452 11014 12480 17682
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 6460 3528 6512 3534
rect 4066 3496 4122 3505
rect 6460 3470 6512 3476
rect 4066 3431 4122 3440
rect 4080 3194 4108 3431
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 2964 2032 3016 2038
rect 2964 1974 3016 1980
rect 3528 1465 3556 2042
rect 3514 1456 3570 1465
rect 3514 1391 3570 1400
rect 3896 800 3924 2790
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 6472 2514 6500 3470
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5184 800 5212 2382
rect 6656 1306 6684 2518
rect 6932 2514 6960 3334
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6472 1278 6684 1306
rect 6472 800 6500 1278
rect 7116 800 7144 3878
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7300 3058 7328 3470
rect 7484 3126 7512 4422
rect 13556 4146 13584 18566
rect 13648 18358 13676 19110
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13740 17678 13768 19314
rect 14292 19310 14320 19654
rect 14936 19514 14964 19994
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 14016 17270 14044 18158
rect 14384 17882 14412 18294
rect 14936 18086 14964 19450
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 8312 3738 8340 4014
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 9140 3534 9168 4014
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 9232 3602 9260 3878
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 800 7788 2926
rect 9416 2774 9444 3538
rect 9968 3194 9996 3878
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10152 3126 10180 3402
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 11532 3058 11560 3470
rect 11716 3126 11744 3878
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 9048 2746 9444 2774
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9048 800 9076 2746
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9600 2106 9628 2586
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 2106 9720 2246
rect 9588 2100 9640 2106
rect 9588 2042 9640 2048
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 10980 800 11008 2858
rect 12360 2582 12388 3538
rect 13464 2854 13492 4082
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13832 3058 13860 3470
rect 14016 3126 14044 3878
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11716 2038 11744 2450
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 14200 800 14228 2926
rect 14844 800 14872 2926
rect 15028 2446 15056 30670
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15120 24750 15148 25842
rect 15304 25838 15332 26318
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 15304 25498 15332 25774
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 15120 23594 15148 24686
rect 15212 24410 15240 25162
rect 15304 24682 15332 25434
rect 15292 24676 15344 24682
rect 15292 24618 15344 24624
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15212 22098 15240 22374
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15120 19786 15148 20198
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15120 19446 15148 19722
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 15212 19310 15240 19926
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15212 18358 15240 18702
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15120 17814 15148 18022
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15304 13802 15332 22034
rect 15396 18154 15424 31726
rect 15580 31482 15608 31758
rect 15764 31754 15792 45526
rect 15948 37466 15976 47534
rect 16132 46918 16160 49200
rect 17420 47410 17448 49200
rect 16684 47382 17448 47410
rect 16580 47048 16632 47054
rect 16580 46990 16632 46996
rect 16592 46918 16620 46990
rect 16120 46912 16172 46918
rect 16120 46854 16172 46860
rect 16580 46912 16632 46918
rect 16580 46854 16632 46860
rect 16488 38344 16540 38350
rect 16488 38286 16540 38292
rect 16500 37466 16528 38286
rect 15936 37460 15988 37466
rect 15936 37402 15988 37408
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 15936 37256 15988 37262
rect 15936 37198 15988 37204
rect 16028 37256 16080 37262
rect 16028 37198 16080 37204
rect 15844 37120 15896 37126
rect 15844 37062 15896 37068
rect 15856 36174 15884 37062
rect 15948 36582 15976 37198
rect 15936 36576 15988 36582
rect 15936 36518 15988 36524
rect 15844 36168 15896 36174
rect 15844 36110 15896 36116
rect 16040 34610 16068 37198
rect 16212 36576 16264 36582
rect 16212 36518 16264 36524
rect 16224 36242 16252 36518
rect 16212 36236 16264 36242
rect 16212 36178 16264 36184
rect 16120 36168 16172 36174
rect 16120 36110 16172 36116
rect 16132 36038 16160 36110
rect 16120 36032 16172 36038
rect 16120 35974 16172 35980
rect 16028 34604 16080 34610
rect 16028 34546 16080 34552
rect 15844 33856 15896 33862
rect 15844 33798 15896 33804
rect 15856 33658 15884 33798
rect 15844 33652 15896 33658
rect 15844 33594 15896 33600
rect 15856 32910 15884 33594
rect 16224 33454 16252 36178
rect 16396 33856 16448 33862
rect 16396 33798 16448 33804
rect 16408 33590 16436 33798
rect 16396 33584 16448 33590
rect 16396 33526 16448 33532
rect 16212 33448 16264 33454
rect 16212 33390 16264 33396
rect 16396 33448 16448 33454
rect 16396 33390 16448 33396
rect 16488 33448 16540 33454
rect 16488 33390 16540 33396
rect 15844 32904 15896 32910
rect 15844 32846 15896 32852
rect 16224 32842 16252 33390
rect 16408 32910 16436 33390
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 16212 32836 16264 32842
rect 16212 32778 16264 32784
rect 16224 32434 16252 32778
rect 16408 32502 16436 32846
rect 16396 32496 16448 32502
rect 16396 32438 16448 32444
rect 16212 32428 16264 32434
rect 16212 32370 16264 32376
rect 16500 31822 16528 33390
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 15764 31726 15884 31754
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 15660 31408 15712 31414
rect 15660 31350 15712 31356
rect 15672 30938 15700 31350
rect 15660 30932 15712 30938
rect 15660 30874 15712 30880
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15764 27538 15792 28358
rect 15856 28014 15884 31726
rect 16396 31136 16448 31142
rect 16396 31078 16448 31084
rect 16408 30666 16436 31078
rect 16592 30818 16620 32302
rect 16684 30938 16712 47382
rect 17408 47116 17460 47122
rect 17408 47058 17460 47064
rect 17314 37904 17370 37913
rect 17314 37839 17316 37848
rect 17368 37839 17370 37848
rect 17316 37810 17368 37816
rect 16856 37664 16908 37670
rect 16856 37606 16908 37612
rect 16868 37330 16896 37606
rect 16856 37324 16908 37330
rect 16856 37266 16908 37272
rect 16764 37188 16816 37194
rect 16764 37130 16816 37136
rect 16776 36106 16804 37130
rect 16764 36100 16816 36106
rect 16764 36042 16816 36048
rect 16776 35766 16804 36042
rect 16764 35760 16816 35766
rect 16764 35702 16816 35708
rect 16776 35154 16804 35702
rect 16764 35148 16816 35154
rect 16764 35090 16816 35096
rect 17040 35012 17092 35018
rect 17040 34954 17092 34960
rect 17052 34746 17080 34954
rect 17040 34740 17092 34746
rect 17040 34682 17092 34688
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 17040 34196 17092 34202
rect 17040 34138 17092 34144
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16868 32774 16896 33458
rect 17052 33318 17080 34138
rect 17236 34134 17264 34546
rect 17224 34128 17276 34134
rect 17224 34070 17276 34076
rect 17040 33312 17092 33318
rect 17040 33254 17092 33260
rect 17132 33312 17184 33318
rect 17132 33254 17184 33260
rect 17144 32910 17172 33254
rect 17328 33046 17356 34546
rect 17224 33040 17276 33046
rect 17224 32982 17276 32988
rect 17316 33040 17368 33046
rect 17316 32982 17368 32988
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16868 32042 16896 32710
rect 16868 32014 16988 32042
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16868 31278 16896 31826
rect 16960 31822 16988 32014
rect 17236 31822 17264 32982
rect 17328 32910 17356 32982
rect 17316 32904 17368 32910
rect 17316 32846 17368 32852
rect 17316 32768 17368 32774
rect 17316 32710 17368 32716
rect 17328 32570 17356 32710
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 16948 31816 17000 31822
rect 17224 31816 17276 31822
rect 17000 31764 17080 31770
rect 16948 31758 17080 31764
rect 17224 31758 17276 31764
rect 16960 31742 17080 31758
rect 17052 31346 17080 31742
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 16856 31272 16908 31278
rect 16856 31214 16908 31220
rect 16672 30932 16724 30938
rect 16672 30874 16724 30880
rect 16592 30790 16804 30818
rect 16396 30660 16448 30666
rect 16396 30602 16448 30608
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16316 29646 16344 30534
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16316 29034 16344 29582
rect 16408 29578 16436 30602
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16592 29714 16620 30534
rect 16580 29708 16632 29714
rect 16580 29650 16632 29656
rect 16488 29640 16540 29646
rect 16488 29582 16540 29588
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16304 29028 16356 29034
rect 16304 28970 16356 28976
rect 15844 28008 15896 28014
rect 15844 27950 15896 27956
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15580 24886 15608 25094
rect 15568 24880 15620 24886
rect 15568 24822 15620 24828
rect 15856 23730 15884 25842
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15948 25226 15976 25638
rect 16316 25430 16344 26182
rect 16304 25424 16356 25430
rect 16304 25366 16356 25372
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15948 23254 15976 24142
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 16316 22030 16344 25366
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16316 20942 16344 21966
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16408 21622 16436 21830
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15488 18834 15516 19654
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15672 17678 15700 18226
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15672 17202 15700 17614
rect 15948 17202 15976 20878
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16316 19786 16344 20334
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16658 15884 16934
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15948 16114 15976 17138
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16408 3398 16436 3538
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16500 2582 16528 29582
rect 16776 24138 16804 30790
rect 16868 30394 16896 31214
rect 17040 31204 17092 31210
rect 17040 31146 17092 31152
rect 17052 30802 17080 31146
rect 17316 31136 17368 31142
rect 17316 31078 17368 31084
rect 17328 30938 17356 31078
rect 17132 30932 17184 30938
rect 17132 30874 17184 30880
rect 17316 30932 17368 30938
rect 17316 30874 17368 30880
rect 17040 30796 17092 30802
rect 17040 30738 17092 30744
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 16868 29510 16896 30330
rect 16948 30184 17000 30190
rect 16948 30126 17000 30132
rect 16960 29850 16988 30126
rect 17052 30054 17080 30738
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 16948 29844 17000 29850
rect 16948 29786 17000 29792
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 17052 28014 17080 29990
rect 17040 28008 17092 28014
rect 17040 27950 17092 27956
rect 17052 27062 17080 27950
rect 17040 27056 17092 27062
rect 17040 26998 17092 27004
rect 17144 26926 17172 30874
rect 17420 29646 17448 47058
rect 18604 47048 18656 47054
rect 18604 46990 18656 46996
rect 17500 38004 17552 38010
rect 17500 37946 17552 37952
rect 18512 38004 18564 38010
rect 18512 37946 18564 37952
rect 17512 37890 17540 37946
rect 17684 37936 17736 37942
rect 17512 37884 17684 37890
rect 17512 37878 17736 37884
rect 17512 37862 17724 37878
rect 18144 37868 18196 37874
rect 18144 37810 18196 37816
rect 18420 37868 18472 37874
rect 18420 37810 18472 37816
rect 18156 36922 18184 37810
rect 18432 37126 18460 37810
rect 18524 37670 18552 37946
rect 18512 37664 18564 37670
rect 18512 37606 18564 37612
rect 18420 37120 18472 37126
rect 18420 37062 18472 37068
rect 18144 36916 18196 36922
rect 18144 36858 18196 36864
rect 18432 36786 18460 37062
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18144 36712 18196 36718
rect 18144 36654 18196 36660
rect 18052 36644 18104 36650
rect 18052 36586 18104 36592
rect 18064 35562 18092 36586
rect 18156 35630 18184 36654
rect 18432 35630 18460 36722
rect 18512 35692 18564 35698
rect 18512 35634 18564 35640
rect 18144 35624 18196 35630
rect 18144 35566 18196 35572
rect 18420 35624 18472 35630
rect 18420 35566 18472 35572
rect 18052 35556 18104 35562
rect 18052 35498 18104 35504
rect 17500 35488 17552 35494
rect 17500 35430 17552 35436
rect 17684 35488 17736 35494
rect 17684 35430 17736 35436
rect 17512 35018 17540 35430
rect 17500 35012 17552 35018
rect 17500 34954 17552 34960
rect 17592 34468 17644 34474
rect 17592 34410 17644 34416
rect 17604 34202 17632 34410
rect 17592 34196 17644 34202
rect 17592 34138 17644 34144
rect 17696 33998 17724 35430
rect 17776 34604 17828 34610
rect 17776 34546 17828 34552
rect 17788 34202 17816 34546
rect 17776 34196 17828 34202
rect 17776 34138 17828 34144
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17788 32910 17816 34138
rect 17868 33516 17920 33522
rect 17868 33458 17920 33464
rect 17880 33114 17908 33458
rect 17868 33108 17920 33114
rect 17868 33050 17920 33056
rect 17500 32904 17552 32910
rect 17500 32846 17552 32852
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 17512 32502 17540 32846
rect 17776 32768 17828 32774
rect 17776 32710 17828 32716
rect 17788 32502 17816 32710
rect 17500 32496 17552 32502
rect 17500 32438 17552 32444
rect 17776 32496 17828 32502
rect 17776 32438 17828 32444
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17880 32026 17908 32166
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 17500 31952 17552 31958
rect 17500 31894 17552 31900
rect 17684 31952 17736 31958
rect 17684 31894 17736 31900
rect 17512 31754 17540 31894
rect 17696 31754 17724 31894
rect 17512 31726 17724 31754
rect 17512 30734 17540 31726
rect 17880 30802 17908 31962
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 17868 30796 17920 30802
rect 17868 30738 17920 30744
rect 17500 30728 17552 30734
rect 17500 30670 17552 30676
rect 17972 30326 18000 31758
rect 18064 31142 18092 35498
rect 18432 34678 18460 35566
rect 18524 34950 18552 35634
rect 18616 35222 18644 46990
rect 18708 46918 18736 49200
rect 19996 47818 20024 49200
rect 19996 47790 20208 47818
rect 20076 47592 20128 47598
rect 20076 47534 20128 47540
rect 20088 47122 20116 47534
rect 20076 47116 20128 47122
rect 20076 47058 20128 47064
rect 19432 46980 19484 46986
rect 19432 46922 19484 46928
rect 19984 46980 20036 46986
rect 19984 46922 20036 46928
rect 18696 46912 18748 46918
rect 18696 46854 18748 46860
rect 19444 41414 19472 46922
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19996 45554 20024 46922
rect 20180 46918 20208 47790
rect 20260 47592 20312 47598
rect 20260 47534 20312 47540
rect 20272 47190 20300 47534
rect 20260 47184 20312 47190
rect 20260 47126 20312 47132
rect 20352 47184 20404 47190
rect 20352 47126 20404 47132
rect 20168 46912 20220 46918
rect 20168 46854 20220 46860
rect 20076 46504 20128 46510
rect 20076 46446 20128 46452
rect 20088 46170 20116 46446
rect 20076 46164 20128 46170
rect 20076 46106 20128 46112
rect 19996 45526 20116 45554
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19352 41386 19472 41414
rect 19352 38962 19380 41386
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19984 39432 20036 39438
rect 19984 39374 20036 39380
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19996 38962 20024 39374
rect 19340 38956 19392 38962
rect 19340 38898 19392 38904
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 18972 38208 19024 38214
rect 19352 38185 19380 38898
rect 19984 38208 20036 38214
rect 18972 38150 19024 38156
rect 19338 38176 19394 38185
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18708 37913 18736 37946
rect 18694 37904 18750 37913
rect 18694 37839 18750 37848
rect 18984 37330 19012 38150
rect 19984 38150 20036 38156
rect 19338 38111 19394 38120
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19524 37964 19748 37992
rect 19248 37936 19300 37942
rect 19246 37904 19248 37913
rect 19300 37904 19302 37913
rect 19524 37890 19552 37964
rect 19444 37874 19552 37890
rect 19246 37839 19302 37848
rect 19432 37868 19552 37874
rect 19484 37862 19552 37868
rect 19432 37810 19484 37816
rect 19294 37800 19346 37806
rect 19346 37768 19394 37777
rect 19294 37742 19338 37748
rect 19306 37726 19338 37742
rect 19338 37703 19394 37712
rect 19616 37732 19668 37738
rect 19616 37674 19668 37680
rect 19248 37664 19300 37670
rect 19300 37624 19472 37652
rect 19248 37606 19300 37612
rect 19340 37460 19392 37466
rect 19340 37402 19392 37408
rect 18972 37324 19024 37330
rect 18972 37266 19024 37272
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 19260 36650 19288 37198
rect 19352 36718 19380 37402
rect 19444 36854 19472 37624
rect 19628 37466 19656 37674
rect 19616 37460 19668 37466
rect 19616 37402 19668 37408
rect 19720 37262 19748 37964
rect 19800 37936 19852 37942
rect 19800 37878 19852 37884
rect 19708 37256 19760 37262
rect 19708 37198 19760 37204
rect 19812 37194 19840 37878
rect 19996 37738 20024 38150
rect 19984 37732 20036 37738
rect 19984 37674 20036 37680
rect 19800 37188 19852 37194
rect 19800 37130 19852 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 19340 36712 19392 36718
rect 19340 36654 19392 36660
rect 19248 36644 19300 36650
rect 19248 36586 19300 36592
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19800 35624 19852 35630
rect 19800 35566 19852 35572
rect 19812 35290 19840 35566
rect 19800 35284 19852 35290
rect 19800 35226 19852 35232
rect 18604 35216 18656 35222
rect 18604 35158 18656 35164
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18420 34672 18472 34678
rect 18420 34614 18472 34620
rect 18524 34610 18552 34886
rect 19444 34678 19472 35022
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19432 34672 19484 34678
rect 19432 34614 19484 34620
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 19996 34406 20024 34954
rect 18788 34400 18840 34406
rect 18788 34342 18840 34348
rect 19432 34400 19484 34406
rect 19432 34342 19484 34348
rect 19984 34400 20036 34406
rect 19984 34342 20036 34348
rect 18512 33924 18564 33930
rect 18512 33866 18564 33872
rect 18524 32910 18552 33866
rect 18800 33454 18828 34342
rect 19338 33824 19394 33833
rect 19338 33759 19394 33768
rect 18788 33448 18840 33454
rect 18788 33390 18840 33396
rect 18512 32904 18564 32910
rect 18432 32864 18512 32892
rect 18432 31890 18460 32864
rect 18512 32846 18564 32852
rect 18512 32768 18564 32774
rect 18512 32710 18564 32716
rect 18524 32502 18552 32710
rect 18512 32496 18564 32502
rect 18512 32438 18564 32444
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 18064 30870 18092 31078
rect 18052 30864 18104 30870
rect 18052 30806 18104 30812
rect 18340 30734 18368 31282
rect 18432 30938 18460 31826
rect 18420 30932 18472 30938
rect 18420 30874 18472 30880
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18788 30728 18840 30734
rect 18788 30670 18840 30676
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 17328 29170 17356 29446
rect 18144 29232 18196 29238
rect 18142 29200 18144 29209
rect 18196 29200 18198 29209
rect 17316 29164 17368 29170
rect 17316 29106 17368 29112
rect 17408 29164 17460 29170
rect 18142 29135 18198 29144
rect 17408 29106 17460 29112
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 17236 28558 17264 29038
rect 17420 28994 17448 29106
rect 17420 28966 17540 28994
rect 17512 28762 17540 28966
rect 17960 28960 18012 28966
rect 17960 28902 18012 28908
rect 17500 28756 17552 28762
rect 17500 28698 17552 28704
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17236 28218 17264 28494
rect 17224 28212 17276 28218
rect 17224 28154 17276 28160
rect 17972 28014 18000 28902
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 16856 26920 16908 26926
rect 16856 26862 16908 26868
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 16868 26586 16896 26862
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 16960 24818 16988 26250
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17144 25498 17172 25842
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17420 25498 17448 25638
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 17144 24818 17172 25434
rect 17420 25294 17448 25434
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 23730 16712 24006
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16960 23322 16988 24142
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 17236 22094 17264 25230
rect 17604 23662 17632 27338
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 18064 25362 18092 25842
rect 18248 25770 18276 28426
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 18616 27606 18644 28086
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 18696 27464 18748 27470
rect 18696 27406 18748 27412
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 18524 25974 18552 26318
rect 18708 26314 18736 27406
rect 18800 26790 18828 30670
rect 19156 28620 19208 28626
rect 19156 28562 19208 28568
rect 19168 27946 19196 28562
rect 19352 28506 19380 33759
rect 19444 29288 19472 34342
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19708 32360 19760 32366
rect 19708 32302 19760 32308
rect 19720 31822 19748 32302
rect 19996 32026 20024 32846
rect 19984 32020 20036 32026
rect 19984 31962 20036 31968
rect 19708 31816 19760 31822
rect 19708 31758 19760 31764
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19984 29572 20036 29578
rect 19984 29514 20036 29520
rect 19996 29481 20024 29514
rect 19982 29472 20038 29481
rect 19574 29404 19882 29424
rect 19982 29407 20038 29416
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19444 29260 19564 29288
rect 19536 28694 19564 29260
rect 19996 29170 20024 29407
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19800 28756 19852 28762
rect 19800 28698 19852 28704
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 19524 28688 19576 28694
rect 19524 28630 19576 28636
rect 19260 28478 19380 28506
rect 19156 27940 19208 27946
rect 19156 27882 19208 27888
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18800 26518 18828 26726
rect 18788 26512 18840 26518
rect 18788 26454 18840 26460
rect 18984 26450 19012 26862
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 19260 26382 19288 28478
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19352 27062 19380 28358
rect 19444 27962 19472 28630
rect 19812 28626 19840 28698
rect 19800 28620 19852 28626
rect 19800 28562 19852 28568
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19996 28150 20024 28426
rect 19984 28144 20036 28150
rect 19984 28086 20036 28092
rect 19444 27934 19564 27962
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19444 27674 19472 27814
rect 19536 27674 19564 27934
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19984 27056 20036 27062
rect 19984 26998 20036 27004
rect 19996 26586 20024 26998
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 18696 26308 18748 26314
rect 18696 26250 18748 26256
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18236 25764 18288 25770
rect 18236 25706 18288 25712
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 17684 24608 17736 24614
rect 17684 24550 17736 24556
rect 17696 24138 17724 24550
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17328 23254 17356 23462
rect 17316 23248 17368 23254
rect 17316 23190 17368 23196
rect 17328 23118 17356 23190
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 18248 22642 18276 25706
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19444 24954 19472 25162
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 19260 24206 19288 24618
rect 19536 24614 19564 24754
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19536 24206 19564 24550
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18616 23594 18644 24006
rect 19260 23866 19288 24142
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 19352 23322 19380 24074
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23730 19472 24006
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19444 22982 19472 23666
rect 19996 23662 20024 24550
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19536 23118 19564 23258
rect 19996 23118 20024 23598
rect 19524 23112 19576 23118
rect 19524 23054 19576 23060
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 17144 22066 17264 22094
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16592 21418 16620 21898
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16868 21622 16896 21830
rect 16856 21616 16908 21622
rect 16856 21558 16908 21564
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16592 20806 16620 21014
rect 17144 20942 17172 22066
rect 18248 21962 18276 22578
rect 18236 21956 18288 21962
rect 18236 21898 18288 21904
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 17316 21072 17368 21078
rect 17316 21014 17368 21020
rect 17328 20942 17356 21014
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 17040 20868 17092 20874
rect 17040 20810 17092 20816
rect 17592 20868 17644 20874
rect 17592 20810 17644 20816
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16592 17678 16620 20742
rect 16776 20482 16804 20742
rect 16684 20454 16804 20482
rect 16856 20460 16908 20466
rect 16684 18290 16712 20454
rect 16856 20402 16908 20408
rect 16868 20262 16896 20402
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16868 19378 16896 20198
rect 16960 19922 16988 20742
rect 17052 20534 17080 20810
rect 17040 20528 17092 20534
rect 17040 20470 17092 20476
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17236 19922 17264 20198
rect 17604 19922 17632 20810
rect 18064 20466 18092 21626
rect 18248 20942 18276 21898
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 18328 21072 18380 21078
rect 18328 21014 18380 21020
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17880 20058 17908 20402
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 18064 19718 18092 20402
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18156 19446 18184 20742
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16960 18970 16988 19382
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16764 18692 16816 18698
rect 16764 18634 16816 18640
rect 16776 18358 16804 18634
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16684 17746 16712 18226
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17696 17882 17724 18158
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17328 16726 17356 17478
rect 17512 17202 17540 17614
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16684 15434 16712 15982
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17236 3738 17264 4082
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 3738 17356 4014
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3058 16712 3334
rect 16776 3194 16804 3470
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15488 800 15516 2382
rect 15580 2038 15608 2382
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15568 2032 15620 2038
rect 15568 1974 15620 1980
rect 16132 800 16160 2314
rect 17420 800 17448 16662
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17512 6866 17540 16458
rect 18340 12434 18368 21014
rect 18616 20874 18644 21830
rect 19352 21622 19380 21830
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19444 21026 19472 22918
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19996 21690 20024 22034
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19260 20998 19472 21026
rect 19260 20942 19288 20998
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 18604 20868 18656 20874
rect 18604 20810 18656 20816
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19800 20528 19852 20534
rect 19892 20528 19944 20534
rect 19800 20470 19852 20476
rect 19890 20496 19892 20505
rect 19944 20496 19946 20505
rect 19812 20262 19840 20470
rect 19890 20431 19946 20440
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19812 20058 19840 20198
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19996 19854 20024 21422
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19156 19780 19208 19786
rect 19156 19722 19208 19728
rect 19168 19514 19196 19722
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18616 17882 18644 18294
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18708 17116 18736 17682
rect 18788 17128 18840 17134
rect 18708 17088 18788 17116
rect 18524 16794 18552 17070
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18708 16590 18736 17088
rect 18788 17070 18840 17076
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18340 12406 18736 12434
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 17604 2650 17632 4082
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17696 3534 17724 3878
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17788 2446 17816 3334
rect 17880 3058 17908 3878
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17972 3194 18000 3470
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 18248 2446 18276 3946
rect 18340 2650 18368 4082
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18524 3058 18552 3334
rect 18616 3194 18644 3470
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18708 800 18736 12406
rect 19076 5166 19104 19314
rect 19168 17678 19196 19314
rect 19444 18154 19472 19790
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19444 17678 19472 18090
rect 19812 17882 19840 18158
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19168 16114 19196 17614
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19444 16250 19472 17206
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19536 16522 19564 17002
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16590 19748 16934
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19168 15502 19196 16050
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20088 12434 20116 45526
rect 20364 40118 20392 47126
rect 20640 46510 20668 49200
rect 21088 47048 21140 47054
rect 21088 46990 21140 46996
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 21100 46034 21128 46990
rect 21284 46034 21312 49200
rect 21824 47252 21876 47258
rect 21824 47194 21876 47200
rect 21088 46028 21140 46034
rect 21088 45970 21140 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 20628 45960 20680 45966
rect 20628 45902 20680 45908
rect 20352 40112 20404 40118
rect 20352 40054 20404 40060
rect 20536 40112 20588 40118
rect 20536 40054 20588 40060
rect 20548 39914 20576 40054
rect 20536 39908 20588 39914
rect 20536 39850 20588 39856
rect 20352 39840 20404 39846
rect 20352 39782 20404 39788
rect 20260 39296 20312 39302
rect 20260 39238 20312 39244
rect 20272 38962 20300 39238
rect 20260 38956 20312 38962
rect 20260 38898 20312 38904
rect 20168 37936 20220 37942
rect 20166 37904 20168 37913
rect 20220 37904 20222 37913
rect 20166 37839 20222 37848
rect 20168 37800 20220 37806
rect 20168 37742 20220 37748
rect 20180 37330 20208 37742
rect 20168 37324 20220 37330
rect 20168 37266 20220 37272
rect 20168 36168 20220 36174
rect 20272 36156 20300 38898
rect 20220 36128 20300 36156
rect 20168 36110 20220 36116
rect 20180 31686 20208 36110
rect 20260 35624 20312 35630
rect 20260 35566 20312 35572
rect 20272 34950 20300 35566
rect 20260 34944 20312 34950
rect 20260 34886 20312 34892
rect 20272 34610 20300 34886
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20260 32836 20312 32842
rect 20260 32778 20312 32784
rect 20272 32570 20300 32778
rect 20260 32564 20312 32570
rect 20260 32506 20312 32512
rect 20364 32434 20392 39782
rect 20444 38820 20496 38826
rect 20444 38762 20496 38768
rect 20456 37874 20484 38762
rect 20548 38457 20576 39850
rect 20534 38448 20590 38457
rect 20534 38383 20590 38392
rect 20536 38276 20588 38282
rect 20536 38218 20588 38224
rect 20548 38010 20576 38218
rect 20536 38004 20588 38010
rect 20536 37946 20588 37952
rect 20534 37904 20590 37913
rect 20444 37868 20496 37874
rect 20534 37839 20590 37848
rect 20444 37810 20496 37816
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20456 33658 20484 34886
rect 20548 33998 20576 37839
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20548 33658 20576 33934
rect 20444 33652 20496 33658
rect 20444 33594 20496 33600
rect 20536 33652 20588 33658
rect 20536 33594 20588 33600
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20168 31680 20220 31686
rect 20168 31622 20220 31628
rect 20180 31346 20208 31622
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20168 31136 20220 31142
rect 20168 31078 20220 31084
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20180 30666 20208 31078
rect 20168 30660 20220 30666
rect 20168 30602 20220 30608
rect 20456 30394 20484 31078
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 20548 30394 20576 30738
rect 20444 30388 20496 30394
rect 20444 30330 20496 30336
rect 20536 30388 20588 30394
rect 20536 30330 20588 30336
rect 20534 30288 20590 30297
rect 20534 30223 20536 30232
rect 20588 30223 20590 30232
rect 20536 30194 20588 30200
rect 20352 30116 20404 30122
rect 20352 30058 20404 30064
rect 20444 30116 20496 30122
rect 20444 30058 20496 30064
rect 20168 29844 20220 29850
rect 20168 29786 20220 29792
rect 20180 28626 20208 29786
rect 20364 29170 20392 30058
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 20180 27538 20208 28562
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 23798 20208 24754
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 20180 21146 20208 23598
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20180 20534 20208 21082
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20180 17542 20208 19994
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20088 12406 20208 12434
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19352 4298 19380 4762
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19260 4270 19380 4298
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18800 3466 18828 3946
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 19260 2258 19288 4270
rect 20180 4214 20208 12406
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19352 2774 19380 4082
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 3058 19472 3470
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19706 3088 19762 3097
rect 19432 3052 19484 3058
rect 19996 3074 20024 3334
rect 19706 3023 19762 3032
rect 19812 3046 20024 3074
rect 19432 2994 19484 3000
rect 19720 2990 19748 3023
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19352 2746 19748 2774
rect 19720 2650 19748 2746
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19812 2446 19840 3046
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 19904 2360 19932 2926
rect 19996 2428 20024 2926
rect 20088 2650 20116 4082
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20180 2990 20208 4014
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20272 2650 20300 29106
rect 20456 29102 20484 30058
rect 20444 29096 20496 29102
rect 20444 29038 20496 29044
rect 20548 29034 20576 30194
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20364 23662 20392 24074
rect 20456 23866 20484 24142
rect 20548 24070 20576 24890
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20548 23866 20576 24006
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 20456 20330 20484 23802
rect 20548 23118 20576 23802
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20640 21962 20668 45902
rect 21088 45892 21140 45898
rect 21088 45834 21140 45840
rect 21100 45626 21128 45834
rect 21088 45620 21140 45626
rect 21088 45562 21140 45568
rect 21836 41414 21864 47194
rect 22008 47048 22060 47054
rect 22008 46990 22060 46996
rect 24584 47048 24636 47054
rect 24584 46990 24636 46996
rect 22020 46646 22048 46990
rect 22008 46640 22060 46646
rect 22008 46582 22060 46588
rect 24596 46578 24624 46990
rect 24584 46572 24636 46578
rect 24584 46514 24636 46520
rect 25148 46510 25176 49200
rect 25504 47048 25556 47054
rect 25504 46990 25556 46996
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25516 46034 25544 46990
rect 25792 46034 25820 49200
rect 25504 46028 25556 46034
rect 25504 45970 25556 45976
rect 25780 46028 25832 46034
rect 25780 45970 25832 45976
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25424 45626 25452 45834
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 26712 45554 26740 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49200 31014 50000
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49314 38098 50000
rect 37986 49286 38424 49314
rect 37986 49200 38098 49286
rect 28264 47592 28316 47598
rect 28264 47534 28316 47540
rect 27804 46980 27856 46986
rect 27804 46922 27856 46928
rect 26436 45526 26740 45554
rect 25136 44396 25188 44402
rect 25136 44338 25188 44344
rect 25148 41414 25176 44338
rect 26436 41414 26464 45526
rect 27252 45280 27304 45286
rect 27252 45222 27304 45228
rect 27264 44946 27292 45222
rect 27252 44940 27304 44946
rect 27252 44882 27304 44888
rect 27068 44872 27120 44878
rect 27068 44814 27120 44820
rect 27080 44538 27108 44814
rect 27068 44532 27120 44538
rect 27068 44474 27120 44480
rect 21836 41386 21956 41414
rect 25148 41386 25268 41414
rect 26436 41386 26556 41414
rect 21364 39432 21416 39438
rect 21364 39374 21416 39380
rect 21376 38418 21404 39374
rect 20812 38412 20864 38418
rect 20812 38354 20864 38360
rect 21364 38412 21416 38418
rect 21364 38354 21416 38360
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20732 36650 20760 37198
rect 20720 36644 20772 36650
rect 20720 36586 20772 36592
rect 20824 35834 20852 38354
rect 21272 38208 21324 38214
rect 21272 38150 21324 38156
rect 21284 37670 21312 38150
rect 20904 37664 20956 37670
rect 20904 37606 20956 37612
rect 21272 37664 21324 37670
rect 21272 37606 21324 37612
rect 20916 37466 20944 37606
rect 20904 37460 20956 37466
rect 20904 37402 20956 37408
rect 21284 37330 21312 37606
rect 21272 37324 21324 37330
rect 21272 37266 21324 37272
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 20812 35828 20864 35834
rect 20812 35770 20864 35776
rect 20720 35080 20772 35086
rect 20718 35048 20720 35057
rect 20772 35048 20774 35057
rect 20718 34983 20774 34992
rect 20824 34746 20852 35770
rect 20916 35698 20944 35974
rect 20904 35692 20956 35698
rect 20904 35634 20956 35640
rect 21088 35488 21140 35494
rect 21088 35430 21140 35436
rect 21272 35488 21324 35494
rect 21272 35430 21324 35436
rect 21100 35290 21128 35430
rect 21088 35284 21140 35290
rect 21088 35226 21140 35232
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 20720 34672 20772 34678
rect 20720 34614 20772 34620
rect 20904 34672 20956 34678
rect 20904 34614 20956 34620
rect 20732 34406 20760 34614
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20824 34218 20852 34546
rect 20732 34190 20852 34218
rect 20732 33998 20760 34190
rect 20720 33992 20772 33998
rect 20720 33934 20772 33940
rect 20732 31414 20760 33934
rect 20916 33318 20944 34614
rect 21100 34542 21128 35226
rect 21180 35148 21232 35154
rect 21180 35090 21232 35096
rect 21192 34950 21220 35090
rect 21284 35086 21312 35430
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 21272 35080 21324 35086
rect 21272 35022 21324 35028
rect 21180 34944 21232 34950
rect 21180 34886 21232 34892
rect 21192 34610 21220 34886
rect 21180 34604 21232 34610
rect 21180 34546 21232 34552
rect 20996 34536 21048 34542
rect 20996 34478 21048 34484
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21008 34406 21036 34478
rect 21468 34474 21496 35090
rect 21732 34944 21784 34950
rect 21732 34886 21784 34892
rect 21456 34468 21508 34474
rect 21456 34410 21508 34416
rect 20996 34400 21048 34406
rect 20996 34342 21048 34348
rect 21548 34400 21600 34406
rect 21548 34342 21600 34348
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 20812 32496 20864 32502
rect 20812 32438 20864 32444
rect 20824 31822 20852 32438
rect 20916 31958 20944 33254
rect 20996 33108 21048 33114
rect 20996 33050 21048 33056
rect 21008 32502 21036 33050
rect 21088 32768 21140 32774
rect 21088 32710 21140 32716
rect 20996 32496 21048 32502
rect 20996 32438 21048 32444
rect 21100 32434 21128 32710
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 20996 32292 21048 32298
rect 20996 32234 21048 32240
rect 21008 31958 21036 32234
rect 20904 31952 20956 31958
rect 20904 31894 20956 31900
rect 20996 31952 21048 31958
rect 20996 31894 21048 31900
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20720 31408 20772 31414
rect 20720 31350 20772 31356
rect 20732 30410 20760 31350
rect 20824 30802 20852 31758
rect 20904 31748 20956 31754
rect 20904 31690 20956 31696
rect 20916 31142 20944 31690
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20916 30938 20944 31078
rect 20904 30932 20956 30938
rect 20904 30874 20956 30880
rect 20812 30796 20864 30802
rect 20812 30738 20864 30744
rect 21008 30598 21036 31282
rect 21272 30796 21324 30802
rect 21272 30738 21324 30744
rect 20812 30592 20864 30598
rect 20810 30560 20812 30569
rect 20996 30592 21048 30598
rect 20864 30560 20866 30569
rect 20996 30534 21048 30540
rect 20810 30495 20866 30504
rect 20732 30382 20852 30410
rect 20720 30320 20772 30326
rect 20720 30262 20772 30268
rect 20732 29714 20760 30262
rect 20824 30258 20852 30382
rect 21008 30326 21036 30534
rect 20996 30320 21048 30326
rect 20996 30262 21048 30268
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 21180 30252 21232 30258
rect 21180 30194 21232 30200
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 21100 28082 21128 29582
rect 21192 28218 21220 30194
rect 21284 29850 21312 30738
rect 21456 30592 21508 30598
rect 21456 30534 21508 30540
rect 21468 29850 21496 30534
rect 21560 29850 21588 34342
rect 21744 34066 21772 34886
rect 21732 34060 21784 34066
rect 21732 34002 21784 34008
rect 21744 31754 21772 34002
rect 21824 32768 21876 32774
rect 21824 32710 21876 32716
rect 21836 32502 21864 32710
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 21744 31726 21864 31754
rect 21640 30728 21692 30734
rect 21640 30670 21692 30676
rect 21272 29844 21324 29850
rect 21272 29786 21324 29792
rect 21456 29844 21508 29850
rect 21456 29786 21508 29792
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21560 29714 21588 29786
rect 21652 29714 21680 30670
rect 21548 29708 21600 29714
rect 21548 29650 21600 29656
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 21732 29572 21784 29578
rect 21732 29514 21784 29520
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21180 28212 21232 28218
rect 21180 28154 21232 28160
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 20732 27130 20760 28018
rect 21008 27674 21036 28018
rect 21088 27872 21140 27878
rect 21086 27840 21088 27849
rect 21140 27840 21142 27849
rect 21086 27775 21142 27784
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21008 27538 21036 27610
rect 21100 27606 21128 27775
rect 21088 27600 21140 27606
rect 21088 27542 21140 27548
rect 20996 27532 21048 27538
rect 20996 27474 21048 27480
rect 21088 27464 21140 27470
rect 21192 27452 21220 28154
rect 21468 28150 21496 29446
rect 21744 28694 21772 29514
rect 21836 29050 21864 31726
rect 21928 29170 21956 41386
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 22100 40384 22152 40390
rect 22100 40326 22152 40332
rect 22112 39506 22140 40326
rect 22940 40186 22968 40462
rect 22928 40180 22980 40186
rect 22928 40122 22980 40128
rect 23112 39976 23164 39982
rect 23112 39918 23164 39924
rect 22100 39500 22152 39506
rect 22100 39442 22152 39448
rect 22100 39364 22152 39370
rect 22100 39306 22152 39312
rect 22112 39098 22140 39306
rect 22928 39296 22980 39302
rect 22928 39238 22980 39244
rect 22100 39092 22152 39098
rect 22100 39034 22152 39040
rect 22940 38962 22968 39238
rect 23124 39098 23152 39918
rect 23112 39092 23164 39098
rect 23112 39034 23164 39040
rect 22928 38956 22980 38962
rect 22928 38898 22980 38904
rect 22560 38888 22612 38894
rect 22560 38830 22612 38836
rect 22192 38276 22244 38282
rect 22192 38218 22244 38224
rect 22204 36922 22232 38218
rect 22572 37126 22600 38830
rect 22836 38208 22888 38214
rect 22836 38150 22888 38156
rect 22848 37874 22876 38150
rect 22940 37890 22968 38898
rect 23480 38752 23532 38758
rect 23480 38694 23532 38700
rect 23492 38282 23520 38694
rect 23480 38276 23532 38282
rect 23480 38218 23532 38224
rect 24768 38276 24820 38282
rect 24768 38218 24820 38224
rect 23204 38208 23256 38214
rect 23204 38150 23256 38156
rect 22940 37874 23060 37890
rect 23216 37874 23244 38150
rect 24780 38010 24808 38218
rect 24768 38004 24820 38010
rect 24768 37946 24820 37952
rect 22836 37868 22888 37874
rect 22940 37868 23072 37874
rect 22940 37862 23020 37868
rect 22836 37810 22888 37816
rect 23020 37810 23072 37816
rect 23204 37868 23256 37874
rect 23204 37810 23256 37816
rect 24952 37868 25004 37874
rect 24952 37810 25004 37816
rect 22744 37800 22796 37806
rect 22744 37742 22796 37748
rect 22560 37120 22612 37126
rect 22560 37062 22612 37068
rect 22192 36916 22244 36922
rect 22192 36858 22244 36864
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 22572 36174 22600 36518
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 22192 36100 22244 36106
rect 22192 36042 22244 36048
rect 22204 35766 22232 36042
rect 22376 36032 22428 36038
rect 22376 35974 22428 35980
rect 22192 35760 22244 35766
rect 22192 35702 22244 35708
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22296 34610 22324 35634
rect 22388 35290 22416 35974
rect 22756 35698 22784 37742
rect 22848 37210 22876 37810
rect 23110 37768 23166 37777
rect 23110 37703 23166 37712
rect 22848 37182 23060 37210
rect 23032 36786 23060 37182
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 22848 36378 22876 36722
rect 22836 36372 22888 36378
rect 22836 36314 22888 36320
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 23032 35494 23060 36722
rect 23124 36106 23152 37703
rect 23204 37664 23256 37670
rect 23204 37606 23256 37612
rect 23296 37664 23348 37670
rect 23296 37606 23348 37612
rect 23572 37664 23624 37670
rect 23572 37606 23624 37612
rect 23216 37262 23244 37606
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 23204 36848 23256 36854
rect 23204 36790 23256 36796
rect 23112 36100 23164 36106
rect 23112 36042 23164 36048
rect 22468 35488 22520 35494
rect 22468 35430 22520 35436
rect 23020 35488 23072 35494
rect 23020 35430 23072 35436
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22388 35018 22416 35226
rect 22480 35154 22508 35430
rect 22468 35148 22520 35154
rect 22468 35090 22520 35096
rect 22376 35012 22428 35018
rect 22376 34954 22428 34960
rect 23124 34950 23152 36042
rect 23112 34944 23164 34950
rect 23112 34886 23164 34892
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22192 33924 22244 33930
rect 22192 33866 22244 33872
rect 22008 33584 22060 33590
rect 22060 33544 22140 33572
rect 22008 33526 22060 33532
rect 22112 33114 22140 33544
rect 22204 33522 22232 33866
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22480 33590 22508 33798
rect 22468 33584 22520 33590
rect 22468 33526 22520 33532
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 22204 31686 22232 32846
rect 23112 32496 23164 32502
rect 23112 32438 23164 32444
rect 23124 31754 23152 32438
rect 23112 31748 23164 31754
rect 23112 31690 23164 31696
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22572 30734 22600 31622
rect 23216 31362 23244 36790
rect 23308 36582 23336 37606
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23400 36582 23428 37198
rect 23296 36576 23348 36582
rect 23296 36518 23348 36524
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23296 36100 23348 36106
rect 23296 36042 23348 36048
rect 23308 35714 23336 36042
rect 23400 35834 23428 36518
rect 23584 36242 23612 37606
rect 24964 37466 24992 37810
rect 24952 37460 25004 37466
rect 24952 37402 25004 37408
rect 24124 37188 24176 37194
rect 24124 37130 24176 37136
rect 24136 36922 24164 37130
rect 24216 37120 24268 37126
rect 24216 37062 24268 37068
rect 24952 37120 25004 37126
rect 24952 37062 25004 37068
rect 24124 36916 24176 36922
rect 24124 36858 24176 36864
rect 23756 36848 23808 36854
rect 23756 36790 23808 36796
rect 23572 36236 23624 36242
rect 23572 36178 23624 36184
rect 23388 35828 23440 35834
rect 23388 35770 23440 35776
rect 23572 35760 23624 35766
rect 23570 35728 23572 35737
rect 23624 35728 23626 35737
rect 23308 35698 23520 35714
rect 23308 35692 23532 35698
rect 23308 35686 23480 35692
rect 23570 35663 23626 35672
rect 23480 35634 23532 35640
rect 23768 35086 23796 36790
rect 24124 36780 24176 36786
rect 24124 36722 24176 36728
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 23756 35080 23808 35086
rect 23756 35022 23808 35028
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23480 34400 23532 34406
rect 23480 34342 23532 34348
rect 23492 33998 23520 34342
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23676 33046 23704 34478
rect 23756 33856 23808 33862
rect 23756 33798 23808 33804
rect 23768 33590 23796 33798
rect 23756 33584 23808 33590
rect 23756 33526 23808 33532
rect 23664 33040 23716 33046
rect 23664 32982 23716 32988
rect 23480 32972 23532 32978
rect 23480 32914 23532 32920
rect 23492 32026 23520 32914
rect 23480 32020 23532 32026
rect 23480 31962 23532 31968
rect 23572 31952 23624 31958
rect 23572 31894 23624 31900
rect 23216 31334 23336 31362
rect 23584 31346 23612 31894
rect 23204 31272 23256 31278
rect 23204 31214 23256 31220
rect 22560 30728 22612 30734
rect 22560 30670 22612 30676
rect 23216 30666 23244 31214
rect 23204 30660 23256 30666
rect 23204 30602 23256 30608
rect 22100 30592 22152 30598
rect 22100 30534 22152 30540
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 21916 29164 21968 29170
rect 21916 29106 21968 29112
rect 21836 29022 21956 29050
rect 21732 28688 21784 28694
rect 21732 28630 21784 28636
rect 21456 28144 21508 28150
rect 21456 28086 21508 28092
rect 21468 27674 21496 28086
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 21824 27532 21876 27538
rect 21824 27474 21876 27480
rect 21272 27464 21324 27470
rect 21192 27424 21272 27452
rect 21088 27406 21140 27412
rect 21272 27406 21324 27412
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20732 24886 20760 25230
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 20732 24410 20760 24822
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20916 24274 20944 24754
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20916 23118 20944 24210
rect 21100 23866 21128 27406
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 21376 25294 21404 27270
rect 21836 27062 21864 27474
rect 21928 27470 21956 29022
rect 22112 28626 22140 30534
rect 22756 30326 22784 30534
rect 22744 30320 22796 30326
rect 22744 30262 22796 30268
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22848 29850 22876 30126
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22480 28994 22508 29582
rect 22296 28966 22508 28994
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22008 27940 22060 27946
rect 22008 27882 22060 27888
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 22020 27062 22048 27882
rect 22204 27130 22232 28086
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 21824 27056 21876 27062
rect 21824 26998 21876 27004
rect 22008 27056 22060 27062
rect 22008 26998 22060 27004
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22204 25906 22232 26250
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21192 24682 21220 25230
rect 21180 24676 21232 24682
rect 21180 24618 21232 24624
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21284 24274 21312 24550
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 21376 22710 21404 25230
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 21560 24274 21588 25094
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21836 23730 21864 24754
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21928 23798 21956 24006
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21824 23520 21876 23526
rect 21824 23462 21876 23468
rect 21836 23186 21864 23462
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 20548 19802 20576 21626
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 19854 20760 20742
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20456 19774 20576 19802
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20364 17270 20392 19722
rect 20456 17678 20484 19774
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20548 19378 20576 19654
rect 20640 19446 20668 19654
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20732 19394 20760 19790
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20732 19366 20852 19394
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20364 17066 20392 17206
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16590 20392 17002
rect 20548 16998 20576 19314
rect 20732 17270 20760 19366
rect 20824 19310 20852 19366
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20824 16522 20852 17478
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20916 16182 20944 21898
rect 22204 21554 22232 21966
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21652 20942 21680 21422
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21744 19854 21772 20198
rect 21836 19922 21864 20402
rect 21824 19916 21876 19922
rect 21824 19858 21876 19864
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21836 19446 21864 19654
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21836 18970 21864 19246
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21008 16658 21036 17206
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 21836 16250 21864 17070
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 22020 16114 22048 18702
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22112 16794 22140 17070
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22296 12434 22324 28966
rect 22664 28558 22692 29582
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 23112 27872 23164 27878
rect 23112 27814 23164 27820
rect 23124 27674 23152 27814
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22572 26042 22600 26250
rect 22560 26036 22612 26042
rect 22560 25978 22612 25984
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 22572 15706 22600 17206
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22480 12986 22508 13194
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22204 12406 22324 12434
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22112 4690 22140 5170
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20824 4146 20852 4422
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20364 2990 20392 4082
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 3534 20760 3878
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20640 3126 20668 3334
rect 20732 3194 20760 3334
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20824 2854 20852 3130
rect 20916 2854 20944 4218
rect 21100 3602 21128 4558
rect 21376 4282 21404 4558
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21284 4134 21496 4162
rect 21284 4078 21312 4134
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 21008 3482 21036 3538
rect 21376 3482 21404 4014
rect 21468 3534 21496 4134
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21836 3534 21864 3878
rect 21008 3454 21404 3482
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21928 3176 21956 3878
rect 22020 3602 22048 3946
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 21836 3148 21956 3176
rect 21836 3097 21864 3148
rect 21822 3088 21878 3097
rect 21822 3023 21878 3032
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20076 2440 20128 2446
rect 19996 2400 20076 2428
rect 20076 2382 20128 2388
rect 20628 2372 20680 2378
rect 19904 2332 20024 2360
rect 19260 2230 19380 2258
rect 19352 800 19380 2230
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2332
rect 20628 2314 20680 2320
rect 20640 800 20668 2314
rect 21928 800 21956 2994
rect 22112 2854 22140 4082
rect 22204 3194 22232 12406
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22190 2952 22246 2961
rect 22190 2887 22192 2896
rect 22244 2887 22246 2896
rect 22192 2858 22244 2864
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22296 2514 22324 4966
rect 22388 4758 22416 12786
rect 22664 12434 22692 26862
rect 23124 26586 23152 27406
rect 23216 27334 23244 30602
rect 23308 29510 23336 31334
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23756 31204 23808 31210
rect 23756 31146 23808 31152
rect 23664 30796 23716 30802
rect 23664 30738 23716 30744
rect 23388 30116 23440 30122
rect 23388 30058 23440 30064
rect 23400 29578 23428 30058
rect 23676 30054 23704 30738
rect 23768 30598 23796 31146
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23768 29714 23796 29990
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23204 27328 23256 27334
rect 23204 27270 23256 27276
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 23112 26444 23164 26450
rect 23112 26386 23164 26392
rect 23124 26042 23152 26386
rect 23112 26036 23164 26042
rect 23112 25978 23164 25984
rect 22928 25900 22980 25906
rect 22928 25842 22980 25848
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22848 23866 22876 24074
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22756 23254 22784 23666
rect 22744 23248 22796 23254
rect 22744 23190 22796 23196
rect 22756 22642 22784 23190
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22848 22778 22876 23054
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22756 21418 22784 21898
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22756 14890 22784 21354
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22848 13394 22876 20742
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22664 12406 22784 12434
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22388 4078 22416 4558
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22480 4146 22508 4422
rect 22664 4282 22692 4558
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22756 4214 22784 12406
rect 22940 5030 22968 25842
rect 23216 21554 23244 27270
rect 23308 26994 23336 29446
rect 23388 28076 23440 28082
rect 23664 28076 23716 28082
rect 23388 28018 23440 28024
rect 23584 28036 23664 28064
rect 23400 27878 23428 28018
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23388 27600 23440 27606
rect 23388 27542 23440 27548
rect 23400 27402 23428 27542
rect 23388 27396 23440 27402
rect 23388 27338 23440 27344
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 23308 26874 23336 26930
rect 23308 26846 23428 26874
rect 23400 25906 23428 26846
rect 23584 26586 23612 28036
rect 23664 28018 23716 28024
rect 23754 27840 23810 27849
rect 23754 27775 23810 27784
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23676 25906 23704 27610
rect 23768 27538 23796 27775
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 23768 25974 23796 27270
rect 23756 25968 23808 25974
rect 23756 25910 23808 25916
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23400 23322 23428 24686
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23388 22092 23440 22098
rect 23860 22094 23888 36110
rect 24136 35834 24164 36722
rect 24124 35828 24176 35834
rect 24124 35770 24176 35776
rect 24124 35012 24176 35018
rect 24124 34954 24176 34960
rect 23940 33312 23992 33318
rect 23940 33254 23992 33260
rect 23952 32910 23980 33254
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 24136 32230 24164 34954
rect 24228 32570 24256 37062
rect 24964 36786 24992 37062
rect 25044 36848 25096 36854
rect 25044 36790 25096 36796
rect 24952 36780 25004 36786
rect 24952 36722 25004 36728
rect 24860 36712 24912 36718
rect 24860 36654 24912 36660
rect 24768 36100 24820 36106
rect 24768 36042 24820 36048
rect 24780 35698 24808 36042
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 24676 35624 24728 35630
rect 24676 35566 24728 35572
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 24412 33998 24440 35022
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24308 33652 24360 33658
rect 24308 33594 24360 33600
rect 24216 32564 24268 32570
rect 24216 32506 24268 32512
rect 24124 32224 24176 32230
rect 24124 32166 24176 32172
rect 24136 31482 24164 32166
rect 24228 31958 24256 32506
rect 24216 31952 24268 31958
rect 24216 31894 24268 31900
rect 24124 31476 24176 31482
rect 24124 31418 24176 31424
rect 24320 29646 24348 33594
rect 24412 32570 24440 33934
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24400 32564 24452 32570
rect 24400 32506 24452 32512
rect 24400 31952 24452 31958
rect 24400 31894 24452 31900
rect 24412 30258 24440 31894
rect 24596 31498 24624 33798
rect 24504 31470 24624 31498
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24412 29782 24440 30194
rect 24400 29776 24452 29782
rect 24400 29718 24452 29724
rect 24308 29640 24360 29646
rect 24308 29582 24360 29588
rect 23940 29572 23992 29578
rect 23940 29514 23992 29520
rect 23952 29170 23980 29514
rect 23940 29164 23992 29170
rect 23940 29106 23992 29112
rect 24320 28422 24348 29582
rect 24504 29034 24532 31470
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24596 30870 24624 31282
rect 24688 31142 24716 35566
rect 24780 34542 24808 35634
rect 24872 35494 24900 36654
rect 25056 36378 25084 36790
rect 25240 36582 25268 41386
rect 25688 38276 25740 38282
rect 25688 38218 25740 38224
rect 25700 38010 25728 38218
rect 25964 38208 26016 38214
rect 25964 38150 26016 38156
rect 25688 38004 25740 38010
rect 25688 37946 25740 37952
rect 25976 37806 26004 38150
rect 25964 37800 26016 37806
rect 25964 37742 26016 37748
rect 25504 37392 25556 37398
rect 25504 37334 25556 37340
rect 25228 36576 25280 36582
rect 25228 36518 25280 36524
rect 25044 36372 25096 36378
rect 25044 36314 25096 36320
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24768 34536 24820 34542
rect 24768 34478 24820 34484
rect 25044 34468 25096 34474
rect 25044 34410 25096 34416
rect 25056 34202 25084 34410
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25044 34196 25096 34202
rect 25044 34138 25096 34144
rect 24768 32836 24820 32842
rect 24768 32778 24820 32784
rect 24676 31136 24728 31142
rect 24676 31078 24728 31084
rect 24584 30864 24636 30870
rect 24584 30806 24636 30812
rect 24596 30326 24624 30806
rect 24584 30320 24636 30326
rect 24584 30262 24636 30268
rect 24492 29028 24544 29034
rect 24492 28970 24544 28976
rect 24124 28416 24176 28422
rect 24124 28358 24176 28364
rect 24308 28416 24360 28422
rect 24308 28358 24360 28364
rect 24136 27946 24164 28358
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 24124 27940 24176 27946
rect 24124 27882 24176 27888
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24032 27532 24084 27538
rect 24032 27474 24084 27480
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 23952 27130 23980 27338
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23952 26586 23980 27066
rect 24044 26994 24072 27474
rect 24320 27062 24348 27814
rect 24412 27402 24440 27950
rect 24400 27396 24452 27402
rect 24400 27338 24452 27344
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24596 27130 24624 27338
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24308 27056 24360 27062
rect 24308 26998 24360 27004
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 23940 26580 23992 26586
rect 23940 26522 23992 26528
rect 24596 26518 24624 27066
rect 24584 26512 24636 26518
rect 24584 26454 24636 26460
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24504 25838 24532 26250
rect 24492 25832 24544 25838
rect 24492 25774 24544 25780
rect 24504 25294 24532 25774
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24688 25226 24716 28018
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23952 23798 23980 24006
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23860 22066 23980 22094
rect 23388 22034 23440 22040
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 23124 20874 23152 21082
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23216 20505 23244 21490
rect 23400 20806 23428 22034
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23572 20868 23624 20874
rect 23572 20810 23624 20816
rect 23388 20800 23440 20806
rect 23294 20768 23350 20777
rect 23388 20742 23440 20748
rect 23480 20800 23532 20806
rect 23584 20777 23612 20810
rect 23480 20742 23532 20748
rect 23570 20768 23626 20777
rect 23294 20703 23350 20712
rect 23202 20496 23258 20505
rect 23202 20431 23258 20440
rect 23020 18148 23072 18154
rect 23020 18090 23072 18096
rect 23032 15026 23060 18090
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23124 15366 23152 17818
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 23216 15978 23244 17546
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 23216 15706 23244 15914
rect 23308 15706 23336 20703
rect 23492 20602 23520 20742
rect 23570 20703 23626 20712
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23480 19984 23532 19990
rect 23480 19926 23532 19932
rect 23492 18766 23520 19926
rect 23584 19786 23612 20470
rect 23572 19780 23624 19786
rect 23572 19722 23624 19728
rect 23584 19514 23612 19722
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23860 18766 23888 21014
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23860 17610 23888 18702
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23492 16590 23520 17478
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23584 16590 23612 16934
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 23400 15162 23428 15982
rect 23584 15434 23612 16526
rect 23860 15502 23888 17546
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23860 14958 23888 15438
rect 23848 14952 23900 14958
rect 23848 14894 23900 14900
rect 23020 14884 23072 14890
rect 23020 14826 23072 14832
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22744 4208 22796 4214
rect 22744 4150 22796 4156
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 23032 3754 23060 14826
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23112 5092 23164 5098
rect 23112 5034 23164 5040
rect 23124 4146 23152 5034
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22848 3726 23060 3754
rect 23216 3738 23244 4082
rect 23204 3732 23256 3738
rect 22756 3641 22784 3674
rect 22742 3632 22798 3641
rect 22742 3567 22798 3576
rect 22848 3398 22876 3726
rect 23204 3674 23256 3680
rect 22928 3664 22980 3670
rect 22928 3606 22980 3612
rect 22836 3392 22888 3398
rect 22558 3360 22614 3369
rect 22836 3334 22888 3340
rect 22558 3295 22614 3304
rect 22572 3126 22600 3295
rect 22560 3120 22612 3126
rect 22560 3062 22612 3068
rect 22836 3052 22888 3058
rect 22940 3040 22968 3606
rect 22888 3012 22968 3040
rect 22836 2994 22888 3000
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22388 2446 22416 2858
rect 23492 2774 23520 4558
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23216 2746 23520 2774
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22560 1420 22612 1426
rect 22560 1362 22612 1368
rect 22572 800 22600 1362
rect 23216 800 23244 2746
rect 23584 1426 23612 2926
rect 23676 2650 23704 13330
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23768 4146 23796 4626
rect 23860 4146 23888 5170
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23860 2514 23888 3470
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 23952 2106 23980 22066
rect 24688 21554 24716 25162
rect 24780 24682 24808 32778
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 24964 32298 24992 32370
rect 25148 32298 25176 34342
rect 24952 32292 25004 32298
rect 24952 32234 25004 32240
rect 25136 32292 25188 32298
rect 25136 32234 25188 32240
rect 24964 32026 24992 32234
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24952 32020 25004 32026
rect 24952 31962 25004 31968
rect 24872 31872 24900 31962
rect 25148 31940 25176 32234
rect 25056 31912 25176 31940
rect 24872 31844 24992 31872
rect 24860 31748 24912 31754
rect 24860 31690 24912 31696
rect 24872 30938 24900 31690
rect 24964 31686 24992 31844
rect 24952 31680 25004 31686
rect 24952 31622 25004 31628
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24872 27946 24900 30670
rect 24952 29640 25004 29646
rect 24952 29582 25004 29588
rect 24964 29481 24992 29582
rect 24950 29472 25006 29481
rect 24950 29407 25006 29416
rect 25056 28558 25084 31912
rect 25136 31680 25188 31686
rect 25136 31622 25188 31628
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 24860 27940 24912 27946
rect 24860 27882 24912 27888
rect 25056 26382 25084 28494
rect 25148 28014 25176 31622
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 24768 24676 24820 24682
rect 24768 24618 24820 24624
rect 24964 23798 24992 25094
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24964 22030 24992 23054
rect 25240 23050 25268 36518
rect 25516 36378 25544 37334
rect 25596 37324 25648 37330
rect 25596 37266 25648 37272
rect 25504 36372 25556 36378
rect 25504 36314 25556 36320
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25516 35698 25544 36110
rect 25504 35692 25556 35698
rect 25504 35634 25556 35640
rect 25412 34060 25464 34066
rect 25412 34002 25464 34008
rect 25424 33658 25452 34002
rect 25412 33652 25464 33658
rect 25412 33594 25464 33600
rect 25320 33380 25372 33386
rect 25320 33322 25372 33328
rect 25332 30734 25360 33322
rect 25412 33312 25464 33318
rect 25412 33254 25464 33260
rect 25424 32502 25452 33254
rect 25412 32496 25464 32502
rect 25412 32438 25464 32444
rect 25424 31686 25452 32438
rect 25516 31890 25544 35634
rect 25608 33386 25636 37266
rect 25688 36576 25740 36582
rect 25688 36518 25740 36524
rect 25700 36174 25728 36518
rect 25976 36394 26004 37742
rect 25884 36366 26004 36394
rect 25884 36174 25912 36366
rect 25964 36236 26016 36242
rect 25964 36178 26016 36184
rect 25688 36168 25740 36174
rect 25688 36110 25740 36116
rect 25872 36168 25924 36174
rect 25872 36110 25924 36116
rect 25688 35148 25740 35154
rect 25688 35090 25740 35096
rect 25596 33380 25648 33386
rect 25596 33322 25648 33328
rect 25700 32366 25728 35090
rect 25780 35080 25832 35086
rect 25780 35022 25832 35028
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 25792 33930 25820 35022
rect 25884 34746 25912 35022
rect 25872 34740 25924 34746
rect 25872 34682 25924 34688
rect 25780 33924 25832 33930
rect 25780 33866 25832 33872
rect 25688 32360 25740 32366
rect 25688 32302 25740 32308
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 25504 31884 25556 31890
rect 25504 31826 25556 31832
rect 25412 31680 25464 31686
rect 25412 31622 25464 31628
rect 25792 31346 25820 32166
rect 25976 31754 26004 36178
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26252 35737 26280 35974
rect 26238 35728 26294 35737
rect 26238 35663 26240 35672
rect 26292 35663 26294 35672
rect 26424 35692 26476 35698
rect 26240 35634 26292 35640
rect 26424 35634 26476 35640
rect 26252 35603 26280 35634
rect 26056 35556 26108 35562
rect 26056 35498 26108 35504
rect 26068 34610 26096 35498
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26252 34610 26280 35430
rect 26436 35154 26464 35634
rect 26424 35148 26476 35154
rect 26424 35090 26476 35096
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 26424 34400 26476 34406
rect 26424 34342 26476 34348
rect 26332 33924 26384 33930
rect 26332 33866 26384 33872
rect 26344 33658 26372 33866
rect 26148 33652 26200 33658
rect 26148 33594 26200 33600
rect 26332 33652 26384 33658
rect 26332 33594 26384 33600
rect 26160 33522 26188 33594
rect 26148 33516 26200 33522
rect 26148 33458 26200 33464
rect 26436 33046 26464 34342
rect 26424 33040 26476 33046
rect 26424 32982 26476 32988
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 25884 31726 26004 31754
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 25412 31136 25464 31142
rect 25412 31078 25464 31084
rect 25688 31136 25740 31142
rect 25688 31078 25740 31084
rect 25424 30938 25452 31078
rect 25412 30932 25464 30938
rect 25412 30874 25464 30880
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 25700 30258 25728 31078
rect 25688 30252 25740 30258
rect 25688 30194 25740 30200
rect 25504 30116 25556 30122
rect 25504 30058 25556 30064
rect 25320 29708 25372 29714
rect 25320 29650 25372 29656
rect 25332 29306 25360 29650
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25320 28008 25372 28014
rect 25320 27950 25372 27956
rect 25332 27606 25360 27950
rect 25320 27600 25372 27606
rect 25320 27542 25372 27548
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25332 26586 25360 26998
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25320 25764 25372 25770
rect 25320 25706 25372 25712
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24964 21554 24992 21966
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25148 21554 25176 21898
rect 25240 21690 25268 22986
rect 25228 21684 25280 21690
rect 25228 21626 25280 21632
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24952 21548 25004 21554
rect 24952 21490 25004 21496
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 24400 21412 24452 21418
rect 24400 21354 24452 21360
rect 24412 21010 24440 21354
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24596 21010 24624 21286
rect 24400 21004 24452 21010
rect 24400 20946 24452 20952
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24688 20942 24716 21490
rect 24872 21418 24900 21490
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24780 20602 24808 20742
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24872 20534 24900 21354
rect 24964 20942 24992 21490
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24136 19786 24164 20198
rect 25148 19922 25176 21490
rect 25332 20806 25360 25706
rect 25424 25362 25452 25842
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25412 20936 25464 20942
rect 25412 20878 25464 20884
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25424 20602 25452 20878
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 24044 17814 24072 19314
rect 24308 19304 24360 19310
rect 24308 19246 24360 19252
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24320 18834 24348 19246
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18902 24440 19110
rect 24596 18970 24624 19246
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24400 18896 24452 18902
rect 24400 18838 24452 18844
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 24688 18698 24716 19654
rect 24780 18902 24808 19722
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24872 18970 24900 19382
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24768 18896 24820 18902
rect 24768 18838 24820 18844
rect 24676 18692 24728 18698
rect 24676 18634 24728 18640
rect 24032 17808 24084 17814
rect 24032 17750 24084 17756
rect 24688 17202 24716 18634
rect 24780 18222 24808 18838
rect 25332 18766 25360 20198
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25424 18902 25452 19858
rect 25412 18896 25464 18902
rect 25412 18838 25464 18844
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 24412 16658 24440 16934
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 25136 16040 25188 16046
rect 25136 15982 25188 15988
rect 24320 3942 24348 15982
rect 25148 15706 25176 15982
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25240 15570 25268 16934
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24596 15366 24624 15438
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24596 15026 24624 15302
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 25332 12434 25360 18158
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25424 16250 25452 16594
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25240 12406 25360 12434
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24308 3936 24360 3942
rect 24308 3878 24360 3884
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24492 3460 24544 3466
rect 24492 3402 24544 3408
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 24504 800 24532 3402
rect 24688 2514 24716 3878
rect 24872 3670 24900 4082
rect 25240 4078 25268 12406
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 25226 3632 25282 3641
rect 25226 3567 25228 3576
rect 25280 3567 25282 3576
rect 25228 3538 25280 3544
rect 25332 3466 25360 4422
rect 25412 4072 25464 4078
rect 25412 4014 25464 4020
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25424 2582 25452 4014
rect 25516 4010 25544 30058
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25792 29073 25820 29106
rect 25778 29064 25834 29073
rect 25778 28999 25834 29008
rect 25596 28960 25648 28966
rect 25596 28902 25648 28908
rect 25608 27674 25636 28902
rect 25596 27668 25648 27674
rect 25596 27610 25648 27616
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25688 24268 25740 24274
rect 25688 24210 25740 24216
rect 25596 23588 25648 23594
rect 25596 23530 25648 23536
rect 25608 22982 25636 23530
rect 25700 23254 25728 24210
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25608 22234 25636 22578
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25608 21554 25636 21626
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25700 21010 25728 22374
rect 25688 21004 25740 21010
rect 25688 20946 25740 20952
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25596 15428 25648 15434
rect 25596 15370 25648 15376
rect 25608 14958 25636 15370
rect 25596 14952 25648 14958
rect 25596 14894 25648 14900
rect 25700 4282 25728 20742
rect 25792 14414 25820 25298
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25884 12434 25912 31726
rect 26068 30394 26096 32370
rect 26240 32224 26292 32230
rect 26160 32184 26240 32212
rect 26160 31890 26188 32184
rect 26240 32166 26292 32172
rect 26148 31884 26200 31890
rect 26148 31826 26200 31832
rect 26528 31754 26556 41386
rect 27344 38548 27396 38554
rect 27344 38490 27396 38496
rect 26976 38276 27028 38282
rect 26976 38218 27028 38224
rect 26988 38010 27016 38218
rect 26976 38004 27028 38010
rect 26976 37946 27028 37952
rect 26976 37868 27028 37874
rect 26976 37810 27028 37816
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 26988 37398 27016 37810
rect 27068 37800 27120 37806
rect 27068 37742 27120 37748
rect 26976 37392 27028 37398
rect 26976 37334 27028 37340
rect 27080 36922 27108 37742
rect 27172 37466 27200 37810
rect 27356 37806 27384 38490
rect 27620 38412 27672 38418
rect 27620 38354 27672 38360
rect 27528 37868 27580 37874
rect 27528 37810 27580 37816
rect 27344 37800 27396 37806
rect 27344 37742 27396 37748
rect 27436 37664 27488 37670
rect 27434 37632 27436 37641
rect 27488 37632 27490 37641
rect 27434 37567 27490 37576
rect 27160 37460 27212 37466
rect 27160 37402 27212 37408
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27068 36916 27120 36922
rect 27068 36858 27120 36864
rect 26792 36780 26844 36786
rect 26792 36722 26844 36728
rect 26700 36100 26752 36106
rect 26700 36042 26752 36048
rect 26712 35494 26740 36042
rect 26804 35714 26832 36722
rect 26884 36304 26936 36310
rect 26884 36246 26936 36252
rect 26896 36106 26924 36246
rect 26976 36168 27028 36174
rect 26976 36110 27028 36116
rect 26884 36100 26936 36106
rect 26884 36042 26936 36048
rect 26896 35834 26924 36042
rect 26884 35828 26936 35834
rect 26884 35770 26936 35776
rect 26988 35714 27016 36110
rect 27356 35834 27384 37198
rect 27344 35828 27396 35834
rect 27344 35770 27396 35776
rect 26804 35686 26924 35714
rect 26988 35686 27108 35714
rect 26700 35488 26752 35494
rect 26700 35430 26752 35436
rect 26712 35086 26740 35430
rect 26700 35080 26752 35086
rect 26700 35022 26752 35028
rect 26712 32434 26740 35022
rect 26896 34950 26924 35686
rect 27080 35630 27108 35686
rect 27068 35624 27120 35630
rect 27068 35566 27120 35572
rect 26976 35148 27028 35154
rect 27080 35136 27108 35566
rect 27356 35154 27384 35770
rect 27028 35108 27108 35136
rect 27344 35148 27396 35154
rect 26976 35090 27028 35096
rect 27344 35090 27396 35096
rect 26884 34944 26936 34950
rect 26884 34886 26936 34892
rect 26700 32428 26752 32434
rect 26700 32370 26752 32376
rect 26792 32360 26844 32366
rect 26792 32302 26844 32308
rect 26804 32026 26832 32302
rect 26792 32020 26844 32026
rect 26792 31962 26844 31968
rect 26528 31726 26648 31754
rect 26332 30592 26384 30598
rect 26332 30534 26384 30540
rect 26344 30394 26372 30534
rect 26056 30388 26108 30394
rect 26056 30330 26108 30336
rect 26332 30388 26384 30394
rect 26332 30330 26384 30336
rect 25962 30288 26018 30297
rect 25962 30223 25964 30232
rect 26016 30223 26018 30232
rect 26056 30252 26108 30258
rect 25964 30194 26016 30200
rect 26056 30194 26108 30200
rect 25976 28762 26004 30194
rect 26068 29510 26096 30194
rect 26332 30116 26384 30122
rect 26332 30058 26384 30064
rect 26344 29714 26372 30058
rect 26332 29708 26384 29714
rect 26332 29650 26384 29656
rect 26056 29504 26108 29510
rect 26056 29446 26108 29452
rect 26068 29306 26096 29446
rect 26056 29300 26108 29306
rect 26056 29242 26108 29248
rect 25964 28756 26016 28762
rect 25964 28698 26016 28704
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 26252 28218 26280 28494
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26160 26382 26188 26726
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 25964 25492 26016 25498
rect 25964 25434 26016 25440
rect 25976 25362 26004 25434
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 26160 24818 26188 26318
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 26148 24812 26200 24818
rect 26148 24754 26200 24760
rect 26252 24614 26280 25298
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26056 24268 26108 24274
rect 26056 24210 26108 24216
rect 25964 22160 26016 22166
rect 25964 22102 26016 22108
rect 25976 21690 26004 22102
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 26068 21486 26096 24210
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 26344 23866 26372 24142
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 26252 20602 26280 23666
rect 26436 22030 26464 24550
rect 26528 24138 26556 24754
rect 26516 24132 26568 24138
rect 26516 24074 26568 24080
rect 26528 23730 26556 24074
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26620 23526 26648 31726
rect 26700 30592 26752 30598
rect 26896 30569 26924 34886
rect 26988 34678 27016 35090
rect 27540 35057 27568 37810
rect 27632 36786 27660 38354
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 27724 36922 27752 37062
rect 27712 36916 27764 36922
rect 27712 36858 27764 36864
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 27632 35136 27660 36722
rect 27724 36174 27752 36858
rect 27816 36530 27844 46922
rect 28276 45554 28304 47534
rect 28368 47054 28396 49200
rect 29000 47252 29052 47258
rect 29000 47194 29052 47200
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 28276 45526 28396 45554
rect 28368 41414 28396 45526
rect 29012 41414 29040 47194
rect 29656 47054 29684 49200
rect 30196 47252 30248 47258
rect 30196 47194 30248 47200
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 28368 41386 28488 41414
rect 29012 41386 29132 41414
rect 27896 38752 27948 38758
rect 27896 38694 27948 38700
rect 27908 38282 27936 38694
rect 27896 38276 27948 38282
rect 27896 38218 27948 38224
rect 28356 38208 28408 38214
rect 28356 38150 28408 38156
rect 28368 37262 28396 38150
rect 27896 37256 27948 37262
rect 27896 37198 27948 37204
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 27908 36718 27936 37198
rect 27896 36712 27948 36718
rect 27948 36660 28028 36666
rect 27896 36654 28028 36660
rect 27908 36638 28028 36654
rect 27816 36502 27936 36530
rect 27712 36168 27764 36174
rect 27712 36110 27764 36116
rect 27712 35148 27764 35154
rect 27632 35108 27712 35136
rect 27526 35048 27582 35057
rect 27526 34983 27582 34992
rect 26976 34672 27028 34678
rect 26976 34614 27028 34620
rect 26988 34202 27016 34614
rect 26976 34196 27028 34202
rect 26976 34138 27028 34144
rect 27344 34196 27396 34202
rect 27344 34138 27396 34144
rect 27356 33590 27384 34138
rect 27344 33584 27396 33590
rect 27344 33526 27396 33532
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 26700 30534 26752 30540
rect 26882 30560 26938 30569
rect 26712 30326 26740 30534
rect 26882 30495 26938 30504
rect 26700 30320 26752 30326
rect 26700 30262 26752 30268
rect 26896 29306 26924 30495
rect 26988 30258 27016 33458
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 27264 31754 27292 31826
rect 27540 31822 27568 34983
rect 27632 34066 27660 35108
rect 27712 35090 27764 35096
rect 27620 34060 27672 34066
rect 27620 34002 27672 34008
rect 27632 33658 27660 34002
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27620 33652 27672 33658
rect 27620 33594 27672 33600
rect 27632 32570 27660 33594
rect 27620 32564 27672 32570
rect 27620 32506 27672 32512
rect 27724 32230 27752 33934
rect 27804 33516 27856 33522
rect 27804 33458 27856 33464
rect 27816 32842 27844 33458
rect 27804 32836 27856 32842
rect 27804 32778 27856 32784
rect 27712 32224 27764 32230
rect 27712 32166 27764 32172
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 27528 31816 27580 31822
rect 27528 31758 27580 31764
rect 27172 31726 27292 31754
rect 27068 30660 27120 30666
rect 27068 30602 27120 30608
rect 27080 30326 27108 30602
rect 27068 30320 27120 30326
rect 27068 30262 27120 30268
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 26884 29300 26936 29306
rect 26884 29242 26936 29248
rect 26974 29064 27030 29073
rect 26974 28999 26976 29008
rect 27028 28999 27030 29008
rect 26976 28970 27028 28976
rect 26976 24608 27028 24614
rect 26976 24550 27028 24556
rect 26988 23730 27016 24550
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26700 22160 26752 22166
rect 26700 22102 26752 22108
rect 26424 22024 26476 22030
rect 26424 21966 26476 21972
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26252 20466 26280 20538
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26436 19378 26464 21966
rect 26712 20874 26740 22102
rect 27172 22094 27200 31726
rect 27356 29850 27384 31758
rect 27528 31680 27580 31686
rect 27528 31622 27580 31628
rect 27436 31340 27488 31346
rect 27436 31282 27488 31288
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 27448 29186 27476 31282
rect 27356 29158 27476 29186
rect 27252 27464 27304 27470
rect 27252 27406 27304 27412
rect 27264 27130 27292 27406
rect 27252 27124 27304 27130
rect 27252 27066 27304 27072
rect 27356 26382 27384 29158
rect 27436 29096 27488 29102
rect 27436 29038 27488 29044
rect 27448 28558 27476 29038
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 27448 27402 27476 28494
rect 27540 28082 27568 31622
rect 27712 31136 27764 31142
rect 27712 31078 27764 31084
rect 27724 30394 27752 31078
rect 27816 30734 27844 32778
rect 27804 30728 27856 30734
rect 27804 30670 27856 30676
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27436 27396 27488 27402
rect 27436 27338 27488 27344
rect 27344 26376 27396 26382
rect 27344 26318 27396 26324
rect 27252 23656 27304 23662
rect 27252 23598 27304 23604
rect 27264 23322 27292 23598
rect 27252 23316 27304 23322
rect 27252 23258 27304 23264
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27356 22642 27384 22918
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27172 22066 27292 22094
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 26700 20868 26752 20874
rect 26700 20810 26752 20816
rect 26988 20466 27016 21626
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 27172 21146 27200 21286
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 26988 19854 27016 20402
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26436 18630 26464 19314
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 27080 18698 27108 19110
rect 27068 18692 27120 18698
rect 27068 18634 27120 18640
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26436 17202 26464 18566
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 27068 17196 27120 17202
rect 27068 17138 27120 17144
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 26056 16992 26108 16998
rect 26056 16934 26108 16940
rect 26068 16522 26096 16934
rect 26436 16658 26464 17138
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26160 16114 26188 16594
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26712 15502 26740 16390
rect 27080 16114 27108 17138
rect 27172 16114 27200 17138
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 26700 15496 26752 15502
rect 26700 15438 26752 15444
rect 25884 12406 26004 12434
rect 25976 9674 26004 12406
rect 25976 9646 26096 9674
rect 25688 4276 25740 4282
rect 25688 4218 25740 4224
rect 25596 4208 25648 4214
rect 25596 4150 25648 4156
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 25608 3126 25636 4150
rect 25596 3120 25648 3126
rect 25596 3062 25648 3068
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 25792 2854 25820 2994
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 26068 2650 26096 9646
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 26146 2952 26202 2961
rect 26252 2922 26280 2994
rect 26146 2887 26202 2896
rect 26240 2916 26292 2922
rect 26160 2854 26188 2887
rect 26240 2858 26292 2864
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 26056 2644 26108 2650
rect 26056 2586 26108 2592
rect 25412 2576 25464 2582
rect 25412 2518 25464 2524
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 800 25176 2450
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26436 800 26464 2382
rect 27080 800 27108 2994
rect 27172 2514 27200 16050
rect 27264 7698 27292 22066
rect 27356 21554 27384 22578
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27356 16726 27384 17546
rect 27344 16720 27396 16726
rect 27344 16662 27396 16668
rect 27356 12434 27384 16662
rect 27356 12406 27476 12434
rect 27264 7670 27384 7698
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 27264 3194 27292 3470
rect 27356 3194 27384 7670
rect 27448 3942 27476 12406
rect 27540 8838 27568 28018
rect 27632 27674 27660 29038
rect 27804 28960 27856 28966
rect 27804 28902 27856 28908
rect 27816 28558 27844 28902
rect 27804 28552 27856 28558
rect 27804 28494 27856 28500
rect 27620 27668 27672 27674
rect 27620 27610 27672 27616
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27632 26518 27660 26930
rect 27908 26874 27936 36502
rect 28000 36378 28028 36638
rect 27988 36372 28040 36378
rect 27988 36314 28040 36320
rect 28264 36168 28316 36174
rect 28264 36110 28316 36116
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 28000 32774 28028 33798
rect 28276 32892 28304 36110
rect 28092 32864 28304 32892
rect 27988 32768 28040 32774
rect 27988 32710 28040 32716
rect 27988 31816 28040 31822
rect 28092 31804 28120 32864
rect 28264 32496 28316 32502
rect 28264 32438 28316 32444
rect 28040 31776 28120 31804
rect 27988 31758 28040 31764
rect 28000 31210 28028 31758
rect 27988 31204 28040 31210
rect 27988 31146 28040 31152
rect 28000 28966 28028 31146
rect 28276 30326 28304 32438
rect 28356 32292 28408 32298
rect 28356 32234 28408 32240
rect 28368 31958 28396 32234
rect 28356 31952 28408 31958
rect 28356 31894 28408 31900
rect 28460 31754 28488 41386
rect 28816 38956 28868 38962
rect 28816 38898 28868 38904
rect 28828 37398 28856 38898
rect 28816 37392 28868 37398
rect 28816 37334 28868 37340
rect 29000 36848 29052 36854
rect 29000 36790 29052 36796
rect 28816 36576 28868 36582
rect 28816 36518 28868 36524
rect 28828 36242 28856 36518
rect 28816 36236 28868 36242
rect 28816 36178 28868 36184
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28552 35698 28580 35974
rect 28540 35692 28592 35698
rect 28540 35634 28592 35640
rect 28828 35630 28856 36178
rect 29012 35834 29040 36790
rect 29000 35828 29052 35834
rect 29000 35770 29052 35776
rect 29000 35692 29052 35698
rect 29000 35634 29052 35640
rect 28816 35624 28868 35630
rect 28816 35566 28868 35572
rect 28908 35624 28960 35630
rect 28908 35566 28960 35572
rect 28816 34128 28868 34134
rect 28816 34070 28868 34076
rect 28828 33658 28856 34070
rect 28816 33652 28868 33658
rect 28816 33594 28868 33600
rect 28724 32360 28776 32366
rect 28724 32302 28776 32308
rect 28540 32224 28592 32230
rect 28540 32166 28592 32172
rect 28552 31890 28580 32166
rect 28736 31890 28764 32302
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 28724 31884 28776 31890
rect 28724 31826 28776 31832
rect 28368 31726 28488 31754
rect 28632 31748 28684 31754
rect 28264 30320 28316 30326
rect 28264 30262 28316 30268
rect 27988 28960 28040 28966
rect 27988 28902 28040 28908
rect 28172 28960 28224 28966
rect 28172 28902 28224 28908
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 28000 27538 28028 28562
rect 28184 28558 28212 28902
rect 28172 28552 28224 28558
rect 28172 28494 28224 28500
rect 28264 28484 28316 28490
rect 28264 28426 28316 28432
rect 27988 27532 28040 27538
rect 27988 27474 28040 27480
rect 28000 26994 28028 27474
rect 28172 27464 28224 27470
rect 28276 27452 28304 28426
rect 28224 27424 28304 27452
rect 28172 27406 28224 27412
rect 28184 27130 28212 27406
rect 28172 27124 28224 27130
rect 28172 27066 28224 27072
rect 28368 27010 28396 31726
rect 28632 31690 28684 31696
rect 28644 31482 28672 31690
rect 28632 31476 28684 31482
rect 28632 31418 28684 31424
rect 28632 31340 28684 31346
rect 28736 31328 28764 31826
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28828 31346 28856 31758
rect 28684 31300 28764 31328
rect 28816 31340 28868 31346
rect 28632 31282 28684 31288
rect 28816 31282 28868 31288
rect 28724 31204 28776 31210
rect 28724 31146 28776 31152
rect 28736 30734 28764 31146
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 28540 29708 28592 29714
rect 28540 29650 28592 29656
rect 28448 29572 28500 29578
rect 28448 29514 28500 29520
rect 28460 28234 28488 29514
rect 28552 29170 28580 29650
rect 28736 29578 28764 30670
rect 28724 29572 28776 29578
rect 28724 29514 28776 29520
rect 28816 29572 28868 29578
rect 28816 29514 28868 29520
rect 28828 29238 28856 29514
rect 28816 29232 28868 29238
rect 28816 29174 28868 29180
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 28552 28490 28580 29106
rect 28632 28688 28684 28694
rect 28632 28630 28684 28636
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28460 28206 28580 28234
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28460 27674 28488 28018
rect 28552 28014 28580 28206
rect 28644 28150 28672 28630
rect 28724 28552 28776 28558
rect 28828 28540 28856 29174
rect 28776 28512 28856 28540
rect 28724 28494 28776 28500
rect 28632 28144 28684 28150
rect 28632 28086 28684 28092
rect 28540 28008 28592 28014
rect 28592 27956 28672 27962
rect 28540 27950 28672 27956
rect 28552 27934 28672 27950
rect 28540 27872 28592 27878
rect 28540 27814 28592 27820
rect 28448 27668 28500 27674
rect 28448 27610 28500 27616
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 28092 26982 28396 27010
rect 27724 26846 27936 26874
rect 27620 26512 27672 26518
rect 27620 26454 27672 26460
rect 27632 24818 27660 26454
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27724 21350 27752 26846
rect 27896 24608 27948 24614
rect 27896 24550 27948 24556
rect 27908 24138 27936 24550
rect 27896 24132 27948 24138
rect 27896 24074 27948 24080
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 28000 22098 28028 23598
rect 27988 22092 28040 22098
rect 27988 22034 28040 22040
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27436 3392 27488 3398
rect 27434 3360 27436 3369
rect 27488 3360 27490 3369
rect 27434 3295 27490 3304
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 27632 2990 27660 20742
rect 28092 19514 28120 26982
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 28368 26586 28396 26862
rect 28356 26580 28408 26586
rect 28356 26522 28408 26528
rect 28552 26382 28580 27814
rect 28644 27402 28672 27934
rect 28816 27464 28868 27470
rect 28816 27406 28868 27412
rect 28632 27396 28684 27402
rect 28632 27338 28684 27344
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28632 25832 28684 25838
rect 28632 25774 28684 25780
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 28552 23798 28580 24550
rect 28540 23792 28592 23798
rect 28540 23734 28592 23740
rect 28644 23662 28672 25774
rect 28724 24744 28776 24750
rect 28724 24686 28776 24692
rect 28736 24274 28764 24686
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28632 23656 28684 23662
rect 28632 23598 28684 23604
rect 28448 23180 28500 23186
rect 28448 23122 28500 23128
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28276 22778 28304 23054
rect 28460 23050 28488 23122
rect 28448 23044 28500 23050
rect 28448 22986 28500 22992
rect 28264 22772 28316 22778
rect 28264 22714 28316 22720
rect 28276 21554 28304 22714
rect 28460 22710 28488 22986
rect 28448 22704 28500 22710
rect 28448 22646 28500 22652
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28552 20942 28580 21898
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 28644 21146 28672 21422
rect 28632 21140 28684 21146
rect 28632 21082 28684 21088
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28828 20330 28856 27406
rect 28816 20324 28868 20330
rect 28816 20266 28868 20272
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28092 18442 28120 19450
rect 28632 19440 28684 19446
rect 28632 19382 28684 19388
rect 28448 19236 28500 19242
rect 28448 19178 28500 19184
rect 28460 18766 28488 19178
rect 28540 18828 28592 18834
rect 28540 18770 28592 18776
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28000 18414 28120 18442
rect 28000 18358 28028 18414
rect 27988 18352 28040 18358
rect 27988 18294 28040 18300
rect 28080 18352 28132 18358
rect 28080 18294 28132 18300
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27724 17610 27752 18226
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27816 17678 27844 18022
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27816 16590 27844 17614
rect 28092 17610 28120 18294
rect 28172 18216 28224 18222
rect 28172 18158 28224 18164
rect 28080 17604 28132 17610
rect 28080 17546 28132 17552
rect 28184 17542 28212 18158
rect 28460 18154 28488 18702
rect 28448 18148 28500 18154
rect 28448 18090 28500 18096
rect 28448 17604 28500 17610
rect 28448 17546 28500 17552
rect 27896 17536 27948 17542
rect 27896 17478 27948 17484
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 28264 17536 28316 17542
rect 28264 17478 28316 17484
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27816 4078 27844 16526
rect 27908 16114 27936 17478
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 28000 16726 28028 17138
rect 27988 16720 28040 16726
rect 27988 16662 28040 16668
rect 28092 16250 28120 17138
rect 28184 16454 28212 17478
rect 28276 17338 28304 17478
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 28276 16658 28304 17274
rect 28460 17270 28488 17546
rect 28448 17264 28500 17270
rect 28448 17206 28500 17212
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 28080 16244 28132 16250
rect 28080 16186 28132 16192
rect 28184 16182 28212 16390
rect 28552 16250 28580 18770
rect 28644 18766 28672 19382
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28540 16244 28592 16250
rect 28540 16186 28592 16192
rect 28172 16176 28224 16182
rect 28172 16118 28224 16124
rect 27896 16108 27948 16114
rect 27896 16050 27948 16056
rect 27804 4072 27856 4078
rect 27804 4014 27856 4020
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 27724 3126 27752 3878
rect 27816 3466 27844 4014
rect 27804 3460 27856 3466
rect 27804 3402 27856 3408
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 28920 2582 28948 35566
rect 29012 30054 29040 35634
rect 29104 31754 29132 41386
rect 29460 37256 29512 37262
rect 29460 37198 29512 37204
rect 29184 37120 29236 37126
rect 29184 37062 29236 37068
rect 29196 36854 29224 37062
rect 29184 36848 29236 36854
rect 29184 36790 29236 36796
rect 29276 36712 29328 36718
rect 29276 36654 29328 36660
rect 29288 35834 29316 36654
rect 29276 35828 29328 35834
rect 29276 35770 29328 35776
rect 29368 35828 29420 35834
rect 29368 35770 29420 35776
rect 29184 35692 29236 35698
rect 29184 35634 29236 35640
rect 29196 34474 29224 35634
rect 29380 34746 29408 35770
rect 29368 34740 29420 34746
rect 29368 34682 29420 34688
rect 29184 34468 29236 34474
rect 29184 34410 29236 34416
rect 29196 33402 29224 34410
rect 29368 33856 29420 33862
rect 29368 33798 29420 33804
rect 29380 33522 29408 33798
rect 29368 33516 29420 33522
rect 29368 33458 29420 33464
rect 29472 33402 29500 37198
rect 29644 35760 29696 35766
rect 29644 35702 29696 35708
rect 29196 33374 29316 33402
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 29196 32298 29224 33254
rect 29288 33114 29316 33374
rect 29380 33374 29500 33402
rect 29552 33380 29604 33386
rect 29276 33108 29328 33114
rect 29276 33050 29328 33056
rect 29184 32292 29236 32298
rect 29184 32234 29236 32240
rect 29196 32026 29224 32234
rect 29184 32020 29236 32026
rect 29184 31962 29236 31968
rect 29380 31754 29408 33374
rect 29552 33322 29604 33328
rect 29564 32570 29592 33322
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29104 31726 29224 31754
rect 29000 30048 29052 30054
rect 29000 29990 29052 29996
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29012 28422 29040 28698
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29000 23180 29052 23186
rect 29000 23122 29052 23128
rect 29012 22710 29040 23122
rect 29000 22704 29052 22710
rect 29000 22646 29052 22652
rect 29000 21480 29052 21486
rect 29000 21422 29052 21428
rect 29012 20534 29040 21422
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 29196 19990 29224 31726
rect 29288 31726 29408 31754
rect 29288 25294 29316 31726
rect 29656 30870 29684 35702
rect 30208 35698 30236 47194
rect 30944 47054 30972 49200
rect 30932 47048 30984 47054
rect 30932 46990 30984 46996
rect 32232 46442 32260 49200
rect 35440 47524 35492 47530
rect 35440 47466 35492 47472
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 32312 46504 32364 46510
rect 32312 46446 32364 46452
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32324 46170 32352 46446
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 32312 46164 32364 46170
rect 32312 46106 32364 46112
rect 31760 45960 31812 45966
rect 31760 45902 31812 45908
rect 31024 45484 31076 45490
rect 31024 45426 31076 45432
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 29932 34950 29960 35634
rect 30932 35488 30984 35494
rect 30932 35430 30984 35436
rect 30012 35284 30064 35290
rect 30012 35226 30064 35232
rect 29920 34944 29972 34950
rect 29920 34886 29972 34892
rect 29932 34610 29960 34886
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 29840 33590 29868 34478
rect 30024 33590 30052 35226
rect 30748 35012 30800 35018
rect 30748 34954 30800 34960
rect 30760 34746 30788 34954
rect 30748 34740 30800 34746
rect 30748 34682 30800 34688
rect 30840 34672 30892 34678
rect 30840 34614 30892 34620
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 30116 33930 30144 34546
rect 30852 33930 30880 34614
rect 30944 34610 30972 35430
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30104 33924 30156 33930
rect 30104 33866 30156 33872
rect 30840 33924 30892 33930
rect 30840 33866 30892 33872
rect 29828 33584 29880 33590
rect 29828 33526 29880 33532
rect 30012 33584 30064 33590
rect 30012 33526 30064 33532
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29748 32910 29776 33458
rect 29840 32978 29868 33526
rect 29828 32972 29880 32978
rect 29828 32914 29880 32920
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29644 30864 29696 30870
rect 29644 30806 29696 30812
rect 29552 30796 29604 30802
rect 29552 30738 29604 30744
rect 29368 30184 29420 30190
rect 29368 30126 29420 30132
rect 29380 29782 29408 30126
rect 29368 29776 29420 29782
rect 29368 29718 29420 29724
rect 29380 29102 29408 29718
rect 29460 29164 29512 29170
rect 29460 29106 29512 29112
rect 29368 29096 29420 29102
rect 29368 29038 29420 29044
rect 29472 28694 29500 29106
rect 29460 28688 29512 28694
rect 29460 28630 29512 28636
rect 29564 28626 29592 30738
rect 29644 30592 29696 30598
rect 29644 30534 29696 30540
rect 29656 30258 29684 30534
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29748 29850 29776 32846
rect 29840 32434 29868 32914
rect 29920 32496 29972 32502
rect 29920 32438 29972 32444
rect 29828 32428 29880 32434
rect 29828 32370 29880 32376
rect 29840 31822 29868 32370
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 29932 31278 29960 32438
rect 30116 32230 30144 33866
rect 30852 33454 30880 33866
rect 30840 33448 30892 33454
rect 30840 33390 30892 33396
rect 30104 32224 30156 32230
rect 30104 32166 30156 32172
rect 30380 32224 30432 32230
rect 30380 32166 30432 32172
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30024 31346 30052 31758
rect 30116 31482 30144 32166
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 30104 31476 30156 31482
rect 30104 31418 30156 31424
rect 30012 31340 30064 31346
rect 30012 31282 30064 31288
rect 29920 31272 29972 31278
rect 29920 31214 29972 31220
rect 29932 30938 29960 31214
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 29920 30932 29972 30938
rect 29920 30874 29972 30880
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29840 30190 29868 30670
rect 29932 30258 29960 30874
rect 30012 30864 30064 30870
rect 30012 30806 30064 30812
rect 30024 30734 30052 30806
rect 30116 30734 30144 31078
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29828 30184 29880 30190
rect 29828 30126 29880 30132
rect 29736 29844 29788 29850
rect 29736 29786 29788 29792
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29920 29640 29972 29646
rect 29920 29582 29972 29588
rect 29840 29102 29868 29582
rect 29932 29306 29960 29582
rect 30024 29306 30052 30670
rect 30300 29306 30328 31962
rect 30392 31754 30420 32166
rect 30380 31748 30432 31754
rect 30380 31690 30432 31696
rect 30392 31482 30420 31690
rect 30380 31476 30432 31482
rect 30380 31418 30432 31424
rect 30380 29776 30432 29782
rect 30380 29718 30432 29724
rect 29920 29300 29972 29306
rect 29920 29242 29972 29248
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 30288 29300 30340 29306
rect 30288 29242 30340 29248
rect 30012 29164 30064 29170
rect 30012 29106 30064 29112
rect 29828 29096 29880 29102
rect 29828 29038 29880 29044
rect 29552 28620 29604 28626
rect 29552 28562 29604 28568
rect 29552 27464 29604 27470
rect 29552 27406 29604 27412
rect 29564 26518 29592 27406
rect 29644 27056 29696 27062
rect 29644 26998 29696 27004
rect 29656 26586 29684 26998
rect 29644 26580 29696 26586
rect 29644 26522 29696 26528
rect 29552 26512 29604 26518
rect 29552 26454 29604 26460
rect 29564 26382 29592 26454
rect 29552 26376 29604 26382
rect 29552 26318 29604 26324
rect 29920 25832 29972 25838
rect 29920 25774 29972 25780
rect 29276 25288 29328 25294
rect 29276 25230 29328 25236
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29564 23254 29592 24142
rect 29656 23730 29684 25230
rect 29932 24954 29960 25774
rect 29920 24948 29972 24954
rect 29920 24890 29972 24896
rect 29736 24064 29788 24070
rect 29736 24006 29788 24012
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29644 23724 29696 23730
rect 29644 23666 29696 23672
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29552 23248 29604 23254
rect 29552 23190 29604 23196
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29564 22234 29592 22510
rect 29552 22228 29604 22234
rect 29552 22170 29604 22176
rect 29656 22030 29684 23462
rect 29748 22710 29776 24006
rect 29840 23866 29868 24006
rect 29828 23860 29880 23866
rect 29828 23802 29880 23808
rect 29736 22704 29788 22710
rect 29736 22646 29788 22652
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29656 21554 29684 21966
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29184 19984 29236 19990
rect 29184 19926 29236 19932
rect 29564 19718 29592 20878
rect 29736 20868 29788 20874
rect 29736 20810 29788 20816
rect 29748 20602 29776 20810
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29656 19514 29684 19790
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29288 18698 29316 19246
rect 29276 18692 29328 18698
rect 29276 18634 29328 18640
rect 29184 18080 29236 18086
rect 29184 18022 29236 18028
rect 29196 17202 29224 18022
rect 29748 17338 29776 20402
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 29932 18766 29960 19654
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 29920 18216 29972 18222
rect 29920 18158 29972 18164
rect 29932 17882 29960 18158
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29748 3602 29776 17274
rect 30024 12714 30052 29106
rect 30288 29028 30340 29034
rect 30288 28970 30340 28976
rect 30300 28762 30328 28970
rect 30392 28966 30420 29718
rect 30852 29646 30880 33390
rect 30840 29640 30892 29646
rect 30840 29582 30892 29588
rect 30932 29640 30984 29646
rect 30932 29582 30984 29588
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30380 28960 30432 28966
rect 30380 28902 30432 28908
rect 30288 28756 30340 28762
rect 30288 28698 30340 28704
rect 30300 28014 30328 28698
rect 30484 28626 30512 29446
rect 30472 28620 30524 28626
rect 30472 28562 30524 28568
rect 30380 28484 30432 28490
rect 30380 28426 30432 28432
rect 30288 28008 30340 28014
rect 30288 27950 30340 27956
rect 30392 27606 30420 28426
rect 30944 28218 30972 29582
rect 30932 28212 30984 28218
rect 30932 28154 30984 28160
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 31036 26450 31064 45426
rect 31772 37330 31800 45902
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 31760 37324 31812 37330
rect 31760 37266 31812 37272
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 32128 35148 32180 35154
rect 32128 35090 32180 35096
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31116 33856 31168 33862
rect 31116 33798 31168 33804
rect 31128 33522 31156 33798
rect 31116 33516 31168 33522
rect 31116 33458 31168 33464
rect 31772 33318 31800 33934
rect 32140 33522 32168 35090
rect 32220 35012 32272 35018
rect 32220 34954 32272 34960
rect 32232 34746 32260 34954
rect 32220 34740 32272 34746
rect 32220 34682 32272 34688
rect 32864 34604 32916 34610
rect 32864 34546 32916 34552
rect 32128 33516 32180 33522
rect 32128 33458 32180 33464
rect 31484 33312 31536 33318
rect 31484 33254 31536 33260
rect 31760 33312 31812 33318
rect 31760 33254 31812 33260
rect 31496 32910 31524 33254
rect 31772 32978 31800 33254
rect 31944 33040 31996 33046
rect 31944 32982 31996 32988
rect 31760 32972 31812 32978
rect 31760 32914 31812 32920
rect 31484 32904 31536 32910
rect 31484 32846 31536 32852
rect 31852 32904 31904 32910
rect 31852 32846 31904 32852
rect 31576 32836 31628 32842
rect 31576 32778 31628 32784
rect 31588 31822 31616 32778
rect 31760 32224 31812 32230
rect 31760 32166 31812 32172
rect 31772 31890 31800 32166
rect 31760 31884 31812 31890
rect 31760 31826 31812 31832
rect 31576 31816 31628 31822
rect 31576 31758 31628 31764
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 31128 30326 31156 30602
rect 31116 30320 31168 30326
rect 31116 30262 31168 30268
rect 31772 29170 31800 31826
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31300 29096 31352 29102
rect 31300 29038 31352 29044
rect 31312 28762 31340 29038
rect 31300 28756 31352 28762
rect 31300 28698 31352 28704
rect 31312 28082 31340 28698
rect 31300 28076 31352 28082
rect 31300 28018 31352 28024
rect 31208 27464 31260 27470
rect 31208 27406 31260 27412
rect 31220 26994 31248 27406
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31024 26444 31076 26450
rect 31024 26386 31076 26392
rect 30380 26376 30432 26382
rect 30380 26318 30432 26324
rect 30104 25424 30156 25430
rect 30104 25366 30156 25372
rect 30116 23118 30144 25366
rect 30392 25294 30420 26318
rect 31220 25974 31248 26930
rect 31484 26444 31536 26450
rect 31484 26386 31536 26392
rect 31208 25968 31260 25974
rect 31208 25910 31260 25916
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30392 25158 30420 25230
rect 30840 25220 30892 25226
rect 30840 25162 30892 25168
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 30392 24818 30420 25094
rect 30380 24812 30432 24818
rect 30432 24772 30512 24800
rect 30380 24754 30432 24760
rect 30484 24206 30512 24772
rect 30564 24336 30616 24342
rect 30564 24278 30616 24284
rect 30472 24200 30524 24206
rect 30472 24142 30524 24148
rect 30380 24132 30432 24138
rect 30380 24074 30432 24080
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30208 22030 30236 22374
rect 30196 22024 30248 22030
rect 30196 21966 30248 21972
rect 30392 20466 30420 24074
rect 30576 22098 30604 24278
rect 30656 23724 30708 23730
rect 30656 23666 30708 23672
rect 30668 22642 30696 23666
rect 30748 23520 30800 23526
rect 30748 23462 30800 23468
rect 30760 23186 30788 23462
rect 30748 23180 30800 23186
rect 30748 23122 30800 23128
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30564 22092 30616 22098
rect 30564 22034 30616 22040
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30484 21894 30512 21966
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30484 19922 30512 21830
rect 30852 20466 30880 25162
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 30944 22778 30972 23666
rect 30932 22772 30984 22778
rect 30932 22714 30984 22720
rect 30840 20460 30892 20466
rect 30840 20402 30892 20408
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30668 19922 30696 20198
rect 30472 19916 30524 19922
rect 30472 19858 30524 19864
rect 30656 19916 30708 19922
rect 30656 19858 30708 19864
rect 31128 19718 31156 24686
rect 31220 21690 31248 25910
rect 31392 25356 31444 25362
rect 31392 25298 31444 25304
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31312 24206 31340 24754
rect 31300 24200 31352 24206
rect 31300 24142 31352 24148
rect 31300 22432 31352 22438
rect 31300 22374 31352 22380
rect 31312 22098 31340 22374
rect 31300 22092 31352 22098
rect 31300 22034 31352 22040
rect 31208 21684 31260 21690
rect 31208 21626 31260 21632
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30392 18154 30420 18770
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 31024 18148 31076 18154
rect 31024 18090 31076 18096
rect 31036 17678 31064 18090
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 30564 16448 30616 16454
rect 30564 16390 30616 16396
rect 30576 15570 30604 16390
rect 30564 15564 30616 15570
rect 30564 15506 30616 15512
rect 30012 12708 30064 12714
rect 30012 12650 30064 12656
rect 30932 3664 30984 3670
rect 30932 3606 30984 3612
rect 29736 3596 29788 3602
rect 29736 3538 29788 3544
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28368 800 28396 2382
rect 29656 800 29684 2382
rect 30944 800 30972 3606
rect 31128 3398 31156 19654
rect 31404 19174 31432 25298
rect 31392 19168 31444 19174
rect 31392 19110 31444 19116
rect 31496 3534 31524 26386
rect 31668 24744 31720 24750
rect 31668 24686 31720 24692
rect 31680 24342 31708 24686
rect 31668 24336 31720 24342
rect 31668 24278 31720 24284
rect 31576 24064 31628 24070
rect 31576 24006 31628 24012
rect 31588 23730 31616 24006
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31588 23050 31616 23666
rect 31576 23044 31628 23050
rect 31576 22986 31628 22992
rect 31668 22092 31720 22098
rect 31668 22034 31720 22040
rect 31680 21962 31708 22034
rect 31668 21956 31720 21962
rect 31668 21898 31720 21904
rect 31760 4752 31812 4758
rect 31760 4694 31812 4700
rect 31484 3528 31536 3534
rect 31484 3470 31536 3476
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 31772 2650 31800 4694
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 31864 2310 31892 32846
rect 31956 32570 31984 32982
rect 32036 32904 32088 32910
rect 32036 32846 32088 32852
rect 31944 32564 31996 32570
rect 31944 32506 31996 32512
rect 32048 31822 32076 32846
rect 32140 32434 32168 33458
rect 32404 33448 32456 33454
rect 32404 33390 32456 33396
rect 32416 33114 32444 33390
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32876 32910 32904 34546
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 33140 33584 33192 33590
rect 33140 33526 33192 33532
rect 33152 33114 33180 33526
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 33140 33108 33192 33114
rect 33140 33050 33192 33056
rect 32864 32904 32916 32910
rect 32784 32864 32864 32892
rect 32128 32428 32180 32434
rect 32128 32370 32180 32376
rect 32404 32360 32456 32366
rect 32404 32302 32456 32308
rect 32416 32026 32444 32302
rect 32404 32020 32456 32026
rect 32404 31962 32456 31968
rect 32784 31822 32812 32864
rect 32864 32846 32916 32852
rect 32864 32496 32916 32502
rect 32864 32438 32916 32444
rect 32876 32026 32904 32438
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 32864 32020 32916 32026
rect 32864 31962 32916 31968
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 32128 31816 32180 31822
rect 32128 31758 32180 31764
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 32140 31346 32168 31758
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 32140 30394 32168 31282
rect 32220 31136 32272 31142
rect 32220 31078 32272 31084
rect 32232 30734 32260 31078
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 32220 30728 32272 30734
rect 32220 30670 32272 30676
rect 32128 30388 32180 30394
rect 32128 30330 32180 30336
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 33140 30184 33192 30190
rect 33140 30126 33192 30132
rect 33152 29850 33180 30126
rect 33140 29844 33192 29850
rect 33140 29786 33192 29792
rect 32956 29640 33008 29646
rect 32956 29582 33008 29588
rect 32772 29572 32824 29578
rect 32772 29514 32824 29520
rect 32784 29102 32812 29514
rect 32312 29096 32364 29102
rect 32312 29038 32364 29044
rect 32496 29096 32548 29102
rect 32496 29038 32548 29044
rect 32772 29096 32824 29102
rect 32772 29038 32824 29044
rect 32220 28552 32272 28558
rect 32220 28494 32272 28500
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 31944 24608 31996 24614
rect 31944 24550 31996 24556
rect 31956 23186 31984 24550
rect 32036 24132 32088 24138
rect 32036 24074 32088 24080
rect 32048 23746 32076 24074
rect 32140 23866 32168 24754
rect 32128 23860 32180 23866
rect 32128 23802 32180 23808
rect 32048 23718 32168 23746
rect 32036 23316 32088 23322
rect 32036 23258 32088 23264
rect 31944 23180 31996 23186
rect 31944 23122 31996 23128
rect 31944 22976 31996 22982
rect 31944 22918 31996 22924
rect 31956 22098 31984 22918
rect 32048 22642 32076 23258
rect 32036 22636 32088 22642
rect 32036 22578 32088 22584
rect 31944 22092 31996 22098
rect 31944 22034 31996 22040
rect 32048 21554 32076 22578
rect 32036 21548 32088 21554
rect 32036 21490 32088 21496
rect 32140 18698 32168 23718
rect 32232 22982 32260 28494
rect 32324 27130 32352 29038
rect 32508 28762 32536 29038
rect 32496 28756 32548 28762
rect 32496 28698 32548 28704
rect 32312 27124 32364 27130
rect 32312 27066 32364 27072
rect 32324 26382 32352 27066
rect 32404 26920 32456 26926
rect 32404 26862 32456 26868
rect 32416 26586 32444 26862
rect 32404 26580 32456 26586
rect 32404 26522 32456 26528
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32508 25498 32536 25842
rect 32496 25492 32548 25498
rect 32496 25434 32548 25440
rect 32404 24744 32456 24750
rect 32404 24686 32456 24692
rect 32416 24426 32444 24686
rect 32772 24608 32824 24614
rect 32772 24550 32824 24556
rect 32324 24410 32444 24426
rect 32312 24404 32444 24410
rect 32364 24398 32444 24404
rect 32496 24404 32548 24410
rect 32312 24346 32364 24352
rect 32496 24346 32548 24352
rect 32508 23662 32536 24346
rect 32784 24206 32812 24550
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 32784 23730 32812 24142
rect 32864 23860 32916 23866
rect 32864 23802 32916 23808
rect 32772 23724 32824 23730
rect 32772 23666 32824 23672
rect 32496 23656 32548 23662
rect 32496 23598 32548 23604
rect 32784 23322 32812 23666
rect 32772 23316 32824 23322
rect 32772 23258 32824 23264
rect 32312 23044 32364 23050
rect 32312 22986 32364 22992
rect 32220 22976 32272 22982
rect 32220 22918 32272 22924
rect 32324 22778 32352 22986
rect 32312 22772 32364 22778
rect 32312 22714 32364 22720
rect 32220 21956 32272 21962
rect 32220 21898 32272 21904
rect 32232 21690 32260 21898
rect 32876 21894 32904 23802
rect 32864 21888 32916 21894
rect 32864 21830 32916 21836
rect 32220 21684 32272 21690
rect 32220 21626 32272 21632
rect 32968 21486 32996 29582
rect 34532 28218 34560 30262
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34520 28212 34572 28218
rect 34520 28154 34572 28160
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 34152 28008 34204 28014
rect 34152 27950 34204 27956
rect 33152 27606 33180 27950
rect 34164 27674 34192 27950
rect 34152 27668 34204 27674
rect 34152 27610 34204 27616
rect 33140 27600 33192 27606
rect 33140 27542 33192 27548
rect 34152 27532 34204 27538
rect 34152 27474 34204 27480
rect 33140 27056 33192 27062
rect 33140 26998 33192 27004
rect 33152 26042 33180 26998
rect 34060 26988 34112 26994
rect 34060 26930 34112 26936
rect 33968 26920 34020 26926
rect 33968 26862 34020 26868
rect 33980 26382 34008 26862
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 33876 26240 33928 26246
rect 33876 26182 33928 26188
rect 33140 26036 33192 26042
rect 33140 25978 33192 25984
rect 33888 25702 33916 26182
rect 33980 25906 34008 26318
rect 34072 26246 34100 26930
rect 34164 26586 34192 27474
rect 34532 27470 34560 28154
rect 34796 28144 34848 28150
rect 34796 28086 34848 28092
rect 34808 27606 34836 28086
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34796 27600 34848 27606
rect 34796 27542 34848 27548
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 34244 27056 34296 27062
rect 34244 26998 34296 27004
rect 34152 26580 34204 26586
rect 34152 26522 34204 26528
rect 34256 26382 34284 26998
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34428 26444 34480 26450
rect 34428 26386 34480 26392
rect 34244 26376 34296 26382
rect 34244 26318 34296 26324
rect 34060 26240 34112 26246
rect 34060 26182 34112 26188
rect 34072 25974 34100 26182
rect 34060 25968 34112 25974
rect 34060 25910 34112 25916
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 34152 25900 34204 25906
rect 34152 25842 34204 25848
rect 33876 25696 33928 25702
rect 33876 25638 33928 25644
rect 33968 25152 34020 25158
rect 33968 25094 34020 25100
rect 33876 24812 33928 24818
rect 33876 24754 33928 24760
rect 33232 24336 33284 24342
rect 33232 24278 33284 24284
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33152 23866 33180 24142
rect 33244 24070 33272 24278
rect 33600 24132 33652 24138
rect 33600 24074 33652 24080
rect 33232 24064 33284 24070
rect 33232 24006 33284 24012
rect 33244 23866 33272 24006
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 33232 23860 33284 23866
rect 33232 23802 33284 23808
rect 33612 23730 33640 24074
rect 33888 24070 33916 24754
rect 33980 24750 34008 25094
rect 34164 24750 34192 25842
rect 34256 25702 34284 26318
rect 34440 25974 34468 26386
rect 34704 26376 34756 26382
rect 34704 26318 34756 26324
rect 34716 26042 34744 26318
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 34428 25968 34480 25974
rect 34428 25910 34480 25916
rect 34440 25702 34468 25910
rect 34808 25906 34836 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34980 26308 35032 26314
rect 34980 26250 35032 26256
rect 34992 26042 35020 26250
rect 34980 26036 35032 26042
rect 34980 25978 35032 25984
rect 35164 25968 35216 25974
rect 35164 25910 35216 25916
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 35176 25770 35204 25910
rect 35164 25764 35216 25770
rect 35164 25706 35216 25712
rect 34244 25696 34296 25702
rect 34244 25638 34296 25644
rect 34428 25696 34480 25702
rect 34428 25638 34480 25644
rect 34520 25696 34572 25702
rect 34520 25638 34572 25644
rect 34256 24954 34284 25638
rect 34532 25226 34560 25638
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 34244 24948 34296 24954
rect 34244 24890 34296 24896
rect 34244 24812 34296 24818
rect 34244 24754 34296 24760
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 34152 24744 34204 24750
rect 34152 24686 34204 24692
rect 34164 24342 34192 24686
rect 34256 24410 34284 24754
rect 35256 24744 35308 24750
rect 34808 24704 35256 24732
rect 34808 24614 34836 24704
rect 35256 24686 35308 24692
rect 34796 24608 34848 24614
rect 34796 24550 34848 24556
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34244 24404 34296 24410
rect 34244 24346 34296 24352
rect 34152 24336 34204 24342
rect 34152 24278 34204 24284
rect 35256 24336 35308 24342
rect 35256 24278 35308 24284
rect 33876 24064 33928 24070
rect 33876 24006 33928 24012
rect 33600 23724 33652 23730
rect 33600 23666 33652 23672
rect 33876 23520 33928 23526
rect 33876 23462 33928 23468
rect 33888 23118 33916 23462
rect 34164 23118 34192 24278
rect 34244 24200 34296 24206
rect 34244 24142 34296 24148
rect 34256 23118 34284 24142
rect 35268 23798 35296 24278
rect 35256 23792 35308 23798
rect 35256 23734 35308 23740
rect 34612 23656 34664 23662
rect 34612 23598 34664 23604
rect 34624 23186 34652 23598
rect 34704 23520 34756 23526
rect 34704 23462 34756 23468
rect 34716 23322 34744 23462
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34704 23316 34756 23322
rect 34704 23258 34756 23264
rect 34612 23180 34664 23186
rect 34612 23122 34664 23128
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 34152 23112 34204 23118
rect 34152 23054 34204 23060
rect 34244 23112 34296 23118
rect 34244 23054 34296 23060
rect 34704 23112 34756 23118
rect 34704 23054 34756 23060
rect 34716 22710 34744 23054
rect 34704 22704 34756 22710
rect 34704 22646 34756 22652
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35452 22234 35480 47466
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38396 45554 38424 49286
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49314 40030 50000
rect 39500 49286 40030 49314
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 39500 45554 39528 49286
rect 39918 49200 40030 49286
rect 40562 49200 40674 50000
rect 41206 49200 41318 50000
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 40132 47456 40184 47462
rect 40132 47398 40184 47404
rect 39948 46096 40000 46102
rect 39948 46038 40000 46044
rect 39960 45966 39988 46038
rect 39948 45960 40000 45966
rect 39948 45902 40000 45908
rect 38396 45526 38608 45554
rect 35532 27464 35584 27470
rect 35532 27406 35584 27412
rect 35544 25906 35572 27406
rect 36636 26376 36688 26382
rect 36636 26318 36688 26324
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 36004 26042 36032 26250
rect 35992 26036 36044 26042
rect 35992 25978 36044 25984
rect 35532 25900 35584 25906
rect 35532 25842 35584 25848
rect 35544 25498 35572 25842
rect 36268 25832 36320 25838
rect 36452 25832 36504 25838
rect 36320 25792 36452 25820
rect 36268 25774 36320 25780
rect 36452 25774 36504 25780
rect 35532 25492 35584 25498
rect 35532 25434 35584 25440
rect 35544 24206 35572 25434
rect 36268 24812 36320 24818
rect 36268 24754 36320 24760
rect 36280 24410 36308 24754
rect 36648 24750 36676 26318
rect 37648 26308 37700 26314
rect 37648 26250 37700 26256
rect 37660 26042 37688 26250
rect 37648 26036 37700 26042
rect 37648 25978 37700 25984
rect 37556 25900 37608 25906
rect 37556 25842 37608 25848
rect 37568 25430 37596 25842
rect 37556 25424 37608 25430
rect 37556 25366 37608 25372
rect 36636 24744 36688 24750
rect 36636 24686 36688 24692
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 38580 24274 38608 45526
rect 38672 45526 39528 45554
rect 38672 44810 38700 45526
rect 38660 44804 38712 44810
rect 38660 44746 38712 44752
rect 39960 38418 39988 45902
rect 39120 38412 39172 38418
rect 39120 38354 39172 38360
rect 39948 38412 40000 38418
rect 39948 38354 40000 38360
rect 39132 25294 39160 38354
rect 40040 25492 40092 25498
rect 40040 25434 40092 25440
rect 39396 25424 39448 25430
rect 39396 25366 39448 25372
rect 39120 25288 39172 25294
rect 39120 25230 39172 25236
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 38764 24410 38792 24754
rect 39028 24608 39080 24614
rect 39028 24550 39080 24556
rect 38752 24404 38804 24410
rect 38752 24346 38804 24352
rect 38568 24268 38620 24274
rect 38568 24210 38620 24216
rect 35532 24200 35584 24206
rect 35532 24142 35584 24148
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 36096 23866 36124 24142
rect 37372 24132 37424 24138
rect 37372 24074 37424 24080
rect 38568 24132 38620 24138
rect 38568 24074 38620 24080
rect 37384 23866 37412 24074
rect 36084 23860 36136 23866
rect 36084 23802 36136 23808
rect 37372 23860 37424 23866
rect 37372 23802 37424 23808
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 37292 22098 37320 23666
rect 37280 22092 37332 22098
rect 37280 22034 37332 22040
rect 35900 22024 35952 22030
rect 35900 21966 35952 21972
rect 34612 21888 34664 21894
rect 34612 21830 34664 21836
rect 34624 21554 34652 21830
rect 35256 21616 35308 21622
rect 35256 21558 35308 21564
rect 34612 21548 34664 21554
rect 34612 21490 34664 21496
rect 32956 21480 33008 21486
rect 32956 21422 33008 21428
rect 35268 21418 35296 21558
rect 35256 21412 35308 21418
rect 35256 21354 35308 21360
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35912 20874 35940 21966
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36188 21010 36216 21422
rect 36176 21004 36228 21010
rect 36176 20946 36228 20952
rect 35532 20868 35584 20874
rect 35532 20810 35584 20816
rect 35900 20868 35952 20874
rect 35900 20810 35952 20816
rect 36360 20868 36412 20874
rect 36360 20810 36412 20816
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 33232 20256 33284 20262
rect 33232 20198 33284 20204
rect 32220 19984 32272 19990
rect 32220 19926 32272 19932
rect 32232 19446 32260 19926
rect 33244 19786 33272 20198
rect 32312 19780 32364 19786
rect 32312 19722 32364 19728
rect 33232 19780 33284 19786
rect 33232 19722 33284 19728
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 32232 18766 32260 19382
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 32128 18692 32180 18698
rect 32128 18634 32180 18640
rect 32048 18290 32076 18634
rect 32220 18352 32272 18358
rect 32220 18294 32272 18300
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 32232 18086 32260 18294
rect 32220 18080 32272 18086
rect 32220 18022 32272 18028
rect 32220 15428 32272 15434
rect 32220 15370 32272 15376
rect 32036 5160 32088 5166
rect 32036 5102 32088 5108
rect 32048 2530 32076 5102
rect 32232 3670 32260 15370
rect 32324 4826 32352 19722
rect 33428 18970 33456 20402
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34152 19780 34204 19786
rect 34152 19722 34204 19728
rect 33600 19508 33652 19514
rect 33600 19450 33652 19456
rect 33612 19242 33640 19450
rect 34164 19310 34192 19722
rect 35544 19310 35572 20810
rect 34152 19304 34204 19310
rect 34152 19246 34204 19252
rect 35532 19304 35584 19310
rect 35532 19246 35584 19252
rect 33600 19236 33652 19242
rect 33600 19178 33652 19184
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 33140 18964 33192 18970
rect 33140 18906 33192 18912
rect 33416 18964 33468 18970
rect 33416 18906 33468 18912
rect 32864 18692 32916 18698
rect 32864 18634 32916 18640
rect 32404 18080 32456 18086
rect 32404 18022 32456 18028
rect 32416 17610 32444 18022
rect 32876 17610 32904 18634
rect 32404 17604 32456 17610
rect 32404 17546 32456 17552
rect 32864 17604 32916 17610
rect 32864 17546 32916 17552
rect 32876 17270 32904 17546
rect 32864 17264 32916 17270
rect 32864 17206 32916 17212
rect 32312 4820 32364 4826
rect 32312 4762 32364 4768
rect 32876 3738 32904 17206
rect 32864 3732 32916 3738
rect 32864 3674 32916 3680
rect 32220 3664 32272 3670
rect 32220 3606 32272 3612
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 32128 3120 32180 3126
rect 32128 3062 32180 3068
rect 32140 2650 32168 3062
rect 32232 3058 32260 3470
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32416 3126 32444 3334
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32220 3052 32272 3058
rect 32220 2994 32272 3000
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 32048 2502 32260 2530
rect 33152 2514 33180 18906
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 31852 2304 31904 2310
rect 31852 2246 31904 2252
rect 32232 800 32260 2502
rect 33140 2508 33192 2514
rect 33140 2450 33192 2456
rect 33520 800 33548 2858
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 36096 800 36124 2314
rect 36188 2038 36216 2790
rect 36372 2650 36400 20810
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36556 19378 36584 19654
rect 36544 19372 36596 19378
rect 36544 19314 36596 19320
rect 37556 19304 37608 19310
rect 37556 19246 37608 19252
rect 36544 17808 36596 17814
rect 36544 17750 36596 17756
rect 36556 17338 36584 17750
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 37004 4548 37056 4554
rect 37004 4490 37056 4496
rect 37016 4282 37044 4490
rect 37004 4276 37056 4282
rect 37004 4218 37056 4224
rect 36728 4140 36780 4146
rect 36728 4082 36780 4088
rect 36740 3194 36768 4082
rect 37568 4078 37596 19246
rect 38580 4690 38608 24074
rect 38764 17746 38792 24346
rect 39040 23798 39068 24550
rect 39028 23792 39080 23798
rect 39028 23734 39080 23740
rect 38752 17740 38804 17746
rect 38752 17682 38804 17688
rect 39132 16726 39160 25230
rect 39408 24818 39436 25366
rect 40052 25226 40080 25434
rect 40040 25220 40092 25226
rect 40040 25162 40092 25168
rect 39396 24812 39448 24818
rect 39396 24754 39448 24760
rect 38660 16720 38712 16726
rect 38660 16662 38712 16668
rect 39120 16720 39172 16726
rect 39120 16662 39172 16668
rect 38672 16114 38700 16662
rect 38660 16108 38712 16114
rect 38660 16050 38712 16056
rect 38568 4684 38620 4690
rect 38568 4626 38620 4632
rect 38580 4214 38608 4626
rect 38660 4548 38712 4554
rect 38660 4490 38712 4496
rect 37648 4208 37700 4214
rect 37648 4150 37700 4156
rect 38568 4208 38620 4214
rect 38568 4150 38620 4156
rect 37556 4072 37608 4078
rect 37556 4014 37608 4020
rect 37568 3602 37596 4014
rect 37556 3596 37608 3602
rect 37556 3538 37608 3544
rect 37660 3398 37688 4150
rect 38476 3936 38528 3942
rect 38476 3878 38528 3884
rect 38488 3534 38516 3878
rect 38672 3738 38700 4490
rect 39408 3738 39436 24754
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 40052 22778 40080 23054
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40144 22438 40172 47398
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 40420 31958 40448 46922
rect 41248 45554 41276 49200
rect 41696 47252 41748 47258
rect 41696 47194 41748 47200
rect 41328 46368 41380 46374
rect 41328 46310 41380 46316
rect 41340 46034 41368 46310
rect 41328 46028 41380 46034
rect 41328 45970 41380 45976
rect 41512 45892 41564 45898
rect 41512 45834 41564 45840
rect 41524 45626 41552 45834
rect 41512 45620 41564 45626
rect 41512 45562 41564 45568
rect 41248 45526 41368 45554
rect 41236 43240 41288 43246
rect 41236 43182 41288 43188
rect 40408 31952 40460 31958
rect 40408 31894 40460 31900
rect 41248 31754 41276 43182
rect 41156 31726 41276 31754
rect 40776 24336 40828 24342
rect 40776 24278 40828 24284
rect 40788 23866 40816 24278
rect 40776 23860 40828 23866
rect 40776 23802 40828 23808
rect 40500 23656 40552 23662
rect 40500 23598 40552 23604
rect 40512 23526 40540 23598
rect 40500 23520 40552 23526
rect 40500 23462 40552 23468
rect 40512 23186 40540 23462
rect 40500 23180 40552 23186
rect 40500 23122 40552 23128
rect 40316 22636 40368 22642
rect 40316 22578 40368 22584
rect 40132 22432 40184 22438
rect 40132 22374 40184 22380
rect 40144 22098 40172 22374
rect 40132 22092 40184 22098
rect 40132 22034 40184 22040
rect 40328 22030 40356 22578
rect 40316 22024 40368 22030
rect 40500 22024 40552 22030
rect 40368 21972 40500 21978
rect 40316 21966 40552 21972
rect 40328 21950 40540 21966
rect 40408 21888 40460 21894
rect 40408 21830 40460 21836
rect 40316 5024 40368 5030
rect 40316 4966 40368 4972
rect 40328 4758 40356 4966
rect 40316 4752 40368 4758
rect 40316 4694 40368 4700
rect 40040 4480 40092 4486
rect 40040 4422 40092 4428
rect 40132 4480 40184 4486
rect 40132 4422 40184 4428
rect 40052 4214 40080 4422
rect 40040 4208 40092 4214
rect 40040 4150 40092 4156
rect 40040 4072 40092 4078
rect 39592 4010 39804 4026
rect 40144 4026 40172 4422
rect 40092 4020 40172 4026
rect 40040 4014 40172 4020
rect 40316 4072 40368 4078
rect 40316 4014 40368 4020
rect 39580 4004 39816 4010
rect 39632 3998 39764 4004
rect 39580 3946 39632 3952
rect 40052 3998 40172 4014
rect 39764 3946 39816 3952
rect 38660 3732 38712 3738
rect 38660 3674 38712 3680
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 40328 3670 40356 4014
rect 40316 3664 40368 3670
rect 40316 3606 40368 3612
rect 38476 3528 38528 3534
rect 38476 3470 38528 3476
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 37648 3392 37700 3398
rect 37648 3334 37700 3340
rect 36728 3188 36780 3194
rect 36728 3130 36780 3136
rect 37660 3058 37688 3334
rect 39316 3194 39344 3470
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39960 3058 39988 3470
rect 40420 3194 40448 21830
rect 41156 18970 41184 31726
rect 41236 24744 41288 24750
rect 41340 24732 41368 45526
rect 41420 45484 41472 45490
rect 41420 45426 41472 45432
rect 41432 44334 41460 45426
rect 41420 44328 41472 44334
rect 41420 44270 41472 44276
rect 41432 25974 41460 44270
rect 41420 25968 41472 25974
rect 41420 25910 41472 25916
rect 41512 25900 41564 25906
rect 41512 25842 41564 25848
rect 41524 25702 41552 25842
rect 41512 25696 41564 25702
rect 41512 25638 41564 25644
rect 41288 24704 41368 24732
rect 41236 24686 41288 24692
rect 41236 24064 41288 24070
rect 41236 24006 41288 24012
rect 41248 23662 41276 24006
rect 41236 23656 41288 23662
rect 41236 23598 41288 23604
rect 41328 19236 41380 19242
rect 41328 19178 41380 19184
rect 41144 18964 41196 18970
rect 41144 18906 41196 18912
rect 41156 18290 41184 18906
rect 41340 18358 41368 19178
rect 41328 18352 41380 18358
rect 41328 18294 41380 18300
rect 41144 18284 41196 18290
rect 41144 18226 41196 18232
rect 41420 17740 41472 17746
rect 41420 17682 41472 17688
rect 41432 16998 41460 17682
rect 41420 16992 41472 16998
rect 41420 16934 41472 16940
rect 41524 11762 41552 25638
rect 41708 25362 41736 47194
rect 41892 46034 41920 49200
rect 42536 46442 42564 49200
rect 43180 47138 43208 49200
rect 43180 47110 43576 47138
rect 42708 47048 42760 47054
rect 42708 46990 42760 46996
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 42628 46170 42656 46446
rect 42616 46164 42668 46170
rect 42616 46106 42668 46112
rect 41880 46028 41932 46034
rect 41880 45970 41932 45976
rect 42720 45554 42748 46990
rect 43352 46980 43404 46986
rect 43352 46922 43404 46928
rect 42800 45554 42852 45558
rect 42720 45552 42852 45554
rect 42720 45526 42800 45552
rect 42800 45494 42852 45500
rect 42800 45416 42852 45422
rect 42800 45358 42852 45364
rect 42812 45082 42840 45358
rect 42800 45076 42852 45082
rect 42800 45018 42852 45024
rect 43076 30796 43128 30802
rect 43076 30738 43128 30744
rect 42156 26240 42208 26246
rect 42156 26182 42208 26188
rect 42168 25362 42196 26182
rect 42340 25696 42392 25702
rect 42340 25638 42392 25644
rect 42352 25362 42380 25638
rect 41696 25356 41748 25362
rect 41696 25298 41748 25304
rect 42156 25356 42208 25362
rect 42156 25298 42208 25304
rect 42340 25356 42392 25362
rect 42340 25298 42392 25304
rect 42984 24200 43036 24206
rect 42984 24142 43036 24148
rect 42524 23724 42576 23730
rect 42524 23666 42576 23672
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42536 22506 42564 23666
rect 42812 22642 42840 23666
rect 42996 22778 43024 24142
rect 42984 22772 43036 22778
rect 42984 22714 43036 22720
rect 42800 22636 42852 22642
rect 42800 22578 42852 22584
rect 42524 22500 42576 22506
rect 42524 22442 42576 22448
rect 42616 20800 42668 20806
rect 42616 20742 42668 20748
rect 42628 20466 42656 20742
rect 42812 20466 42840 22578
rect 43088 21622 43116 30738
rect 43364 30598 43392 46922
rect 43548 45554 43576 47110
rect 43824 47054 43852 49200
rect 44468 47122 44496 49200
rect 44456 47116 44508 47122
rect 44456 47058 44508 47064
rect 43812 47048 43864 47054
rect 43812 46990 43864 46996
rect 45112 45830 45140 49200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 45824 45152 45830
rect 45100 45766 45152 45772
rect 43548 45526 44128 45554
rect 44100 45422 44128 45526
rect 44088 45416 44140 45422
rect 44088 45358 44140 45364
rect 45100 45416 45152 45422
rect 45100 45358 45152 45364
rect 43536 45348 43588 45354
rect 43536 45290 43588 45296
rect 43548 45082 43576 45290
rect 45112 45082 45140 45358
rect 43536 45076 43588 45082
rect 43536 45018 43588 45024
rect 45100 45076 45152 45082
rect 45100 45018 45152 45024
rect 45008 44872 45060 44878
rect 45008 44814 45060 44820
rect 44364 42288 44416 42294
rect 44364 42230 44416 42236
rect 43628 38956 43680 38962
rect 43628 38898 43680 38904
rect 43640 38350 43668 38898
rect 44376 38894 44404 42230
rect 45020 39438 45048 44814
rect 45204 44402 45232 46990
rect 45468 46980 45520 46986
rect 45468 46922 45520 46928
rect 45376 46504 45428 46510
rect 45376 46446 45428 46452
rect 45388 46170 45416 46446
rect 45376 46164 45428 46170
rect 45376 46106 45428 46112
rect 45376 45892 45428 45898
rect 45376 45834 45428 45840
rect 45388 44878 45416 45834
rect 45376 44872 45428 44878
rect 45376 44814 45428 44820
rect 45192 44396 45244 44402
rect 45192 44338 45244 44344
rect 45388 42294 45416 44814
rect 45480 44470 45508 46922
rect 45652 46436 45704 46442
rect 45652 46378 45704 46384
rect 45664 45880 45692 46378
rect 45756 46034 45784 49200
rect 45744 46028 45796 46034
rect 45744 45970 45796 45976
rect 46296 45960 46348 45966
rect 46296 45902 46348 45908
rect 45836 45892 45888 45898
rect 45664 45852 45784 45880
rect 45560 45824 45612 45830
rect 45612 45784 45692 45812
rect 45560 45766 45612 45772
rect 45664 45422 45692 45784
rect 45652 45416 45704 45422
rect 45652 45358 45704 45364
rect 45468 44464 45520 44470
rect 45468 44406 45520 44412
rect 45756 44402 45784 45852
rect 45836 45834 45888 45840
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45376 42288 45428 42294
rect 45376 42230 45428 42236
rect 45848 40118 45876 45834
rect 46308 45014 46336 45902
rect 46400 45626 46428 49200
rect 46754 47696 46810 47705
rect 46754 47631 46810 47640
rect 46768 46510 46796 47631
rect 46848 47252 46900 47258
rect 46848 47194 46900 47200
rect 46860 47025 46888 47194
rect 46846 47016 46902 47025
rect 46846 46951 46902 46960
rect 46756 46504 46808 46510
rect 46756 46446 46808 46452
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 47860 47184 47912 47190
rect 47860 47126 47912 47132
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46388 45620 46440 45626
rect 46388 45562 46440 45568
rect 46492 45082 46520 45834
rect 47492 45280 47544 45286
rect 47492 45222 47544 45228
rect 46480 45076 46532 45082
rect 46480 45018 46532 45024
rect 46296 45008 46348 45014
rect 46296 44950 46348 44956
rect 46204 44804 46256 44810
rect 46204 44746 46256 44752
rect 46480 44804 46532 44810
rect 46480 44746 46532 44752
rect 46216 42226 46244 44746
rect 46492 44538 46520 44746
rect 47032 44736 47084 44742
rect 47032 44678 47084 44684
rect 46480 44532 46532 44538
rect 46480 44474 46532 44480
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 46952 43858 46980 44134
rect 46940 43852 46992 43858
rect 46940 43794 46992 43800
rect 47044 43314 47072 44678
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 46940 42628 46992 42634
rect 46940 42570 46992 42576
rect 46952 42362 46980 42570
rect 46940 42356 46992 42362
rect 46940 42298 46992 42304
rect 46204 42220 46256 42226
rect 46204 42162 46256 42168
rect 46664 42220 46716 42226
rect 46664 42162 46716 42168
rect 46480 42016 46532 42022
rect 46480 41958 46532 41964
rect 46492 41682 46520 41958
rect 46480 41676 46532 41682
rect 46480 41618 46532 41624
rect 45836 40112 45888 40118
rect 45836 40054 45888 40060
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 45008 39432 45060 39438
rect 45008 39374 45060 39380
rect 44364 38888 44416 38894
rect 44364 38830 44416 38836
rect 44640 38888 44692 38894
rect 44640 38830 44692 38836
rect 43628 38344 43680 38350
rect 43628 38286 43680 38292
rect 43640 37874 43668 38286
rect 43628 37868 43680 37874
rect 43628 37810 43680 37816
rect 44272 37868 44324 37874
rect 44272 37810 44324 37816
rect 44284 37466 44312 37810
rect 44272 37460 44324 37466
rect 44272 37402 44324 37408
rect 44284 37262 44312 37402
rect 44088 37256 44140 37262
rect 44088 37198 44140 37204
rect 44272 37256 44324 37262
rect 44272 37198 44324 37204
rect 44100 36854 44128 37198
rect 44088 36848 44140 36854
rect 44088 36790 44140 36796
rect 44376 35894 44404 38830
rect 44376 35866 44588 35894
rect 43352 30592 43404 30598
rect 43352 30534 43404 30540
rect 43720 27668 43772 27674
rect 43720 27610 43772 27616
rect 43732 26450 43760 27610
rect 43720 26444 43772 26450
rect 43720 26386 43772 26392
rect 43996 25220 44048 25226
rect 43996 25162 44048 25168
rect 43168 24200 43220 24206
rect 43168 24142 43220 24148
rect 43180 23322 43208 24142
rect 43536 24064 43588 24070
rect 43536 24006 43588 24012
rect 43548 23730 43576 24006
rect 43536 23724 43588 23730
rect 43536 23666 43588 23672
rect 43168 23316 43220 23322
rect 43168 23258 43220 23264
rect 43444 23180 43496 23186
rect 43444 23122 43496 23128
rect 43456 22642 43484 23122
rect 43536 23112 43588 23118
rect 43536 23054 43588 23060
rect 43444 22636 43496 22642
rect 43444 22578 43496 22584
rect 43548 22574 43576 23054
rect 43720 22976 43772 22982
rect 43720 22918 43772 22924
rect 43732 22778 43760 22918
rect 43720 22772 43772 22778
rect 43720 22714 43772 22720
rect 43536 22568 43588 22574
rect 43536 22510 43588 22516
rect 43260 22024 43312 22030
rect 43444 22024 43496 22030
rect 43260 21966 43312 21972
rect 43364 21972 43444 21978
rect 43364 21966 43496 21972
rect 43076 21616 43128 21622
rect 43076 21558 43128 21564
rect 42892 21548 42944 21554
rect 42892 21490 42944 21496
rect 42904 20942 42932 21490
rect 43088 21078 43116 21558
rect 43168 21344 43220 21350
rect 43168 21286 43220 21292
rect 43076 21072 43128 21078
rect 42996 21020 43076 21026
rect 42996 21014 43128 21020
rect 42996 20998 43116 21014
rect 42892 20936 42944 20942
rect 42892 20878 42944 20884
rect 42616 20460 42668 20466
rect 42616 20402 42668 20408
rect 42800 20460 42852 20466
rect 42800 20402 42852 20408
rect 42904 19922 42932 20878
rect 42892 19916 42944 19922
rect 42892 19858 42944 19864
rect 42996 19854 43024 20998
rect 43076 20936 43128 20942
rect 43076 20878 43128 20884
rect 43088 20602 43116 20878
rect 43076 20596 43128 20602
rect 43076 20538 43128 20544
rect 43180 20398 43208 21286
rect 43272 20466 43300 21966
rect 43364 21950 43484 21966
rect 43364 20602 43392 21950
rect 43444 21888 43496 21894
rect 43444 21830 43496 21836
rect 43456 20942 43484 21830
rect 43444 20936 43496 20942
rect 43444 20878 43496 20884
rect 43352 20596 43404 20602
rect 43352 20538 43404 20544
rect 43260 20460 43312 20466
rect 43260 20402 43312 20408
rect 43168 20392 43220 20398
rect 43168 20334 43220 20340
rect 43272 20262 43300 20402
rect 43260 20256 43312 20262
rect 43260 20198 43312 20204
rect 43364 19990 43392 20538
rect 43352 19984 43404 19990
rect 43352 19926 43404 19932
rect 42984 19848 43036 19854
rect 42984 19790 43036 19796
rect 43260 19848 43312 19854
rect 43260 19790 43312 19796
rect 42800 19168 42852 19174
rect 42800 19110 42852 19116
rect 42812 18834 42840 19110
rect 42800 18828 42852 18834
rect 42800 18770 42852 18776
rect 41604 18148 41656 18154
rect 41604 18090 41656 18096
rect 41616 17746 41644 18090
rect 42616 17876 42668 17882
rect 42616 17818 42668 17824
rect 41604 17740 41656 17746
rect 41604 17682 41656 17688
rect 41880 17740 41932 17746
rect 41880 17682 41932 17688
rect 41892 17270 41920 17682
rect 41880 17264 41932 17270
rect 41880 17206 41932 17212
rect 42248 16992 42300 16998
rect 42248 16934 42300 16940
rect 42260 16046 42288 16934
rect 42628 16658 42656 17818
rect 42616 16652 42668 16658
rect 42616 16594 42668 16600
rect 42892 16516 42944 16522
rect 42892 16458 42944 16464
rect 42904 16250 42932 16458
rect 42892 16244 42944 16250
rect 42892 16186 42944 16192
rect 42248 16040 42300 16046
rect 42248 15982 42300 15988
rect 41512 11756 41564 11762
rect 41512 11698 41564 11704
rect 40868 6724 40920 6730
rect 40868 6666 40920 6672
rect 40880 6458 40908 6666
rect 40868 6452 40920 6458
rect 40868 6394 40920 6400
rect 40868 6316 40920 6322
rect 40868 6258 40920 6264
rect 40880 5370 40908 6258
rect 41880 5772 41932 5778
rect 41880 5714 41932 5720
rect 40868 5364 40920 5370
rect 40868 5306 40920 5312
rect 40500 4616 40552 4622
rect 40500 4558 40552 4564
rect 40512 4162 40540 4558
rect 40512 4134 40632 4162
rect 40500 4072 40552 4078
rect 40500 4014 40552 4020
rect 40512 3466 40540 4014
rect 40604 3670 40632 4134
rect 40592 3664 40644 3670
rect 40592 3606 40644 3612
rect 41892 3602 41920 5714
rect 41972 5636 42024 5642
rect 41972 5578 42024 5584
rect 41984 5234 42012 5578
rect 41972 5228 42024 5234
rect 41972 5170 42024 5176
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 41788 3528 41840 3534
rect 41788 3470 41840 3476
rect 40500 3460 40552 3466
rect 40500 3402 40552 3408
rect 40408 3188 40460 3194
rect 40408 3130 40460 3136
rect 37648 3052 37700 3058
rect 37648 2994 37700 3000
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 39132 2650 39160 2994
rect 40420 2854 40448 3130
rect 40512 2938 40540 3402
rect 41420 3392 41472 3398
rect 41420 3334 41472 3340
rect 40512 2910 40632 2938
rect 40604 2854 40632 2910
rect 40408 2848 40460 2854
rect 40408 2790 40460 2796
rect 40592 2848 40644 2854
rect 40592 2790 40644 2796
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 39948 2440 40000 2446
rect 39948 2382 40000 2388
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 36176 2032 36228 2038
rect 36176 1974 36228 1980
rect 38028 800 38056 2382
rect 39396 2372 39448 2378
rect 39396 2314 39448 2320
rect 39408 1170 39436 2314
rect 39316 1142 39436 1170
rect 39316 800 39344 1142
rect 39960 800 39988 2382
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 41248 800 41276 2382
rect 41432 2378 41460 3334
rect 41696 3120 41748 3126
rect 41524 3068 41696 3074
rect 41524 3062 41748 3068
rect 41524 3058 41736 3062
rect 41512 3052 41736 3058
rect 41564 3046 41736 3052
rect 41512 2994 41564 3000
rect 41800 2990 41828 3470
rect 41788 2984 41840 2990
rect 41788 2926 41840 2932
rect 41800 2650 41828 2926
rect 41788 2644 41840 2650
rect 41788 2586 41840 2592
rect 41984 2514 42012 5170
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 42812 3602 42840 3878
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 43168 3596 43220 3602
rect 43168 3538 43220 3544
rect 42524 3460 42576 3466
rect 42524 3402 42576 3408
rect 42432 3392 42484 3398
rect 42432 3334 42484 3340
rect 42444 3058 42472 3334
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 41972 2508 42024 2514
rect 41972 2450 42024 2456
rect 41420 2372 41472 2378
rect 41420 2314 41472 2320
rect 42536 800 42564 3402
rect 43180 800 43208 3538
rect 43272 2310 43300 19790
rect 43548 6866 43576 22510
rect 43628 20460 43680 20466
rect 43628 20402 43680 20408
rect 43640 20058 43668 20402
rect 43812 20392 43864 20398
rect 43812 20334 43864 20340
rect 43824 20058 43852 20334
rect 43628 20052 43680 20058
rect 43628 19994 43680 20000
rect 43812 20052 43864 20058
rect 43812 19994 43864 20000
rect 43720 18284 43772 18290
rect 43720 18226 43772 18232
rect 43732 17542 43760 18226
rect 43720 17536 43772 17542
rect 43720 17478 43772 17484
rect 43720 16448 43772 16454
rect 43720 16390 43772 16396
rect 43732 16250 43760 16390
rect 43720 16244 43772 16250
rect 43720 16186 43772 16192
rect 43536 6860 43588 6866
rect 43536 6802 43588 6808
rect 43548 5778 43576 6802
rect 43536 5772 43588 5778
rect 43536 5714 43588 5720
rect 43812 3936 43864 3942
rect 43812 3878 43864 3884
rect 43824 3670 43852 3878
rect 43812 3664 43864 3670
rect 43812 3606 43864 3612
rect 44008 3466 44036 25162
rect 44364 21888 44416 21894
rect 44364 21830 44416 21836
rect 44376 21554 44404 21830
rect 44560 21570 44588 35866
rect 44652 23662 44680 38830
rect 44916 37800 44968 37806
rect 44916 37742 44968 37748
rect 44928 24818 44956 37742
rect 44916 24812 44968 24818
rect 44916 24754 44968 24760
rect 44928 24410 44956 24754
rect 44916 24404 44968 24410
rect 44916 24346 44968 24352
rect 44640 23656 44692 23662
rect 44640 23598 44692 23604
rect 44652 22098 44680 23598
rect 44640 22092 44692 22098
rect 44640 22034 44692 22040
rect 44364 21548 44416 21554
rect 44560 21542 44864 21570
rect 44364 21490 44416 21496
rect 44640 21480 44692 21486
rect 44640 21422 44692 21428
rect 44272 21344 44324 21350
rect 44272 21286 44324 21292
rect 44088 20800 44140 20806
rect 44088 20742 44140 20748
rect 44100 20346 44128 20742
rect 44284 20534 44312 21286
rect 44364 20868 44416 20874
rect 44364 20810 44416 20816
rect 44272 20528 44324 20534
rect 44272 20470 44324 20476
rect 44376 20482 44404 20810
rect 44376 20466 44588 20482
rect 44364 20460 44588 20466
rect 44416 20454 44588 20460
rect 44364 20402 44416 20408
rect 44456 20392 44508 20398
rect 44100 20340 44456 20346
rect 44100 20334 44508 20340
rect 44100 20318 44496 20334
rect 44100 18698 44128 20318
rect 44180 20052 44232 20058
rect 44180 19994 44232 20000
rect 44088 18692 44140 18698
rect 44088 18634 44140 18640
rect 44192 17882 44220 19994
rect 44560 19922 44588 20454
rect 44652 20058 44680 21422
rect 44732 20936 44784 20942
rect 44732 20878 44784 20884
rect 44744 20466 44772 20878
rect 44732 20460 44784 20466
rect 44732 20402 44784 20408
rect 44640 20052 44692 20058
rect 44640 19994 44692 20000
rect 44744 19938 44772 20402
rect 44548 19916 44600 19922
rect 44548 19858 44600 19864
rect 44652 19910 44772 19938
rect 44652 19854 44680 19910
rect 44640 19848 44692 19854
rect 44640 19790 44692 19796
rect 44456 18692 44508 18698
rect 44456 18634 44508 18640
rect 44364 18624 44416 18630
rect 44364 18566 44416 18572
rect 44376 18290 44404 18566
rect 44364 18284 44416 18290
rect 44364 18226 44416 18232
rect 44364 18148 44416 18154
rect 44364 18090 44416 18096
rect 44180 17876 44232 17882
rect 44180 17818 44232 17824
rect 44272 17536 44324 17542
rect 44272 17478 44324 17484
rect 44284 17270 44312 17478
rect 44272 17264 44324 17270
rect 44272 17206 44324 17212
rect 44376 17134 44404 18090
rect 44364 17128 44416 17134
rect 44364 17070 44416 17076
rect 44088 16448 44140 16454
rect 44088 16390 44140 16396
rect 44100 16182 44128 16390
rect 44088 16176 44140 16182
rect 44088 16118 44140 16124
rect 43996 3460 44048 3466
rect 43996 3402 44048 3408
rect 44468 3126 44496 18634
rect 44548 17128 44600 17134
rect 44548 17070 44600 17076
rect 44560 16794 44588 17070
rect 44548 16788 44600 16794
rect 44548 16730 44600 16736
rect 44652 6458 44680 19790
rect 44836 18426 44864 21542
rect 44824 18420 44876 18426
rect 44824 18362 44876 18368
rect 44640 6452 44692 6458
rect 44640 6394 44692 6400
rect 44928 4146 44956 24346
rect 45020 24138 45048 39374
rect 45192 39296 45244 39302
rect 45192 39238 45244 39244
rect 45204 39030 45232 39238
rect 45192 39024 45244 39030
rect 45192 38966 45244 38972
rect 46572 38344 46624 38350
rect 46572 38286 46624 38292
rect 45928 38276 45980 38282
rect 45928 38218 45980 38224
rect 45940 37942 45968 38218
rect 45928 37936 45980 37942
rect 45928 37878 45980 37884
rect 45468 37324 45520 37330
rect 45468 37266 45520 37272
rect 45480 28082 45508 37266
rect 45744 30660 45796 30666
rect 45744 30602 45796 30608
rect 45558 28656 45614 28665
rect 45558 28591 45614 28600
rect 45468 28076 45520 28082
rect 45468 28018 45520 28024
rect 45572 27674 45600 28591
rect 45560 27668 45612 27674
rect 45560 27610 45612 27616
rect 45466 26616 45522 26625
rect 45466 26551 45522 26560
rect 45480 25838 45508 26551
rect 45468 25832 45520 25838
rect 45468 25774 45520 25780
rect 45192 25288 45244 25294
rect 45192 25230 45244 25236
rect 45008 24132 45060 24138
rect 45008 24074 45060 24080
rect 45204 22642 45232 25230
rect 45652 25220 45704 25226
rect 45652 25162 45704 25168
rect 45664 24818 45692 25162
rect 45652 24812 45704 24818
rect 45652 24754 45704 24760
rect 45560 24676 45612 24682
rect 45560 24618 45612 24624
rect 45572 23905 45600 24618
rect 45558 23896 45614 23905
rect 45558 23831 45614 23840
rect 45756 23746 45784 30602
rect 45834 30016 45890 30025
rect 45834 29951 45890 29960
rect 45848 23866 45876 29951
rect 45836 23860 45888 23866
rect 45836 23802 45888 23808
rect 45572 23718 45784 23746
rect 45376 22976 45428 22982
rect 45376 22918 45428 22924
rect 45388 22710 45416 22918
rect 45376 22704 45428 22710
rect 45376 22646 45428 22652
rect 45192 22636 45244 22642
rect 45192 22578 45244 22584
rect 45100 22024 45152 22030
rect 45100 21966 45152 21972
rect 45112 21146 45140 21966
rect 45204 21622 45232 22578
rect 45376 22432 45428 22438
rect 45376 22374 45428 22380
rect 45388 22098 45416 22374
rect 45376 22092 45428 22098
rect 45376 22034 45428 22040
rect 45192 21616 45244 21622
rect 45192 21558 45244 21564
rect 45100 21140 45152 21146
rect 45100 21082 45152 21088
rect 45008 19984 45060 19990
rect 45008 19926 45060 19932
rect 45020 19378 45048 19926
rect 45008 19372 45060 19378
rect 45008 19314 45060 19320
rect 45020 16726 45048 19314
rect 45192 18760 45244 18766
rect 45192 18702 45244 18708
rect 45376 18760 45428 18766
rect 45376 18702 45428 18708
rect 45204 18426 45232 18702
rect 45192 18420 45244 18426
rect 45192 18362 45244 18368
rect 45204 17746 45232 18362
rect 45192 17740 45244 17746
rect 45192 17682 45244 17688
rect 45388 17678 45416 18702
rect 45376 17672 45428 17678
rect 45376 17614 45428 17620
rect 45388 17338 45416 17614
rect 45376 17332 45428 17338
rect 45376 17274 45428 17280
rect 45008 16720 45060 16726
rect 45008 16662 45060 16668
rect 45100 16040 45152 16046
rect 45100 15982 45152 15988
rect 44916 4140 44968 4146
rect 44916 4082 44968 4088
rect 44456 3120 44508 3126
rect 44456 3062 44508 3068
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43260 2304 43312 2310
rect 43260 2246 43312 2252
rect 43824 800 43852 2382
rect 45112 800 45140 15982
rect 45572 7954 45600 23718
rect 45744 23044 45796 23050
rect 45744 22986 45796 22992
rect 45756 22574 45784 22986
rect 45744 22568 45796 22574
rect 45744 22510 45796 22516
rect 45756 22098 45784 22510
rect 45744 22092 45796 22098
rect 45744 22034 45796 22040
rect 45652 21480 45704 21486
rect 45652 21422 45704 21428
rect 45664 19786 45692 21422
rect 45756 20398 45784 22034
rect 45744 20392 45796 20398
rect 45744 20334 45796 20340
rect 45652 19780 45704 19786
rect 45652 19722 45704 19728
rect 45652 19372 45704 19378
rect 45652 19314 45704 19320
rect 45664 18465 45692 19314
rect 45650 18456 45706 18465
rect 45650 18391 45706 18400
rect 45756 18340 45784 20334
rect 45940 19718 45968 37878
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46308 31890 46336 32846
rect 46480 32224 46532 32230
rect 46480 32166 46532 32172
rect 46492 31890 46520 32166
rect 46296 31884 46348 31890
rect 46296 31826 46348 31832
rect 46480 31884 46532 31890
rect 46480 31826 46532 31832
rect 46110 31376 46166 31385
rect 46110 31311 46166 31320
rect 46124 21690 46152 31311
rect 46388 25424 46440 25430
rect 46388 25366 46440 25372
rect 46296 24608 46348 24614
rect 46296 24550 46348 24556
rect 46308 24274 46336 24550
rect 46296 24268 46348 24274
rect 46296 24210 46348 24216
rect 46400 24154 46428 25366
rect 46308 24126 46428 24154
rect 46308 23186 46336 24126
rect 46584 23526 46612 38286
rect 46676 35894 46704 42162
rect 47308 40928 47360 40934
rect 47308 40870 47360 40876
rect 46846 39536 46902 39545
rect 46846 39471 46902 39480
rect 46860 39030 46888 39471
rect 46940 39364 46992 39370
rect 46940 39306 46992 39312
rect 46848 39024 46900 39030
rect 46848 38966 46900 38972
rect 46952 38554 46980 39306
rect 47032 38752 47084 38758
rect 47032 38694 47084 38700
rect 46940 38548 46992 38554
rect 46940 38490 46992 38496
rect 47044 36854 47072 38694
rect 47032 36848 47084 36854
rect 47032 36790 47084 36796
rect 47216 36780 47268 36786
rect 47216 36722 47268 36728
rect 47228 35894 47256 36722
rect 47320 36394 47348 40870
rect 47504 36718 47532 45222
rect 47584 44396 47636 44402
rect 47584 44338 47636 44344
rect 47492 36712 47544 36718
rect 47492 36654 47544 36660
rect 47320 36366 47532 36394
rect 46676 35866 46888 35894
rect 47228 35866 47440 35894
rect 46664 32428 46716 32434
rect 46664 32370 46716 32376
rect 46676 25498 46704 32370
rect 46860 29646 46888 35866
rect 47124 34944 47176 34950
rect 47124 34886 47176 34892
rect 47136 32978 47164 34886
rect 47216 33312 47268 33318
rect 47216 33254 47268 33260
rect 47124 32972 47176 32978
rect 47124 32914 47176 32920
rect 47228 32842 47256 33254
rect 47216 32836 47268 32842
rect 47216 32778 47268 32784
rect 46848 29640 46900 29646
rect 46900 29588 47256 29594
rect 46848 29582 47256 29588
rect 46860 29566 47256 29582
rect 46860 29517 46888 29566
rect 47032 29504 47084 29510
rect 47032 29446 47084 29452
rect 46940 28552 46992 28558
rect 46940 28494 46992 28500
rect 46952 27606 46980 28494
rect 46940 27600 46992 27606
rect 46940 27542 46992 27548
rect 46846 25936 46902 25945
rect 46756 25900 46808 25906
rect 46846 25871 46902 25880
rect 46756 25842 46808 25848
rect 46664 25492 46716 25498
rect 46664 25434 46716 25440
rect 46572 23520 46624 23526
rect 46572 23462 46624 23468
rect 46768 23225 46796 25842
rect 46860 25362 46888 25871
rect 46848 25356 46900 25362
rect 46848 25298 46900 25304
rect 47044 23882 47072 29446
rect 47124 26920 47176 26926
rect 47124 26862 47176 26868
rect 46860 23854 47072 23882
rect 46860 23662 46888 23854
rect 46940 23724 46992 23730
rect 46940 23666 46992 23672
rect 46848 23656 46900 23662
rect 46848 23598 46900 23604
rect 46860 23526 46888 23598
rect 46848 23520 46900 23526
rect 46848 23462 46900 23468
rect 46754 23216 46810 23225
rect 46296 23180 46348 23186
rect 46754 23151 46810 23160
rect 46296 23122 46348 23128
rect 46202 22536 46258 22545
rect 46202 22471 46258 22480
rect 46112 21684 46164 21690
rect 46112 21626 46164 21632
rect 46216 21554 46244 22471
rect 46952 21690 46980 23666
rect 47032 23520 47084 23526
rect 47032 23462 47084 23468
rect 47044 23254 47072 23462
rect 47032 23248 47084 23254
rect 47032 23190 47084 23196
rect 46940 21684 46992 21690
rect 46940 21626 46992 21632
rect 46204 21548 46256 21554
rect 46204 21490 46256 21496
rect 46296 20936 46348 20942
rect 46296 20878 46348 20884
rect 46308 20058 46336 20878
rect 46296 20052 46348 20058
rect 46296 19994 46348 20000
rect 45928 19712 45980 19718
rect 45928 19654 45980 19660
rect 46296 19440 46348 19446
rect 46296 19382 46348 19388
rect 46204 19372 46256 19378
rect 46204 19314 46256 19320
rect 46216 18766 46244 19314
rect 46204 18760 46256 18766
rect 46204 18702 46256 18708
rect 46308 18714 46336 19382
rect 46952 19310 46980 21626
rect 47136 19446 47164 26862
rect 47228 24818 47256 29566
rect 47308 28076 47360 28082
rect 47308 28018 47360 28024
rect 47216 24812 47268 24818
rect 47216 24754 47268 24760
rect 47216 23724 47268 23730
rect 47216 23666 47268 23672
rect 47228 21078 47256 23666
rect 47216 21072 47268 21078
rect 47216 21014 47268 21020
rect 47228 20806 47256 21014
rect 47216 20800 47268 20806
rect 47216 20742 47268 20748
rect 47216 19780 47268 19786
rect 47216 19722 47268 19728
rect 47124 19440 47176 19446
rect 47124 19382 47176 19388
rect 46940 19304 46992 19310
rect 46940 19246 46992 19252
rect 47032 19236 47084 19242
rect 47032 19178 47084 19184
rect 47044 18766 47072 19178
rect 47136 18834 47164 19382
rect 47228 18970 47256 19722
rect 47216 18964 47268 18970
rect 47216 18906 47268 18912
rect 47124 18828 47176 18834
rect 47124 18770 47176 18776
rect 47320 18766 47348 28018
rect 47412 19990 47440 35866
rect 47504 24342 47532 36366
rect 47596 32434 47624 44338
rect 47768 43104 47820 43110
rect 47768 43046 47820 43052
rect 47780 42770 47808 43046
rect 47768 42764 47820 42770
rect 47768 42706 47820 42712
rect 47676 41540 47728 41546
rect 47676 41482 47728 41488
rect 47688 40730 47716 41482
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47768 38956 47820 38962
rect 47768 38898 47820 38904
rect 47780 38865 47808 38898
rect 47766 38856 47822 38865
rect 47766 38791 47822 38800
rect 47768 37664 47820 37670
rect 47768 37606 47820 37612
rect 47676 37188 47728 37194
rect 47676 37130 47728 37136
rect 47688 36922 47716 37130
rect 47780 37126 47808 37606
rect 47768 37120 47820 37126
rect 47768 37062 47820 37068
rect 47676 36916 47728 36922
rect 47676 36858 47728 36864
rect 47676 36712 47728 36718
rect 47676 36654 47728 36660
rect 47688 35894 47716 36654
rect 47688 35866 47808 35894
rect 47676 32972 47728 32978
rect 47676 32914 47728 32920
rect 47584 32428 47636 32434
rect 47584 32370 47636 32376
rect 47688 30802 47716 32914
rect 47676 30796 47728 30802
rect 47676 30738 47728 30744
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27538 47716 27814
rect 47676 27532 47728 27538
rect 47676 27474 47728 27480
rect 47584 25696 47636 25702
rect 47584 25638 47636 25644
rect 47492 24336 47544 24342
rect 47492 24278 47544 24284
rect 47492 23588 47544 23594
rect 47492 23530 47544 23536
rect 47504 22438 47532 23530
rect 47596 22642 47624 25638
rect 47676 24608 47728 24614
rect 47676 24550 47728 24556
rect 47688 24274 47716 24550
rect 47676 24268 47728 24274
rect 47676 24210 47728 24216
rect 47676 23520 47728 23526
rect 47676 23462 47728 23468
rect 47688 23186 47716 23462
rect 47780 23322 47808 35866
rect 47872 35834 47900 47126
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47964 46345 47992 46514
rect 48044 46368 48096 46374
rect 47950 46336 48006 46345
rect 48044 46310 48096 46316
rect 47950 46271 48006 46280
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47860 35828 47912 35834
rect 47860 35770 47912 35776
rect 47860 34400 47912 34406
rect 47860 34342 47912 34348
rect 47872 33318 47900 34342
rect 47952 33924 48004 33930
rect 47952 33866 48004 33872
rect 47964 33425 47992 33866
rect 47950 33416 48006 33425
rect 47950 33351 48006 33360
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 47952 32428 48004 32434
rect 47952 32370 48004 32376
rect 47964 32065 47992 32370
rect 47950 32056 48006 32065
rect 47950 31991 48006 32000
rect 48056 26926 48084 46310
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48148 37330 48176 38111
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 48136 35080 48188 35086
rect 48136 35022 48188 35028
rect 48148 34785 48176 35022
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48148 34105 48176 34546
rect 48134 34096 48190 34105
rect 48134 34031 48190 34040
rect 48228 33516 48280 33522
rect 48228 33458 48280 33464
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48148 31890 48176 32671
rect 48136 31884 48188 31890
rect 48136 31826 48188 31832
rect 48240 30598 48268 33458
rect 48228 30592 48280 30598
rect 48228 30534 48280 30540
rect 48136 29640 48188 29646
rect 48136 29582 48188 29588
rect 48148 29345 48176 29582
rect 48134 29336 48190 29345
rect 48134 29271 48190 29280
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48044 26920 48096 26926
rect 48044 26862 48096 26868
rect 48240 26738 48268 30534
rect 48056 26710 48268 26738
rect 47952 24812 48004 24818
rect 47952 24754 48004 24760
rect 47964 24052 47992 24754
rect 48056 24154 48084 26710
rect 48226 25256 48282 25265
rect 48226 25191 48282 25200
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48056 24126 48176 24154
rect 47964 24024 48084 24052
rect 47860 23656 47912 23662
rect 47860 23598 47912 23604
rect 47768 23316 47820 23322
rect 47768 23258 47820 23264
rect 47676 23180 47728 23186
rect 47676 23122 47728 23128
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47676 22568 47728 22574
rect 47676 22510 47728 22516
rect 47492 22432 47544 22438
rect 47492 22374 47544 22380
rect 47504 22094 47532 22374
rect 47504 22066 47624 22094
rect 47596 21622 47624 22066
rect 47688 21894 47716 22510
rect 47872 22098 47900 23598
rect 47952 22636 48004 22642
rect 47952 22578 48004 22584
rect 47860 22092 47912 22098
rect 47860 22034 47912 22040
rect 47964 22030 47992 22578
rect 47768 22024 47820 22030
rect 47768 21966 47820 21972
rect 47952 22024 48004 22030
rect 47952 21966 48004 21972
rect 47676 21888 47728 21894
rect 47676 21830 47728 21836
rect 47584 21616 47636 21622
rect 47584 21558 47636 21564
rect 47688 21434 47716 21830
rect 47780 21622 47808 21966
rect 47860 21888 47912 21894
rect 47860 21830 47912 21836
rect 47950 21856 48006 21865
rect 47872 21690 47900 21830
rect 47950 21791 48006 21800
rect 47860 21684 47912 21690
rect 47860 21626 47912 21632
rect 47768 21616 47820 21622
rect 47768 21558 47820 21564
rect 47596 21406 47716 21434
rect 47400 19984 47452 19990
rect 47400 19926 47452 19932
rect 47400 19712 47452 19718
rect 47400 19654 47452 19660
rect 47412 19378 47440 19654
rect 47492 19508 47544 19514
rect 47492 19450 47544 19456
rect 47400 19372 47452 19378
rect 47400 19314 47452 19320
rect 46388 18760 46440 18766
rect 46308 18708 46388 18714
rect 46308 18702 46440 18708
rect 47032 18760 47084 18766
rect 47032 18702 47084 18708
rect 47308 18760 47360 18766
rect 47308 18702 47360 18708
rect 46112 18692 46164 18698
rect 46308 18686 46428 18702
rect 46112 18634 46164 18640
rect 46124 18358 46152 18634
rect 45664 18312 45784 18340
rect 46112 18352 46164 18358
rect 45664 18222 45692 18312
rect 46112 18294 46164 18300
rect 45652 18216 45704 18222
rect 45652 18158 45704 18164
rect 45664 17270 45692 18158
rect 46400 18086 46428 18686
rect 46480 18624 46532 18630
rect 46480 18566 46532 18572
rect 46388 18080 46440 18086
rect 46388 18022 46440 18028
rect 45652 17264 45704 17270
rect 45652 17206 45704 17212
rect 46020 16516 46072 16522
rect 46020 16458 46072 16464
rect 45652 16244 45704 16250
rect 45652 16186 45704 16192
rect 45664 15745 45692 16186
rect 45650 15736 45706 15745
rect 45650 15671 45706 15680
rect 46032 8265 46060 16458
rect 46400 12434 46428 18022
rect 46492 16522 46520 18566
rect 46756 18284 46808 18290
rect 46756 18226 46808 18232
rect 46768 17202 46796 18226
rect 46756 17196 46808 17202
rect 46756 17138 46808 17144
rect 46480 16516 46532 16522
rect 46480 16458 46532 16464
rect 46400 12406 46612 12434
rect 46480 11552 46532 11558
rect 46480 11494 46532 11500
rect 46492 11218 46520 11494
rect 46480 11212 46532 11218
rect 46480 11154 46532 11160
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46018 8256 46074 8265
rect 46018 8191 46074 8200
rect 45560 7948 45612 7954
rect 45560 7890 45612 7896
rect 45572 5846 45600 7890
rect 46296 7744 46348 7750
rect 46296 7686 46348 7692
rect 46308 7410 46336 7686
rect 46296 7404 46348 7410
rect 46296 7346 46348 7352
rect 45560 5840 45612 5846
rect 45560 5782 45612 5788
rect 46308 4690 46336 7346
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 46388 4208 46440 4214
rect 46388 4150 46440 4156
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3602 46336 3878
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 45204 3058 45232 3470
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 46400 800 46428 4150
rect 46584 2514 46612 12406
rect 46768 7954 46796 17138
rect 46940 16720 46992 16726
rect 46940 16662 46992 16668
rect 46952 11762 46980 16662
rect 46940 11756 46992 11762
rect 46940 11698 46992 11704
rect 46756 7948 46808 7954
rect 46756 7890 46808 7896
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46756 4480 46808 4486
rect 46756 4422 46808 4428
rect 46664 4208 46716 4214
rect 46664 4150 46716 4156
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46676 82 46704 4150
rect 46768 3126 46796 4422
rect 46860 4185 46888 4558
rect 46846 4176 46902 4185
rect 46846 4111 46902 4120
rect 47044 3194 47072 18702
rect 47412 18578 47440 19314
rect 47320 18550 47440 18578
rect 47320 12850 47348 18550
rect 47504 18358 47532 19450
rect 47492 18352 47544 18358
rect 47412 18312 47492 18340
rect 47412 17202 47440 18312
rect 47492 18294 47544 18300
rect 47492 17740 47544 17746
rect 47492 17682 47544 17688
rect 47400 17196 47452 17202
rect 47400 17138 47452 17144
rect 47504 15706 47532 17682
rect 47492 15700 47544 15706
rect 47492 15642 47544 15648
rect 47596 15586 47624 21406
rect 47676 20868 47728 20874
rect 47676 20810 47728 20816
rect 47688 19514 47716 20810
rect 47768 20800 47820 20806
rect 47768 20742 47820 20748
rect 47676 19508 47728 19514
rect 47676 19450 47728 19456
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 47688 17338 47716 17546
rect 47676 17332 47728 17338
rect 47676 17274 47728 17280
rect 47780 17218 47808 20742
rect 47964 20534 47992 21791
rect 47952 20528 48004 20534
rect 47952 20470 48004 20476
rect 48056 18766 48084 24024
rect 48148 22094 48176 24126
rect 48240 23186 48268 25191
rect 48228 23180 48280 23186
rect 48228 23122 48280 23128
rect 48148 22066 48268 22094
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48136 19780 48188 19786
rect 48136 19722 48188 19728
rect 48148 19145 48176 19722
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48044 18760 48096 18766
rect 48044 18702 48096 18708
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 47688 17202 47808 17218
rect 47676 17196 47808 17202
rect 47728 17190 47808 17196
rect 47676 17138 47728 17144
rect 47412 15558 47624 15586
rect 47308 12844 47360 12850
rect 47308 12786 47360 12792
rect 47124 8288 47176 8294
rect 47124 8230 47176 8236
rect 47136 7954 47164 8230
rect 47124 7948 47176 7954
rect 47124 7890 47176 7896
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47320 6866 47348 7511
rect 47412 6866 47440 15558
rect 47688 15450 47716 17138
rect 48148 17105 48176 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 47780 16114 47808 16594
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 48148 16425 48176 16458
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47596 15422 47716 15450
rect 47596 12434 47624 15422
rect 47676 13320 47728 13326
rect 47676 13262 47728 13268
rect 47504 12406 47624 12434
rect 47504 10674 47532 12406
rect 47688 12306 47716 13262
rect 47768 12640 47820 12646
rect 47768 12582 47820 12588
rect 47676 12300 47728 12306
rect 47676 12242 47728 12248
rect 47676 12164 47728 12170
rect 47676 12106 47728 12112
rect 47688 11898 47716 12106
rect 47676 11892 47728 11898
rect 47676 11834 47728 11840
rect 47780 11286 47808 12582
rect 48134 12336 48190 12345
rect 48134 12271 48136 12280
rect 48188 12271 48190 12280
rect 48136 12242 48188 12248
rect 47768 11280 47820 11286
rect 47768 11222 47820 11228
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 47492 10668 47544 10674
rect 47492 10610 47544 10616
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 47400 6860 47452 6866
rect 47400 6802 47452 6808
rect 47504 4554 47532 10610
rect 47676 10464 47728 10470
rect 47676 10406 47728 10412
rect 47688 10130 47716 10406
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 47676 10124 47728 10130
rect 47676 10066 47728 10072
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 47858 9616 47914 9625
rect 47858 9551 47860 9560
rect 47912 9551 47914 9560
rect 47860 9522 47912 9528
rect 48240 9450 48268 22066
rect 48228 9444 48280 9450
rect 48228 9386 48280 9392
rect 47766 8936 47822 8945
rect 47766 8871 47768 8880
rect 47820 8871 47822 8880
rect 47768 8842 47820 8848
rect 48136 8492 48188 8498
rect 48136 8434 48188 8440
rect 47584 7812 47636 7818
rect 47584 7754 47636 7760
rect 47596 7546 47624 7754
rect 47584 7540 47636 7546
rect 47584 7482 47636 7488
rect 48148 6905 48176 8434
rect 48134 6896 48190 6905
rect 48134 6831 48190 6840
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 47964 6225 47992 6258
rect 47950 6216 48006 6225
rect 47950 6151 48006 6160
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 47492 4548 47544 4554
rect 47492 4490 47544 4496
rect 47780 3505 47808 5170
rect 47766 3496 47822 3505
rect 47766 3431 47822 3440
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 47032 3188 47084 3194
rect 47032 3130 47084 3136
rect 46756 3120 46808 3126
rect 46756 3062 46808 3068
rect 48320 3052 48372 3058
rect 48320 2994 48372 3000
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 46756 2372 46808 2378
rect 46756 2314 46808 2320
rect 46768 1465 46796 2314
rect 46754 1456 46810 1465
rect 46754 1391 46810 1400
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 46754 96 46810 105
rect 46676 54 46754 82
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48056 785 48084 2382
rect 48332 800 48360 2994
rect 48976 800 49004 3402
rect 48042 776 48098 785
rect 48042 711 48098 720
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1398 47640 1454 47696
rect 3330 46960 3386 47016
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 1398 42880 1454 42936
rect 1582 35400 1638 35456
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 32680 1638 32736
rect 2778 46280 2834 46336
rect 3422 44920 3478 44976
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1858 32000 1914 32056
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 1858 23160 1914 23216
rect 1858 17720 1914 17776
rect 1858 16360 1914 16416
rect 1398 12280 1454 12336
rect 2778 36760 2834 36816
rect 3330 31320 3386 31376
rect 2226 19080 2282 19136
rect 3330 28600 3386 28656
rect 3514 43560 3570 43616
rect 3698 39480 3754 39536
rect 3054 19760 3110 19816
rect 3422 18420 3478 18456
rect 3422 18400 3424 18420
rect 3424 18400 3476 18420
rect 3476 18400 3478 18420
rect 3054 17040 3110 17096
rect 2778 15000 2834 15056
rect 3422 13640 3478 13696
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3238 7520 3294 7576
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4066 10240 4122 10296
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 14370 37732 14426 37768
rect 14370 37712 14372 37732
rect 14372 37712 14424 37732
rect 14424 37712 14426 37732
rect 14462 29180 14464 29200
rect 14464 29180 14516 29200
rect 14516 29180 14518 29200
rect 14462 29144 14518 29180
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3440 4122 3496
rect 3514 1400 3570 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 17314 37868 17370 37904
rect 17314 37848 17316 37868
rect 17316 37848 17368 37868
rect 17368 37848 17370 37868
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 18694 37848 18750 37904
rect 19338 38120 19394 38176
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19246 37884 19248 37904
rect 19248 37884 19300 37904
rect 19300 37884 19302 37904
rect 19246 37848 19302 37884
rect 19338 37748 19346 37768
rect 19346 37748 19394 37768
rect 19338 37712 19394 37748
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19338 33768 19394 33824
rect 18142 29180 18144 29200
rect 18144 29180 18196 29200
rect 18196 29180 18198 29200
rect 18142 29144 18198 29180
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19982 29416 20038 29472
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19890 20476 19892 20496
rect 19892 20476 19944 20496
rect 19944 20476 19946 20496
rect 19890 20440 19946 20476
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20166 37884 20168 37904
rect 20168 37884 20220 37904
rect 20220 37884 20222 37904
rect 20166 37848 20222 37884
rect 20534 38392 20590 38448
rect 20534 37848 20590 37904
rect 20534 30252 20590 30288
rect 20534 30232 20536 30252
rect 20536 30232 20588 30252
rect 20588 30232 20590 30252
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19706 3032 19762 3088
rect 20718 35028 20720 35048
rect 20720 35028 20772 35048
rect 20772 35028 20774 35048
rect 20718 34992 20774 35028
rect 20810 30540 20812 30560
rect 20812 30540 20864 30560
rect 20864 30540 20866 30560
rect 20810 30504 20866 30540
rect 21086 27820 21088 27840
rect 21088 27820 21140 27840
rect 21140 27820 21142 27840
rect 21086 27784 21142 27820
rect 23110 37712 23166 37768
rect 23570 35708 23572 35728
rect 23572 35708 23624 35728
rect 23624 35708 23626 35728
rect 23570 35672 23626 35708
rect 21822 3032 21878 3088
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22190 2916 22246 2952
rect 22190 2896 22192 2916
rect 22192 2896 22244 2916
rect 22244 2896 22246 2916
rect 23754 27784 23810 27840
rect 23294 20712 23350 20768
rect 23202 20440 23258 20496
rect 23570 20712 23626 20768
rect 22742 3576 22798 3632
rect 22558 3304 22614 3360
rect 24950 29416 25006 29472
rect 26238 35692 26294 35728
rect 26238 35672 26240 35692
rect 26240 35672 26292 35692
rect 26292 35672 26294 35692
rect 25226 3596 25282 3632
rect 25226 3576 25228 3596
rect 25228 3576 25280 3596
rect 25280 3576 25282 3596
rect 25778 29008 25834 29064
rect 27434 37612 27436 37632
rect 27436 37612 27488 37632
rect 27488 37612 27490 37632
rect 27434 37576 27490 37612
rect 25962 30252 26018 30288
rect 25962 30232 25964 30252
rect 25964 30232 26016 30252
rect 26016 30232 26018 30252
rect 27526 34992 27582 35048
rect 26882 30504 26938 30560
rect 26974 29028 27030 29064
rect 26974 29008 26976 29028
rect 26976 29008 27028 29028
rect 27028 29008 27030 29028
rect 26146 2896 26202 2952
rect 27434 3340 27436 3360
rect 27436 3340 27488 3360
rect 27488 3340 27490 3360
rect 27434 3304 27490 3340
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 46754 47640 46810 47696
rect 46846 46960 46902 47016
rect 45558 28600 45614 28656
rect 45466 26560 45522 26616
rect 45558 23840 45614 23896
rect 45834 29960 45890 30016
rect 45650 18400 45706 18456
rect 46110 31320 46166 31376
rect 46846 39480 46902 39536
rect 46846 25880 46902 25936
rect 46754 23160 46810 23216
rect 46202 22480 46258 22536
rect 47766 38800 47822 38856
rect 47950 46280 48006 46336
rect 47950 40840 48006 40896
rect 47950 33360 48006 33416
rect 47950 32000 48006 32056
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48134 34040 48190 34096
rect 48134 32680 48190 32736
rect 48134 29280 48190 29336
rect 48134 27920 48190 27976
rect 48226 25200 48282 25256
rect 48134 24520 48190 24576
rect 47950 21800 48006 21856
rect 45650 15680 45706 15736
rect 46018 8200 46074 8256
rect 2870 720 2926 776
rect 46846 4120 46902 4176
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 47306 7520 47362 7576
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12300 48190 12336
rect 48134 12280 48136 12300
rect 48136 12280 48188 12300
rect 48188 12280 48190 12300
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 47858 9580 47914 9616
rect 47858 9560 47860 9580
rect 47860 9560 47912 9580
rect 47912 9560 47914 9580
rect 47766 8900 47822 8936
rect 47766 8880 47768 8900
rect 47768 8880 47820 8900
rect 47820 8880 47822 8900
rect 48134 6840 48190 6896
rect 47950 6160 48006 6216
rect 47766 3440 47822 3496
rect 46754 1400 46810 1456
rect 46754 40 46810 96
rect 48042 720 48098 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47548 800 47638
rect 1393 47635 1459 47638
rect 46749 47698 46815 47701
rect 49200 47698 50000 47788
rect 46749 47696 50000 47698
rect 46749 47640 46754 47696
rect 46810 47640 50000 47696
rect 46749 47638 50000 47640
rect 46749 47635 46815 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3325 47018 3391 47021
rect 0 47016 3391 47018
rect 0 46960 3330 47016
rect 3386 46960 3391 47016
rect 0 46958 3391 46960
rect 0 46868 800 46958
rect 3325 46955 3391 46958
rect 46841 47018 46907 47021
rect 49200 47018 50000 47108
rect 46841 47016 50000 47018
rect 46841 46960 46846 47016
rect 46902 46960 50000 47016
rect 46841 46958 50000 46960
rect 46841 46955 46907 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3417 44978 3483 44981
rect 0 44976 3483 44978
rect 0 44920 3422 44976
rect 3478 44920 3483 44976
rect 0 44918 3483 44920
rect 0 44828 800 44918
rect 3417 44915 3483 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3509 43618 3575 43621
rect 0 43616 3575 43618
rect 0 43560 3514 43616
rect 3570 43560 3575 43616
rect 0 43558 3575 43560
rect 0 43468 800 43558
rect 3509 43555 3575 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3693 39538 3759 39541
rect 0 39536 3759 39538
rect 0 39480 3698 39536
rect 3754 39480 3759 39536
rect 0 39478 3759 39480
rect 0 39388 800 39478
rect 3693 39475 3759 39478
rect 46841 39538 46907 39541
rect 49200 39538 50000 39628
rect 46841 39536 50000 39538
rect 46841 39480 46846 39536
rect 46902 39480 50000 39536
rect 46841 39478 50000 39480
rect 46841 39475 46907 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47761 38858 47827 38861
rect 49200 38858 50000 38948
rect 47761 38856 50000 38858
rect 47761 38800 47766 38856
rect 47822 38800 50000 38856
rect 47761 38798 50000 38800
rect 47761 38795 47827 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 20529 38450 20595 38453
rect 20486 38448 20595 38450
rect 20486 38392 20534 38448
rect 20590 38392 20595 38448
rect 20486 38387 20595 38392
rect 0 38028 800 38268
rect 19333 38180 19399 38181
rect 19333 38176 19380 38180
rect 19444 38178 19450 38180
rect 19333 38120 19338 38176
rect 19333 38116 19380 38120
rect 19444 38118 19490 38178
rect 19444 38116 19450 38118
rect 19333 38115 19399 38116
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 20486 37909 20546 38387
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 49200 38028 50000 38118
rect 17309 37906 17375 37909
rect 18689 37906 18755 37909
rect 17309 37904 18755 37906
rect 17309 37848 17314 37904
rect 17370 37848 18694 37904
rect 18750 37848 18755 37904
rect 17309 37846 18755 37848
rect 17309 37843 17375 37846
rect 18689 37843 18755 37846
rect 19241 37906 19307 37909
rect 20161 37906 20227 37909
rect 19241 37904 20227 37906
rect 19241 37848 19246 37904
rect 19302 37848 20166 37904
rect 20222 37848 20227 37904
rect 19241 37846 20227 37848
rect 20486 37904 20595 37909
rect 20486 37848 20534 37904
rect 20590 37848 20595 37904
rect 20486 37846 20595 37848
rect 19241 37843 19307 37846
rect 20161 37843 20227 37846
rect 20529 37843 20595 37846
rect 14365 37770 14431 37773
rect 19333 37770 19399 37773
rect 23105 37770 23171 37773
rect 14365 37768 17970 37770
rect 14365 37712 14370 37768
rect 14426 37712 17970 37768
rect 14365 37710 17970 37712
rect 14365 37707 14431 37710
rect 17910 37634 17970 37710
rect 19333 37768 23171 37770
rect 19333 37712 19338 37768
rect 19394 37712 23110 37768
rect 23166 37712 23171 37768
rect 19333 37710 23171 37712
rect 19333 37707 19399 37710
rect 23105 37707 23171 37710
rect 27429 37634 27495 37637
rect 17910 37632 27495 37634
rect 0 37348 800 37588
rect 17910 37576 27434 37632
rect 27490 37576 27495 37632
rect 17910 37574 27495 37576
rect 27429 37571 27495 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 23565 35730 23631 35733
rect 26233 35730 26299 35733
rect 23565 35728 26299 35730
rect 23565 35672 23570 35728
rect 23626 35672 26238 35728
rect 26294 35672 26299 35728
rect 23565 35670 26299 35672
rect 23565 35667 23631 35670
rect 26233 35667 26299 35670
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 20713 35050 20779 35053
rect 27521 35050 27587 35053
rect 20713 35048 27587 35050
rect 20713 34992 20718 35048
rect 20774 34992 27526 35048
rect 27582 34992 27587 35048
rect 20713 34990 27587 34992
rect 20713 34987 20779 34990
rect 27521 34987 27587 34990
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48129 34098 48195 34101
rect 49200 34098 50000 34188
rect 48129 34096 50000 34098
rect 48129 34040 48134 34096
rect 48190 34040 50000 34096
rect 48129 34038 50000 34040
rect 48129 34035 48195 34038
rect 49200 33948 50000 34038
rect 19333 33828 19399 33829
rect 19333 33824 19380 33828
rect 19444 33826 19450 33828
rect 19333 33768 19338 33824
rect 19333 33764 19380 33768
rect 19444 33766 19490 33826
rect 19444 33764 19450 33766
rect 19333 33763 19399 33764
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 47945 33418 48011 33421
rect 49200 33418 50000 33508
rect 47945 33416 50000 33418
rect 47945 33360 47950 33416
rect 48006 33360 50000 33416
rect 47945 33358 50000 33360
rect 47945 33355 48011 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 47945 32058 48011 32061
rect 49200 32058 50000 32148
rect 47945 32056 50000 32058
rect 47945 32000 47950 32056
rect 48006 32000 50000 32056
rect 47945 31998 50000 32000
rect 47945 31995 48011 31998
rect 49200 31908 50000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3325 31378 3391 31381
rect 0 31376 3391 31378
rect 0 31320 3330 31376
rect 3386 31320 3391 31376
rect 0 31318 3391 31320
rect 0 31228 800 31318
rect 3325 31315 3391 31318
rect 46105 31378 46171 31381
rect 49200 31378 50000 31468
rect 46105 31376 50000 31378
rect 46105 31320 46110 31376
rect 46166 31320 50000 31376
rect 46105 31318 50000 31320
rect 46105 31315 46171 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 20805 30562 20871 30565
rect 26877 30562 26943 30565
rect 20805 30560 26943 30562
rect 20805 30504 20810 30560
rect 20866 30504 26882 30560
rect 26938 30504 26943 30560
rect 49200 30548 50000 30788
rect 20805 30502 26943 30504
rect 20805 30499 20871 30502
rect 26877 30499 26943 30502
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 20529 30290 20595 30293
rect 25957 30290 26023 30293
rect 20529 30288 26023 30290
rect 20529 30232 20534 30288
rect 20590 30232 25962 30288
rect 26018 30232 26023 30288
rect 20529 30230 26023 30232
rect 20529 30227 20595 30230
rect 25957 30227 26023 30230
rect 0 29868 800 30108
rect 45829 30018 45895 30021
rect 49200 30018 50000 30108
rect 45829 30016 50000 30018
rect 45829 29960 45834 30016
rect 45890 29960 50000 30016
rect 45829 29958 50000 29960
rect 45829 29955 45895 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19977 29474 20043 29477
rect 24945 29474 25011 29477
rect 19977 29472 25011 29474
rect 19977 29416 19982 29472
rect 20038 29416 24950 29472
rect 25006 29416 25011 29472
rect 19977 29414 25011 29416
rect 19977 29411 20043 29414
rect 24945 29411 25011 29414
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 48129 29338 48195 29341
rect 49200 29338 50000 29428
rect 48129 29336 50000 29338
rect 48129 29280 48134 29336
rect 48190 29280 50000 29336
rect 48129 29278 50000 29280
rect 48129 29275 48195 29278
rect 14457 29202 14523 29205
rect 18137 29202 18203 29205
rect 14457 29200 18203 29202
rect 14457 29144 14462 29200
rect 14518 29144 18142 29200
rect 18198 29144 18203 29200
rect 49200 29188 50000 29278
rect 14457 29142 18203 29144
rect 14457 29139 14523 29142
rect 18137 29139 18203 29142
rect 25773 29066 25839 29069
rect 26969 29066 27035 29069
rect 25773 29064 27035 29066
rect 25773 29008 25778 29064
rect 25834 29008 26974 29064
rect 27030 29008 27035 29064
rect 25773 29006 27035 29008
rect 25773 29003 25839 29006
rect 26969 29003 27035 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3325 28658 3391 28661
rect 0 28656 3391 28658
rect 0 28600 3330 28656
rect 3386 28600 3391 28656
rect 0 28598 3391 28600
rect 0 28508 800 28598
rect 3325 28595 3391 28598
rect 45553 28658 45619 28661
rect 49200 28658 50000 28748
rect 45553 28656 50000 28658
rect 45553 28600 45558 28656
rect 45614 28600 50000 28656
rect 45553 28598 50000 28600
rect 45553 28595 45619 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 21081 27842 21147 27845
rect 23749 27842 23815 27845
rect 21081 27840 23815 27842
rect 21081 27784 21086 27840
rect 21142 27784 23754 27840
rect 23810 27784 23815 27840
rect 49200 27828 50000 27918
rect 21081 27782 23815 27784
rect 21081 27779 21147 27782
rect 23749 27779 23815 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 45461 26618 45527 26621
rect 49200 26618 50000 26708
rect 45461 26616 50000 26618
rect 45461 26560 45466 26616
rect 45522 26560 50000 26616
rect 45461 26558 50000 26560
rect 45461 26555 45527 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 46841 25938 46907 25941
rect 49200 25938 50000 26028
rect 46841 25936 50000 25938
rect 46841 25880 46846 25936
rect 46902 25880 50000 25936
rect 46841 25878 50000 25880
rect 46841 25875 46907 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 48221 25258 48287 25261
rect 49200 25258 50000 25348
rect 48221 25256 50000 25258
rect 48221 25200 48226 25256
rect 48282 25200 50000 25256
rect 48221 25198 50000 25200
rect 48221 25195 48287 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 45553 23898 45619 23901
rect 49200 23898 50000 23988
rect 45553 23896 50000 23898
rect 45553 23840 45558 23896
rect 45614 23840 50000 23896
rect 45553 23838 50000 23840
rect 45553 23835 45619 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 46749 23218 46815 23221
rect 49200 23218 50000 23308
rect 46749 23216 50000 23218
rect 46749 23160 46754 23216
rect 46810 23160 50000 23216
rect 46749 23158 50000 23160
rect 46749 23155 46815 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46197 22538 46263 22541
rect 49200 22538 50000 22628
rect 46197 22536 50000 22538
rect 46197 22480 46202 22536
rect 46258 22480 50000 22536
rect 46197 22478 50000 22480
rect 46197 22475 46263 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 47945 21858 48011 21861
rect 49200 21858 50000 21948
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 23289 20770 23355 20773
rect 23565 20770 23631 20773
rect 23289 20768 23631 20770
rect 23289 20712 23294 20768
rect 23350 20712 23570 20768
rect 23626 20712 23631 20768
rect 23289 20710 23631 20712
rect 23289 20707 23355 20710
rect 23565 20707 23631 20710
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 19885 20498 19951 20501
rect 23197 20498 23263 20501
rect 19885 20496 23263 20498
rect 19885 20440 19890 20496
rect 19946 20440 23202 20496
rect 23258 20440 23263 20496
rect 19885 20438 23263 20440
rect 19885 20435 19951 20438
rect 23197 20435 23263 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3049 19818 3115 19821
rect 0 19816 3115 19818
rect 0 19760 3054 19816
rect 3110 19760 3115 19816
rect 0 19758 3115 19760
rect 0 19668 800 19758
rect 3049 19755 3115 19758
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3417 18458 3483 18461
rect 0 18456 3483 18458
rect 0 18400 3422 18456
rect 3478 18400 3483 18456
rect 0 18398 3483 18400
rect 0 18308 800 18398
rect 3417 18395 3483 18398
rect 45645 18458 45711 18461
rect 49200 18458 50000 18548
rect 45645 18456 50000 18458
rect 45645 18400 45650 18456
rect 45706 18400 50000 18456
rect 45645 18398 50000 18400
rect 45645 18395 45711 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1853 17778 1919 17781
rect 0 17776 1919 17778
rect 0 17720 1858 17776
rect 1914 17720 1919 17776
rect 0 17718 1919 17720
rect 0 17628 800 17718
rect 1853 17715 1919 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3049 17098 3115 17101
rect 0 17096 3115 17098
rect 0 17040 3054 17096
rect 3110 17040 3115 17096
rect 0 17038 3115 17040
rect 0 16948 800 17038
rect 3049 17035 3115 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45645 15738 45711 15741
rect 49200 15738 50000 15828
rect 45645 15736 50000 15738
rect 45645 15680 45650 15736
rect 45706 15680 50000 15736
rect 45645 15678 50000 15680
rect 45645 15675 45711 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13548 800 13638
rect 3417 13635 3483 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 4061 10298 4127 10301
rect 0 10296 4127 10298
rect 0 10240 4066 10296
rect 4122 10240 4127 10296
rect 0 10238 4127 10240
rect 0 10148 800 10238
rect 4061 10235 4127 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 47853 9618 47919 9621
rect 49200 9618 50000 9708
rect 47853 9616 50000 9618
rect 47853 9560 47858 9616
rect 47914 9560 50000 9616
rect 47853 9558 50000 9560
rect 47853 9555 47919 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 46013 8258 46079 8261
rect 49200 8258 50000 8348
rect 46013 8256 50000 8258
rect 46013 8200 46018 8256
rect 46074 8200 50000 8256
rect 46013 8198 50000 8200
rect 46013 8195 46079 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3233 7578 3299 7581
rect 0 7576 3299 7578
rect 0 7520 3238 7576
rect 3294 7520 3299 7576
rect 0 7518 3299 7520
rect 0 7428 800 7518
rect 3233 7515 3299 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6748 800 6838
rect 4061 6835 4127 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 47945 6218 48011 6221
rect 49200 6218 50000 6308
rect 47945 6216 50000 6218
rect 47945 6160 47950 6216
rect 48006 6160 50000 6216
rect 47945 6158 50000 6160
rect 47945 6155 48011 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 49200 4028 50000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 22737 3634 22803 3637
rect 25221 3634 25287 3637
rect 22737 3632 25287 3634
rect 0 3498 800 3588
rect 22737 3576 22742 3632
rect 22798 3576 25226 3632
rect 25282 3576 25287 3632
rect 22737 3574 25287 3576
rect 22737 3571 22803 3574
rect 25221 3571 25287 3574
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3348 800 3438
rect 4061 3435 4127 3438
rect 47761 3498 47827 3501
rect 49200 3498 50000 3588
rect 47761 3496 50000 3498
rect 47761 3440 47766 3496
rect 47822 3440 50000 3496
rect 47761 3438 50000 3440
rect 47761 3435 47827 3438
rect 22553 3362 22619 3365
rect 27429 3362 27495 3365
rect 22553 3360 27495 3362
rect 22553 3304 22558 3360
rect 22614 3304 27434 3360
rect 27490 3304 27495 3360
rect 49200 3348 50000 3438
rect 22553 3302 27495 3304
rect 22553 3299 22619 3302
rect 27429 3299 27495 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 19701 3090 19767 3093
rect 21817 3090 21883 3093
rect 19701 3088 21883 3090
rect 19701 3032 19706 3088
rect 19762 3032 21822 3088
rect 21878 3032 21883 3088
rect 19701 3030 21883 3032
rect 19701 3027 19767 3030
rect 21817 3027 21883 3030
rect 22185 2954 22251 2957
rect 26141 2954 26207 2957
rect 22185 2952 26207 2954
rect 0 2668 800 2908
rect 22185 2896 22190 2952
rect 22246 2896 26146 2952
rect 26202 2896 26207 2952
rect 22185 2894 26207 2896
rect 22185 2891 22251 2894
rect 26141 2891 26207 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1308 800 1398
rect 3509 1395 3575 1398
rect 46749 1458 46815 1461
rect 49200 1458 50000 1548
rect 46749 1456 50000 1458
rect 46749 1400 46754 1456
rect 46810 1400 50000 1456
rect 46749 1398 50000 1400
rect 46749 1395 46815 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 48037 778 48103 781
rect 49200 778 50000 868
rect 48037 776 50000 778
rect 48037 720 48042 776
rect 48098 720 50000 776
rect 48037 718 50000 720
rect 48037 715 48103 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19380 38176 19444 38180
rect 19380 38120 19394 38176
rect 19394 38120 19444 38176
rect 19380 38116 19444 38120
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19380 33824 19444 33828
rect 19380 33768 19394 33824
rect 19394 33768 19444 33824
rect 19380 33764 19444 33768
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19379 38180 19445 38181
rect 19379 38116 19380 38180
rect 19444 38116 19445 38180
rect 19379 38115 19445 38116
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 19382 33829 19442 38115
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19379 33828 19445 33829
rect 19379 33764 19380 33828
rect 19444 33764 19445 33828
rect 19379 33763 19445 33764
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33488 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 45908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 22540 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform -1 0 35696 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 40296 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 36432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 23920 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform 1 0 22172 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1644511149
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_200
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_207 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_242
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1644511149
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1644511149
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_314
timestamp 1644511149
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_412
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1644511149
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_88
timestamp 1644511149
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_96
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_172
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_180
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1644511149
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_257
timestamp 1644511149
transform 1 0 24748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_265
timestamp 1644511149
transform 1 0 25484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_289
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_301
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_313
timestamp 1644511149
transform 1 0 29900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_325
timestamp 1644511149
transform 1 0 31004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1644511149
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_359
timestamp 1644511149
transform 1 0 34132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_371
timestamp 1644511149
transform 1 0 35236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_423
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_434
timestamp 1644511149
transform 1 0 41032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_116
timestamp 1644511149
transform 1 0 11776 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_148
timestamp 1644511149
transform 1 0 14720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_156
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1644511149
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1644511149
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_228
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_239
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_261
timestamp 1644511149
transform 1 0 25116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_278
timestamp 1644511149
transform 1 0 26680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1644511149
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_329
timestamp 1644511149
transform 1 0 31372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_337
timestamp 1644511149
transform 1 0 32108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_341
timestamp 1644511149
transform 1 0 32476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_353
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1644511149
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_405
timestamp 1644511149
transform 1 0 38364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_409
timestamp 1644511149
transform 1 0 38732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1644511149
transform 1 0 40572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_441
timestamp 1644511149
transform 1 0 41676 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_449
timestamp 1644511149
transform 1 0 42412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1644511149
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_96
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_122
timestamp 1644511149
transform 1 0 12328 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp 1644511149
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 1644511149
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_190
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_198
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_209
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1644511149
transform 1 0 24840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_262
timestamp 1644511149
transform 1 0 25208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_408
timestamp 1644511149
transform 1 0 38640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_419
timestamp 1644511149
transform 1 0 39652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1644511149
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_458
timestamp 1644511149
transform 1 0 43240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_465
timestamp 1644511149
transform 1 0 43884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_477
timestamp 1644511149
transform 1 0 44988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_499
timestamp 1644511149
transform 1 0 47012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1644511149
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1644511149
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_383
timestamp 1644511149
transform 1 0 36340 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_386
timestamp 1644511149
transform 1 0 36616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_425
timestamp 1644511149
transform 1 0 40204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_432
timestamp 1644511149
transform 1 0 40848 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_444
timestamp 1644511149
transform 1 0 41952 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_456
timestamp 1644511149
transform 1 0 43056 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_468
timestamp 1644511149
transform 1 0 44160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_235
timestamp 1644511149
transform 1 0 22724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_247
timestamp 1644511149
transform 1 0 23828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_259
timestamp 1644511149
transform 1 0 24932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1644511149
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_431
timestamp 1644511149
transform 1 0 40756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1644511149
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_441
timestamp 1644511149
transform 1 0 41676 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_455
timestamp 1644511149
transform 1 0 42964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_467
timestamp 1644511149
transform 1 0 44068 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_433
timestamp 1644511149
transform 1 0 40940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_445
timestamp 1644511149
transform 1 0 42044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_425
timestamp 1644511149
transform 1 0 40204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_428
timestamp 1644511149
transform 1 0 40480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_443
timestamp 1644511149
transform 1 0 41860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_455
timestamp 1644511149
transform 1 0 42964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_467
timestamp 1644511149
transform 1 0 44068 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_489
timestamp 1644511149
transform 1 0 46092 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1644511149
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_481
timestamp 1644511149
transform 1 0 45356 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_495
timestamp 1644511149
transform 1 0 46644 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_505
timestamp 1644511149
transform 1 0 47564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1644511149
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_493
timestamp 1644511149
transform 1 0 46460 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_498
timestamp 1644511149
transform 1 0 46920 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1644511149
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_234
timestamp 1644511149
transform 1 0 22632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_246
timestamp 1644511149
transform 1 0 23736 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_258
timestamp 1644511149
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1644511149
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1644511149
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_507
timestamp 1644511149
transform 1 0 47748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_515
timestamp 1644511149
transform 1 0 48484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1644511149
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_244
timestamp 1644511149
transform 1 0 23552 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_258
timestamp 1644511149
transform 1 0 24840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_270
timestamp 1644511149
transform 1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1644511149
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_227
timestamp 1644511149
transform 1 0 21988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_235
timestamp 1644511149
transform 1 0 22724 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_256
timestamp 1644511149
transform 1 0 24656 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_262
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_284
timestamp 1644511149
transform 1 0 27232 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_296
timestamp 1644511149
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_317
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1644511149
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1644511149
transform 1 0 33396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_507
timestamp 1644511149
transform 1 0 47748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1644511149
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_200
timestamp 1644511149
transform 1 0 19504 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_212
timestamp 1644511149
transform 1 0 20608 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_229
timestamp 1644511149
transform 1 0 22172 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_256
timestamp 1644511149
transform 1 0 24656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_285
timestamp 1644511149
transform 1 0 27324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_299
timestamp 1644511149
transform 1 0 28612 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_311
timestamp 1644511149
transform 1 0 29716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_323
timestamp 1644511149
transform 1 0 30820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_456
timestamp 1644511149
transform 1 0 43056 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_464
timestamp 1644511149
transform 1 0 43792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_486
timestamp 1644511149
transform 1 0 45816 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_498
timestamp 1644511149
transform 1 0 46920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 1644511149
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_179
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_187
timestamp 1644511149
transform 1 0 18308 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_204
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_273
timestamp 1644511149
transform 1 0 26220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_280
timestamp 1644511149
transform 1 0 26864 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_288
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_293
timestamp 1644511149
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1644511149
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_330
timestamp 1644511149
transform 1 0 31464 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_342
timestamp 1644511149
transform 1 0 32568 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_354
timestamp 1644511149
transform 1 0 33672 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1644511149
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_472
timestamp 1644511149
transform 1 0 44528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_480
timestamp 1644511149
transform 1 0 45264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_488
timestamp 1644511149
transform 1 0 46000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_119
timestamp 1644511149
transform 1 0 12052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_131
timestamp 1644511149
transform 1 0 13156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_142
timestamp 1644511149
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_154
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1644511149
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_177
timestamp 1644511149
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_214
timestamp 1644511149
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1644511149
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1644511149
transform 1 0 23644 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_253
timestamp 1644511149
transform 1 0 24380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_266
timestamp 1644511149
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_285
timestamp 1644511149
transform 1 0 27324 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_296
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1644511149
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1644511149
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_488
timestamp 1644511149
transform 1 0 46000 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_499
timestamp 1644511149
transform 1 0 47012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_146
timestamp 1644511149
transform 1 0 14536 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_158
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_180
timestamp 1644511149
transform 1 0 17664 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_188
timestamp 1644511149
transform 1 0 18400 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_204
timestamp 1644511149
transform 1 0 19872 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_210
timestamp 1644511149
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_214
timestamp 1644511149
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_226
timestamp 1644511149
transform 1 0 21896 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_238
timestamp 1644511149
transform 1 0 23000 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1644511149
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_281
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_287
timestamp 1644511149
transform 1 0 27508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_298
timestamp 1644511149
transform 1 0 28520 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1644511149
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_318
timestamp 1644511149
transform 1 0 30360 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_324
timestamp 1644511149
transform 1 0 30912 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_346
timestamp 1644511149
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1644511149
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_437
timestamp 1644511149
transform 1 0 41308 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_459
timestamp 1644511149
transform 1 0 43332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_470
timestamp 1644511149
transform 1 0 44344 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_485
timestamp 1644511149
transform 1 0 45724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1644511149
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_119
timestamp 1644511149
transform 1 0 12052 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1644511149
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1644511149
transform 1 0 16928 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_200
timestamp 1644511149
transform 1 0 19504 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_212
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_233
timestamp 1644511149
transform 1 0 22540 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_238
timestamp 1644511149
transform 1 0 23000 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_263
timestamp 1644511149
transform 1 0 25300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_275
timestamp 1644511149
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp 1644511149
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1644511149
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_303
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_343
timestamp 1644511149
transform 1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_350
timestamp 1644511149
transform 1 0 33304 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_362
timestamp 1644511149
transform 1 0 34408 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_374
timestamp 1644511149
transform 1 0 35512 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1644511149
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_444
timestamp 1644511149
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_475
timestamp 1644511149
transform 1 0 44804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_510
timestamp 1644511149
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_173
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_185
timestamp 1644511149
transform 1 0 18124 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1644511149
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_217
timestamp 1644511149
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_223
timestamp 1644511149
transform 1 0 21620 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1644511149
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_260
timestamp 1644511149
transform 1 0 25024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_284
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_296
timestamp 1644511149
transform 1 0 28336 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1644511149
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_316
timestamp 1644511149
transform 1 0 30176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_320
timestamp 1644511149
transform 1 0 30544 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_342
timestamp 1644511149
transform 1 0 32568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_352
timestamp 1644511149
transform 1 0 33488 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1644511149
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_482
timestamp 1644511149
transform 1 0 45448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_498
timestamp 1644511149
transform 1 0 46920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_505
timestamp 1644511149
transform 1 0 47564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_151
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1644511149
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1644511149
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_196
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_203
timestamp 1644511149
transform 1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1644511149
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_248
timestamp 1644511149
transform 1 0 23920 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_272
timestamp 1644511149
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_284
timestamp 1644511149
transform 1 0 27232 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_292
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_295
timestamp 1644511149
transform 1 0 28244 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_302
timestamp 1644511149
transform 1 0 28888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_311
timestamp 1644511149
transform 1 0 29716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_323
timestamp 1644511149
transform 1 0 30820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_350
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_354
timestamp 1644511149
transform 1 0 33672 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_366
timestamp 1644511149
transform 1 0 34776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_378
timestamp 1644511149
transform 1 0 35880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1644511149
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_455
timestamp 1644511149
transform 1 0 42964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_459
timestamp 1644511149
transform 1 0 43332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_471
timestamp 1644511149
transform 1 0 44436 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_479
timestamp 1644511149
transform 1 0 45172 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_496
timestamp 1644511149
transform 1 0 46736 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1644511149
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1644511149
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1644511149
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1644511149
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1644511149
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1644511149
transform 1 0 20884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_223
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1644511149
transform 1 0 21988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_239
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_243
timestamp 1644511149
transform 1 0 23460 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_257
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_275
timestamp 1644511149
transform 1 0 26404 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_287
timestamp 1644511149
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_312
timestamp 1644511149
transform 1 0 29808 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_318
timestamp 1644511149
transform 1 0 30360 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_340
timestamp 1644511149
transform 1 0 32384 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_346
timestamp 1644511149
transform 1 0 32936 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1644511149
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_453
timestamp 1644511149
transform 1 0 42780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_459
timestamp 1644511149
transform 1 0 43332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_463
timestamp 1644511149
transform 1 0 43700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_467
timestamp 1644511149
transform 1 0 44068 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_480
timestamp 1644511149
transform 1 0 45264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_487
timestamp 1644511149
transform 1 0 45908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_121
timestamp 1644511149
transform 1 0 12236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_145
timestamp 1644511149
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_155
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_173
timestamp 1644511149
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_185
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_210
timestamp 1644511149
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1644511149
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_229
timestamp 1644511149
transform 1 0 22172 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_241
timestamp 1644511149
transform 1 0 23276 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_247
timestamp 1644511149
transform 1 0 23828 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_253
timestamp 1644511149
transform 1 0 24380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1644511149
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1644511149
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_285
timestamp 1644511149
transform 1 0 27324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_297
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_303
timestamp 1644511149
transform 1 0 28980 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_307
timestamp 1644511149
transform 1 0 29348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_322
timestamp 1644511149
transform 1 0 30728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1644511149
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_352
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_364
timestamp 1644511149
transform 1 0 34592 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_376
timestamp 1644511149
transform 1 0 35696 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_452
timestamp 1644511149
transform 1 0 42688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_463
timestamp 1644511149
transform 1 0 43700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_512
timestamp 1644511149
transform 1 0 48208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_160
timestamp 1644511149
transform 1 0 15824 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_180
timestamp 1644511149
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_218
timestamp 1644511149
transform 1 0 21160 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1644511149
transform 1 0 21988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_239
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1644511149
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_260
timestamp 1644511149
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_294
timestamp 1644511149
transform 1 0 28152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_330
timestamp 1644511149
transform 1 0 31464 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_342
timestamp 1644511149
transform 1 0 32568 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1644511149
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_386
timestamp 1644511149
transform 1 0 36616 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_398
timestamp 1644511149
transform 1 0 37720 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_410
timestamp 1644511149
transform 1 0 38824 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1644511149
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_451
timestamp 1644511149
transform 1 0 42596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_468
timestamp 1644511149
transform 1 0 44160 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_482
timestamp 1644511149
transform 1 0 45448 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_490
timestamp 1644511149
transform 1 0 46184 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_134
timestamp 1644511149
transform 1 0 13432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_142
timestamp 1644511149
transform 1 0 14168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_190
timestamp 1644511149
transform 1 0 18584 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_198
timestamp 1644511149
transform 1 0 19320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_235
timestamp 1644511149
transform 1 0 22724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_243
timestamp 1644511149
transform 1 0 23460 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_263
timestamp 1644511149
transform 1 0 25300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_274
timestamp 1644511149
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_289
timestamp 1644511149
transform 1 0 27692 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_316
timestamp 1644511149
transform 1 0 30176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_320
timestamp 1644511149
transform 1 0 30544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_340
timestamp 1644511149
transform 1 0 32384 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_360
timestamp 1644511149
transform 1 0 34224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_365
timestamp 1644511149
transform 1 0 34684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_382
timestamp 1644511149
transform 1 0 36248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1644511149
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_458
timestamp 1644511149
transform 1 0 43240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_462
timestamp 1644511149
transform 1 0 43608 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_466
timestamp 1644511149
transform 1 0 43976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_483
timestamp 1644511149
transform 1 0 45540 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_489
timestamp 1644511149
transform 1 0 46092 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_510
timestamp 1644511149
transform 1 0 48024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_113
timestamp 1644511149
transform 1 0 11500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1644511149
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1644511149
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_200
timestamp 1644511149
transform 1 0 19504 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_217
timestamp 1644511149
transform 1 0 21068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_229
timestamp 1644511149
transform 1 0 22172 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_263
timestamp 1644511149
transform 1 0 25300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_273
timestamp 1644511149
transform 1 0 26220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1644511149
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_313
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_324
timestamp 1644511149
transform 1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_348
timestamp 1644511149
transform 1 0 33120 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_372
timestamp 1644511149
transform 1 0 35328 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_376
timestamp 1644511149
transform 1 0 35696 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_388
timestamp 1644511149
transform 1 0 36800 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_400
timestamp 1644511149
transform 1 0 37904 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_412
timestamp 1644511149
transform 1 0 39008 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_430
timestamp 1644511149
transform 1 0 40664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_442
timestamp 1644511149
transform 1 0 41768 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_454
timestamp 1644511149
transform 1 0 42872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_458
timestamp 1644511149
transform 1 0 43240 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_462
timestamp 1644511149
transform 1 0 43608 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_471
timestamp 1644511149
transform 1 0 44436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_500
timestamp 1644511149
transform 1 0 47104 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_511
timestamp 1644511149
transform 1 0 48116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_515
timestamp 1644511149
transform 1 0 48484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_120
timestamp 1644511149
transform 1 0 12144 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_128
timestamp 1644511149
transform 1 0 12880 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_132
timestamp 1644511149
transform 1 0 13248 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_144
timestamp 1644511149
transform 1 0 14352 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_233
timestamp 1644511149
transform 1 0 22540 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_238
timestamp 1644511149
transform 1 0 23000 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_250
timestamp 1644511149
transform 1 0 24104 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_262
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_267
timestamp 1644511149
transform 1 0 25668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_289
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_295
timestamp 1644511149
transform 1 0 28244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_299
timestamp 1644511149
transform 1 0 28612 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_321
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_325
timestamp 1644511149
transform 1 0 31004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1644511149
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_340
timestamp 1644511149
transform 1 0 32384 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_352
timestamp 1644511149
transform 1 0 33488 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_364
timestamp 1644511149
transform 1 0 34592 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_376
timestamp 1644511149
transform 1 0 35696 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_431
timestamp 1644511149
transform 1 0 40756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_443
timestamp 1644511149
transform 1 0 41860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_454
timestamp 1644511149
transform 1 0 42872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_469
timestamp 1644511149
transform 1 0 44252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_475
timestamp 1644511149
transform 1 0 44804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_160
timestamp 1644511149
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1644511149
transform 1 0 17480 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1644511149
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_204
timestamp 1644511149
transform 1 0 19872 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_214
timestamp 1644511149
transform 1 0 20792 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_220
timestamp 1644511149
transform 1 0 21344 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_241
timestamp 1644511149
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1644511149
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_257
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_270
timestamp 1644511149
transform 1 0 25944 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_279
timestamp 1644511149
transform 1 0 26772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_286
timestamp 1644511149
transform 1 0 27416 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_294
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1644511149
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_319
timestamp 1644511149
transform 1 0 30452 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_353
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1644511149
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_369
timestamp 1644511149
transform 1 0 35052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_381
timestamp 1644511149
transform 1 0 36156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_393
timestamp 1644511149
transform 1 0 37260 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_405
timestamp 1644511149
transform 1 0 38364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_417
timestamp 1644511149
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_424
timestamp 1644511149
transform 1 0 40112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_449
timestamp 1644511149
transform 1 0 42412 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_458
timestamp 1644511149
transform 1 0 43240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_465
timestamp 1644511149
transform 1 0 43884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_473
timestamp 1644511149
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_483
timestamp 1644511149
transform 1 0 45540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_487
timestamp 1644511149
transform 1 0 45908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_120
timestamp 1644511149
transform 1 0 12144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_132
timestamp 1644511149
transform 1 0 13248 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_144
timestamp 1644511149
transform 1 0 14352 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_157
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_189
timestamp 1644511149
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_200
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_206
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1644511149
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1644511149
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_229
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_238
timestamp 1644511149
transform 1 0 23000 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_244
timestamp 1644511149
transform 1 0 23552 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_268
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_301
timestamp 1644511149
transform 1 0 28796 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_309
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_314
timestamp 1644511149
transform 1 0 29992 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_324
timestamp 1644511149
transform 1 0 30912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1644511149
transform 1 0 32476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_357
timestamp 1644511149
transform 1 0 33948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_381
timestamp 1644511149
transform 1 0 36156 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1644511149
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_396
timestamp 1644511149
transform 1 0 37536 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_408
timestamp 1644511149
transform 1 0 38640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_431
timestamp 1644511149
transform 1 0 40756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_442
timestamp 1644511149
transform 1 0 41768 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_455
timestamp 1644511149
transform 1 0 42964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_478
timestamp 1644511149
transform 1 0 45080 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_486
timestamp 1644511149
transform 1 0 45816 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_490
timestamp 1644511149
transform 1 0 46184 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_126
timestamp 1644511149
transform 1 0 12696 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_149
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_163
timestamp 1644511149
transform 1 0 16100 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_171
timestamp 1644511149
transform 1 0 16836 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_214
timestamp 1644511149
transform 1 0 20792 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_218
timestamp 1644511149
transform 1 0 21160 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1644511149
transform 1 0 23092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_258
timestamp 1644511149
transform 1 0 24840 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_273
timestamp 1644511149
transform 1 0 26220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_300
timestamp 1644511149
transform 1 0 28704 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_313
timestamp 1644511149
transform 1 0 29900 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_317
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_330
timestamp 1644511149
transform 1 0 31464 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_343
timestamp 1644511149
transform 1 0 32660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_352
timestamp 1644511149
transform 1 0 33488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_356
timestamp 1644511149
transform 1 0 33856 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_369
timestamp 1644511149
transform 1 0 35052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_373
timestamp 1644511149
transform 1 0 35420 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_380
timestamp 1644511149
transform 1 0 36064 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_388
timestamp 1644511149
transform 1 0 36800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_411
timestamp 1644511149
transform 1 0 38916 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_428
timestamp 1644511149
transform 1 0 40480 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_440
timestamp 1644511149
transform 1 0 41584 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_452
timestamp 1644511149
transform 1 0 42688 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_458
timestamp 1644511149
transform 1 0 43240 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_470
timestamp 1644511149
transform 1 0 44344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1644511149
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1644511149
transform 1 0 13524 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_143
timestamp 1644511149
transform 1 0 14260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_152
timestamp 1644511149
transform 1 0 15088 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_159
timestamp 1644511149
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_174
timestamp 1644511149
transform 1 0 17112 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_178
timestamp 1644511149
transform 1 0 17480 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_182
timestamp 1644511149
transform 1 0 17848 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_194
timestamp 1644511149
transform 1 0 18952 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_204
timestamp 1644511149
transform 1 0 19872 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1644511149
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_229
timestamp 1644511149
transform 1 0 22172 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_243
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_268
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_289
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_300
timestamp 1644511149
transform 1 0 28704 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_308
timestamp 1644511149
transform 1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_314
timestamp 1644511149
transform 1 0 29992 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1644511149
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_340
timestamp 1644511149
transform 1 0 32384 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_352
timestamp 1644511149
transform 1 0 33488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_363
timestamp 1644511149
transform 1 0 34500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1644511149
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_412
timestamp 1644511149
transform 1 0 39008 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_419
timestamp 1644511149
transform 1 0 39652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1644511149
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_479
timestamp 1644511149
transform 1 0 45172 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_491
timestamp 1644511149
transform 1 0 46276 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1644511149
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1644511149
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_167
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_185
timestamp 1644511149
transform 1 0 18124 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_203
timestamp 1644511149
transform 1 0 19780 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_215
timestamp 1644511149
transform 1 0 20884 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_257
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1644511149
transform 1 0 26220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_283
timestamp 1644511149
transform 1 0 27140 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_291
timestamp 1644511149
transform 1 0 27876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 1644511149
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 1644511149
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_338
timestamp 1644511149
transform 1 0 32200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1644511149
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1644511149
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_442
timestamp 1644511149
transform 1 0 41768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_467
timestamp 1644511149
transform 1 0 44068 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_481
timestamp 1644511149
transform 1 0 45356 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_503
timestamp 1644511149
transform 1 0 47380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_510
timestamp 1644511149
transform 1 0 48024 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_119
timestamp 1644511149
transform 1 0 12052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1644511149
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_154
timestamp 1644511149
transform 1 0 15272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_158
timestamp 1644511149
transform 1 0 15640 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1644511149
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1644511149
transform 1 0 17572 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_189
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_201
timestamp 1644511149
transform 1 0 19596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1644511149
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1644511149
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_231
timestamp 1644511149
transform 1 0 22356 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_246
timestamp 1644511149
transform 1 0 23736 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_258
timestamp 1644511149
transform 1 0 24840 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_262
timestamp 1644511149
transform 1 0 25208 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_272
timestamp 1644511149
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_344
timestamp 1644511149
transform 1 0 32752 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_354
timestamp 1644511149
transform 1 0 33672 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_363
timestamp 1644511149
transform 1 0 34500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_370
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_377
timestamp 1644511149
transform 1 0 35788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1644511149
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_399
timestamp 1644511149
transform 1 0 37812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_411
timestamp 1644511149
transform 1 0 38916 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_423
timestamp 1644511149
transform 1 0 40020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_435
timestamp 1644511149
transform 1 0 41124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_442
timestamp 1644511149
transform 1 0 41768 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_512
timestamp 1644511149
transform 1 0 48208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1644511149
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_127
timestamp 1644511149
transform 1 0 12788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1644511149
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1644511149
transform 1 0 14352 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1644511149
transform 1 0 15088 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_156
timestamp 1644511149
transform 1 0 15456 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_181
timestamp 1644511149
transform 1 0 17756 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_187
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_201
timestamp 1644511149
transform 1 0 19596 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_208
timestamp 1644511149
transform 1 0 20240 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_220
timestamp 1644511149
transform 1 0 21344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1644511149
transform 1 0 24840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_295
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_312
timestamp 1644511149
transform 1 0 29808 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_327
timestamp 1644511149
transform 1 0 31188 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_335
timestamp 1644511149
transform 1 0 31924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_344
timestamp 1644511149
transform 1 0 32752 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_352
timestamp 1644511149
transform 1 0 33488 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_385
timestamp 1644511149
transform 1 0 36524 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_393
timestamp 1644511149
transform 1 0 37260 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1644511149
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_126
timestamp 1644511149
transform 1 0 12696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_138
timestamp 1644511149
transform 1 0 13800 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_150
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_190
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_230
timestamp 1644511149
transform 1 0 22264 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_245
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1644511149
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1644511149
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_287
timestamp 1644511149
transform 1 0 27508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_291
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_312
timestamp 1644511149
transform 1 0 29808 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_324
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_357
timestamp 1644511149
transform 1 0 33948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_365
timestamp 1644511149
transform 1 0 34684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_377
timestamp 1644511149
transform 1 0 35788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1644511149
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_149
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_171
timestamp 1644511149
transform 1 0 16836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_183
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_204
timestamp 1644511149
transform 1 0 19872 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_212
timestamp 1644511149
transform 1 0 20608 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_223
timestamp 1644511149
transform 1 0 21620 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_234
timestamp 1644511149
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1644511149
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_258
timestamp 1644511149
transform 1 0 24840 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_266
timestamp 1644511149
transform 1 0 25576 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_293
timestamp 1644511149
transform 1 0 28060 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_314
timestamp 1644511149
transform 1 0 29992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_326
timestamp 1644511149
transform 1 0 31096 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_338
timestamp 1644511149
transform 1 0 32200 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_349
timestamp 1644511149
transform 1 0 33212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_371
timestamp 1644511149
transform 1 0 35236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_383
timestamp 1644511149
transform 1 0 36340 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_395
timestamp 1644511149
transform 1 0 37444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_407
timestamp 1644511149
transform 1 0 38548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_203
timestamp 1644511149
transform 1 0 19780 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_212
timestamp 1644511149
transform 1 0 20608 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1644511149
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_230
timestamp 1644511149
transform 1 0 22264 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_238
timestamp 1644511149
transform 1 0 23000 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1644511149
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_256
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_271
timestamp 1644511149
transform 1 0 26036 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_289
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_302
timestamp 1644511149
transform 1 0 28888 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_321
timestamp 1644511149
transform 1 0 30636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_333
timestamp 1644511149
transform 1 0 31740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_355
timestamp 1644511149
transform 1 0 33764 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_376
timestamp 1644511149
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_149
timestamp 1644511149
transform 1 0 14812 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_154
timestamp 1644511149
transform 1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_161
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_180
timestamp 1644511149
transform 1 0 17664 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_207
timestamp 1644511149
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_219
timestamp 1644511149
transform 1 0 21252 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_231
timestamp 1644511149
transform 1 0 22356 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1644511149
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_261
timestamp 1644511149
transform 1 0 25116 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_267
timestamp 1644511149
transform 1 0 25668 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_272
timestamp 1644511149
transform 1 0 26128 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_280
timestamp 1644511149
transform 1 0 26864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_287
timestamp 1644511149
transform 1 0 27508 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_295
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_329
timestamp 1644511149
transform 1 0 31372 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_337
timestamp 1644511149
transform 1 0 32108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_343
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 1644511149
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_507
timestamp 1644511149
transform 1 0 47748 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_515
timestamp 1644511149
transform 1 0 48484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_175
timestamp 1644511149
transform 1 0 17204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1644511149
transform 1 0 18032 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_196
timestamp 1644511149
transform 1 0 19136 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_204
timestamp 1644511149
transform 1 0 19872 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_210
timestamp 1644511149
transform 1 0 20424 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1644511149
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_265
timestamp 1644511149
transform 1 0 25484 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_290
timestamp 1644511149
transform 1 0 27784 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_299
timestamp 1644511149
transform 1 0 28612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_313
timestamp 1644511149
transform 1 0 29900 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_323
timestamp 1644511149
transform 1 0 30820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_360
timestamp 1644511149
transform 1 0 34224 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_372
timestamp 1644511149
transform 1 0 35328 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1644511149
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_161
timestamp 1644511149
transform 1 0 15916 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1644511149
transform 1 0 16744 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_179
timestamp 1644511149
transform 1 0 17572 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_191
timestamp 1644511149
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_205
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_213
timestamp 1644511149
transform 1 0 20700 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_224
timestamp 1644511149
transform 1 0 21712 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_237
timestamp 1644511149
transform 1 0 22908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1644511149
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_257
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_297
timestamp 1644511149
transform 1 0 28428 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1644511149
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_315
timestamp 1644511149
transform 1 0 30084 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_325
timestamp 1644511149
transform 1 0 31004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_337
timestamp 1644511149
transform 1 0 32108 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_350
timestamp 1644511149
transform 1 0 33304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1644511149
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_145
timestamp 1644511149
transform 1 0 14444 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_189
timestamp 1644511149
transform 1 0 18492 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_197
timestamp 1644511149
transform 1 0 19228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_201
timestamp 1644511149
transform 1 0 19596 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_213
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_247
timestamp 1644511149
transform 1 0 23828 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1644511149
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_284
timestamp 1644511149
transform 1 0 27232 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_292
timestamp 1644511149
transform 1 0 27968 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_296
timestamp 1644511149
transform 1 0 28336 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_314
timestamp 1644511149
transform 1 0 29992 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_326
timestamp 1644511149
transform 1 0 31096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1644511149
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_345
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1644511149
transform 1 0 35972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_160
timestamp 1644511149
transform 1 0 15824 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_178
timestamp 1644511149
transform 1 0 17480 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_186
timestamp 1644511149
transform 1 0 18216 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1644511149
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_227
timestamp 1644511149
transform 1 0 21988 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_236
timestamp 1644511149
transform 1 0 22816 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_260
timestamp 1644511149
transform 1 0 25024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_285
timestamp 1644511149
transform 1 0 27324 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_293
timestamp 1644511149
transform 1 0 28060 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_299
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_316
timestamp 1644511149
transform 1 0 30176 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_322
timestamp 1644511149
transform 1 0 30728 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_343
timestamp 1644511149
transform 1 0 32660 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_355
timestamp 1644511149
transform 1 0 33764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_495
timestamp 1644511149
transform 1 0 46644 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_509
timestamp 1644511149
transform 1 0 47932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_515
timestamp 1644511149
transform 1 0 48484 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_18
timestamp 1644511149
transform 1 0 2760 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_40
timestamp 1644511149
transform 1 0 4784 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1644511149
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_158
timestamp 1644511149
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1644511149
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_176
timestamp 1644511149
transform 1 0 17296 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_186
timestamp 1644511149
transform 1 0 18216 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_198
timestamp 1644511149
transform 1 0 19320 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_209
timestamp 1644511149
transform 1 0 20332 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_218
timestamp 1644511149
transform 1 0 21160 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_251
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_259
timestamp 1644511149
transform 1 0 24932 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_267
timestamp 1644511149
transform 1 0 25668 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1644511149
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_291
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_297
timestamp 1644511149
transform 1 0 28428 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_303
timestamp 1644511149
transform 1 0 28980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_309
timestamp 1644511149
transform 1 0 29532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_314
timestamp 1644511149
transform 1 0 29992 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_322
timestamp 1644511149
transform 1 0 30728 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1644511149
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_340
timestamp 1644511149
transform 1 0 32384 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_352
timestamp 1644511149
transform 1 0 33488 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_364
timestamp 1644511149
transform 1 0 34592 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_376
timestamp 1644511149
transform 1 0 35696 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_148
timestamp 1644511149
transform 1 0 14720 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_156
timestamp 1644511149
transform 1 0 15456 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_161
timestamp 1644511149
transform 1 0 15916 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_176
timestamp 1644511149
transform 1 0 17296 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_183
timestamp 1644511149
transform 1 0 17940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_201
timestamp 1644511149
transform 1 0 19596 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_206
timestamp 1644511149
transform 1 0 20056 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_217
timestamp 1644511149
transform 1 0 21068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_229
timestamp 1644511149
transform 1 0 22172 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_237
timestamp 1644511149
transform 1 0 22908 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1644511149
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_263
timestamp 1644511149
transform 1 0 25300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_270
timestamp 1644511149
transform 1 0 25944 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_278
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_286
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_297
timestamp 1644511149
transform 1 0 28428 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_313
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_329
timestamp 1644511149
transform 1 0 31372 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_339
timestamp 1644511149
transform 1 0 32292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_347
timestamp 1644511149
transform 1 0 33028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1644511149
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_6
timestamp 1644511149
transform 1 0 1656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_174
timestamp 1644511149
transform 1 0 17112 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_198
timestamp 1644511149
transform 1 0 19320 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_210
timestamp 1644511149
transform 1 0 20424 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_262
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_301
timestamp 1644511149
transform 1 0 28796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_310
timestamp 1644511149
transform 1 0 29624 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_319
timestamp 1644511149
transform 1 0 30452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_331
timestamp 1644511149
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_357
timestamp 1644511149
transform 1 0 33948 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_369
timestamp 1644511149
transform 1 0 35052 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_381
timestamp 1644511149
transform 1 0 36156 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_389
timestamp 1644511149
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1644511149
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_14
timestamp 1644511149
transform 1 0 2392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1644511149
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_150
timestamp 1644511149
transform 1 0 14904 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1644511149
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_170
timestamp 1644511149
transform 1 0 16744 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_183
timestamp 1644511149
transform 1 0 17940 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_225
timestamp 1644511149
transform 1 0 21804 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_232
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_238
timestamp 1644511149
transform 1 0 23000 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1644511149
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_285
timestamp 1644511149
transform 1 0 27324 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_297
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1644511149
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_320
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_328
timestamp 1644511149
transform 1 0 31280 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_339
timestamp 1644511149
transform 1 0 32292 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_348
timestamp 1644511149
transform 1 0 33120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1644511149
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_495
timestamp 1644511149
transform 1 0 46644 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_133
timestamp 1644511149
transform 1 0 13340 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_140
timestamp 1644511149
transform 1 0 13984 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_150
timestamp 1644511149
transform 1 0 14904 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_178
timestamp 1644511149
transform 1 0 17480 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_188
timestamp 1644511149
transform 1 0 18400 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_200
timestamp 1644511149
transform 1 0 19504 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_212
timestamp 1644511149
transform 1 0 20608 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_257
timestamp 1644511149
transform 1 0 24748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_262
timestamp 1644511149
transform 1 0 25208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_285
timestamp 1644511149
transform 1 0 27324 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_290
timestamp 1644511149
transform 1 0 27784 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_303
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_316
timestamp 1644511149
transform 1 0 30176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_326
timestamp 1644511149
transform 1 0 31096 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1644511149
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_357
timestamp 1644511149
transform 1 0 33948 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_369
timestamp 1644511149
transform 1 0 35052 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_381
timestamp 1644511149
transform 1 0 36156 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_389
timestamp 1644511149
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_511
timestamp 1644511149
transform 1 0 48116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_515
timestamp 1644511149
transform 1 0 48484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_161
timestamp 1644511149
transform 1 0 15916 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_168
timestamp 1644511149
transform 1 0 16560 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_183
timestamp 1644511149
transform 1 0 17940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_214
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_228
timestamp 1644511149
transform 1 0 22080 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_236
timestamp 1644511149
transform 1 0 22816 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_241
timestamp 1644511149
transform 1 0 23276 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_257
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_285
timestamp 1644511149
transform 1 0 27324 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1644511149
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_315
timestamp 1644511149
transform 1 0 30084 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_328
timestamp 1644511149
transform 1 0 31280 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_340
timestamp 1644511149
transform 1 0 32384 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_352
timestamp 1644511149
transform 1 0 33488 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_507
timestamp 1644511149
transform 1 0 47748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_141
timestamp 1644511149
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_145
timestamp 1644511149
transform 1 0 14444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_156
timestamp 1644511149
transform 1 0 15456 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_184
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_216
timestamp 1644511149
transform 1 0 20976 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_230
timestamp 1644511149
transform 1 0 22264 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_238
timestamp 1644511149
transform 1 0 23000 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_243
timestamp 1644511149
transform 1 0 23460 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_254
timestamp 1644511149
transform 1 0 24472 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_266
timestamp 1644511149
transform 1 0 25576 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_318
timestamp 1644511149
transform 1 0 30360 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_328
timestamp 1644511149
transform 1 0 31280 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_340
timestamp 1644511149
transform 1 0 32384 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_352
timestamp 1644511149
transform 1 0 33488 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_364
timestamp 1644511149
transform 1 0 34592 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_376
timestamp 1644511149
transform 1 0 35696 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_169
timestamp 1644511149
transform 1 0 16652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_190
timestamp 1644511149
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_203
timestamp 1644511149
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_213
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_223
timestamp 1644511149
transform 1 0 21620 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_257
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_274
timestamp 1644511149
transform 1 0 26312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_282
timestamp 1644511149
transform 1 0 27048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_317
timestamp 1644511149
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_338
timestamp 1644511149
transform 1 0 32200 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_350
timestamp 1644511149
transform 1 0 33304 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1644511149
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_173
timestamp 1644511149
transform 1 0 17020 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_177
timestamp 1644511149
transform 1 0 17388 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_187
timestamp 1644511149
transform 1 0 18308 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1644511149
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_233
timestamp 1644511149
transform 1 0 22540 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_243
timestamp 1644511149
transform 1 0 23460 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_251
timestamp 1644511149
transform 1 0 24196 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_255
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_260
timestamp 1644511149
transform 1 0 25024 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_268
timestamp 1644511149
transform 1 0 25760 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_272
timestamp 1644511149
transform 1 0 26128 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1644511149
transform 1 0 27416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_307
timestamp 1644511149
transform 1 0 29348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_319
timestamp 1644511149
transform 1 0 30452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_331
timestamp 1644511149
transform 1 0 31556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_154
timestamp 1644511149
transform 1 0 15272 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_164
timestamp 1644511149
transform 1 0 16192 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_176
timestamp 1644511149
transform 1 0 17296 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_188
timestamp 1644511149
transform 1 0 18400 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_214
timestamp 1644511149
transform 1 0 20792 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_226
timestamp 1644511149
transform 1 0 21896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_232
timestamp 1644511149
transform 1 0 22448 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_244
timestamp 1644511149
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_272
timestamp 1644511149
transform 1 0 26128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_278
timestamp 1644511149
transform 1 0 26680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_285
timestamp 1644511149
transform 1 0 27324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_296
timestamp 1644511149
transform 1 0 28336 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_159
timestamp 1644511149
transform 1 0 15732 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_172
timestamp 1644511149
transform 1 0 16928 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_178
timestamp 1644511149
transform 1 0 17480 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_186
timestamp 1644511149
transform 1 0 18216 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_198
timestamp 1644511149
transform 1 0 19320 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_210
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_233
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_240
timestamp 1644511149
transform 1 0 23184 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_251
timestamp 1644511149
transform 1 0 24196 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_263
timestamp 1644511149
transform 1 0 25300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1644511149
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_290
timestamp 1644511149
transform 1 0 27784 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_296
timestamp 1644511149
transform 1 0 28336 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_508
timestamp 1644511149
transform 1 0 47840 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_163
timestamp 1644511149
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1644511149
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1644511149
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_200
timestamp 1644511149
transform 1 0 19504 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_212
timestamp 1644511149
transform 1 0 20608 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_217
timestamp 1644511149
transform 1 0 21068 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_229
timestamp 1644511149
transform 1 0 22172 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_235
timestamp 1644511149
transform 1 0 22724 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1644511149
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_260
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_272
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_290
timestamp 1644511149
transform 1 0 27784 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_298
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_465
timestamp 1644511149
transform 1 0 43884 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_471
timestamp 1644511149
transform 1 0 44436 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_486
timestamp 1644511149
transform 1 0 45816 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_490
timestamp 1644511149
transform 1 0 46184 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_192
timestamp 1644511149
transform 1 0 18768 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_200
timestamp 1644511149
transform 1 0 19504 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_206
timestamp 1644511149
transform 1 0 20056 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_210
timestamp 1644511149
transform 1 0 20424 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_214
timestamp 1644511149
transform 1 0 20792 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1644511149
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_233
timestamp 1644511149
transform 1 0 22540 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_242
timestamp 1644511149
transform 1 0 23368 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_260
timestamp 1644511149
transform 1 0 25024 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_264
timestamp 1644511149
transform 1 0 25392 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_268
timestamp 1644511149
transform 1 0 25760 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_288
timestamp 1644511149
transform 1 0 27600 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_300
timestamp 1644511149
transform 1 0 28704 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_312
timestamp 1644511149
transform 1 0 29808 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_324
timestamp 1644511149
transform 1 0 30912 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_479
timestamp 1644511149
transform 1 0 45172 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_491
timestamp 1644511149
transform 1 0 46276 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_168
timestamp 1644511149
transform 1 0 16560 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_180
timestamp 1644511149
transform 1 0 17664 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_192
timestamp 1644511149
transform 1 0 18768 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_220
timestamp 1644511149
transform 1 0 21344 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_246
timestamp 1644511149
transform 1 0 23736 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_273
timestamp 1644511149
transform 1 0 26220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_297
timestamp 1644511149
transform 1 0 28428 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_305
timestamp 1644511149
transform 1 0 29164 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_472
timestamp 1644511149
transform 1 0 44528 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_493
timestamp 1644511149
transform 1 0 46460 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_500
timestamp 1644511149
transform 1 0 47104 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_210
timestamp 1644511149
transform 1 0 20424 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1644511149
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_229
timestamp 1644511149
transform 1 0 22172 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_240
timestamp 1644511149
transform 1 0 23184 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_247
timestamp 1644511149
transform 1 0 23828 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_259
timestamp 1644511149
transform 1 0 24932 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_271
timestamp 1644511149
transform 1 0 26036 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_289
timestamp 1644511149
transform 1 0 27692 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_498
timestamp 1644511149
transform 1 0 46920 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_203
timestamp 1644511149
transform 1 0 19780 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_208
timestamp 1644511149
transform 1 0 20240 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_240
timestamp 1644511149
transform 1 0 23184 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_480
timestamp 1644511149
transform 1 0 45264 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_488
timestamp 1644511149
transform 1 0 46000 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_214
timestamp 1644511149
transform 1 0 20792 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1644511149
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_231
timestamp 1644511149
transform 1 0 22356 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_235
timestamp 1644511149
transform 1 0 22724 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_246
timestamp 1644511149
transform 1 0 23736 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_250
timestamp 1644511149
transform 1 0 24104 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_262
timestamp 1644511149
transform 1 0 25208 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_274
timestamp 1644511149
transform 1 0 26312 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_227
timestamp 1644511149
transform 1 0 21988 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_231
timestamp 1644511149
transform 1 0 22356 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_243
timestamp 1644511149
transform 1 0 23460 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_284
timestamp 1644511149
transform 1 0 27232 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_296
timestamp 1644511149
transform 1 0 28336 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_308
timestamp 1644511149
transform 1 0 29440 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_320
timestamp 1644511149
transform 1 0 30544 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_332
timestamp 1644511149
transform 1 0 31648 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_14
timestamp 1644511149
transform 1 0 2392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1644511149
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_281
timestamp 1644511149
transform 1 0 26956 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_303
timestamp 1644511149
transform 1 0 28980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_451
timestamp 1644511149
transform 1 0 42596 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_455
timestamp 1644511149
transform 1 0 42964 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_462
timestamp 1644511149
transform 1 0 43608 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_468
timestamp 1644511149
transform 1 0 44160 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_28
timestamp 1644511149
transform 1 0 3680 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_40
timestamp 1644511149
transform 1 0 4784 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1644511149
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_117
timestamp 1644511149
transform 1 0 11868 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_121
timestamp 1644511149
transform 1 0 12236 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_133
timestamp 1644511149
transform 1 0 13340 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_145
timestamp 1644511149
transform 1 0 14444 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_157
timestamp 1644511149
transform 1 0 15548 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1644511149
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_219
timestamp 1644511149
transform 1 0 21252 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_286
timestamp 1644511149
transform 1 0 27416 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_298
timestamp 1644511149
transform 1 0 28520 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_310
timestamp 1644511149
transform 1 0 29624 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_322
timestamp 1644511149
transform 1 0 30728 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1644511149
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_437
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_472
timestamp 1644511149
transform 1 0 44528 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1644511149
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_509
timestamp 1644511149
transform 1 0 47932 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_515
timestamp 1644511149
transform 1 0 48484 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_7
timestamp 1644511149
transform 1 0 1748 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1644511149
transform 1 0 2116 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1644511149
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_36
timestamp 1644511149
transform 1 0 4416 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_45
timestamp 1644511149
transform 1 0 5244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_57
timestamp 1644511149
transform 1 0 6348 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_69
timestamp 1644511149
transform 1 0 7452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_81
timestamp 1644511149
transform 1 0 8556 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_125
timestamp 1644511149
transform 1 0 12604 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_208
timestamp 1644511149
transform 1 0 20240 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_235
timestamp 1644511149
transform 1 0 22724 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1644511149
transform 1 0 23828 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_336
timestamp 1644511149
transform 1 0 32016 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_348
timestamp 1644511149
transform 1 0 33120 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1644511149
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_458
timestamp 1644511149
transform 1 0 43240 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_465
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1644511149
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_7
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_19
timestamp 1644511149
transform 1 0 2852 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_358
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_370
timestamp 1644511149
transform 1 0 35144 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_382
timestamp 1644511149
transform 1 0 36248 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_390
timestamp 1644511149
transform 1 0 36984 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1644511149
transform 1 0 6900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_151
timestamp 1644511149
transform 1 0 14996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_163
timestamp 1644511149
transform 1 0 16100 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_207
timestamp 1644511149
transform 1 0 20148 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_82_218
timestamp 1644511149
transform 1 0 21160 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_228
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_235
timestamp 1644511149
transform 1 0 22724 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_247
timestamp 1644511149
transform 1 0 23828 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1644511149
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_258
timestamp 1644511149
transform 1 0 24840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_262
timestamp 1644511149
transform 1 0 25208 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_266
timestamp 1644511149
transform 1 0 25576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1644511149
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_323
timestamp 1644511149
transform 1 0 30820 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_328
timestamp 1644511149
transform 1 0 31280 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1644511149
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_453
timestamp 1644511149
transform 1 0 42780 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1644511149
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0597_
timestamp 1644511149
transform 1 0 32568 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0601_
timestamp 1644511149
transform 1 0 30176 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29348 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0603_
timestamp 1644511149
transform 1 0 18400 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0604_
timestamp 1644511149
transform 1 0 16192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0605_
timestamp 1644511149
transform 1 0 17848 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0606_
timestamp 1644511149
transform 1 0 26772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0607_
timestamp 1644511149
transform 1 0 22816 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0608_
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0609_
timestamp 1644511149
transform 1 0 21068 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0611_
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0612_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0615_
timestamp 1644511149
transform 1 0 24932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32568 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0618_
timestamp 1644511149
transform 1 0 21160 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14904 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0620_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0621_
timestamp 1644511149
transform 1 0 18952 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0622_
timestamp 1644511149
transform 1 0 23920 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0623_
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0624_
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0625_
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0626_
timestamp 1644511149
transform 1 0 19320 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0627_
timestamp 1644511149
transform 1 0 20148 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0628_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33028 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0630_
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33580 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1644511149
transform 1 0 32476 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0633_
timestamp 1644511149
transform 1 0 34040 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0634_
timestamp 1644511149
transform 1 0 32108 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1644511149
transform 1 0 35512 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0639_
timestamp 1644511149
transform 1 0 33856 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1644511149
transform 1 0 35144 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0641_
timestamp 1644511149
transform 1 0 32200 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0642_
timestamp 1644511149
transform 1 0 33580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0643_
timestamp 1644511149
transform 1 0 33856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0644_
timestamp 1644511149
transform 1 0 30084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0646_
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0648_
timestamp 1644511149
transform 1 0 31280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1644511149
transform 1 0 29624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0651_
timestamp 1644511149
transform 1 0 28336 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1644511149
transform 1 0 22724 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 1644511149
transform 1 0 19320 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0656_
timestamp 1644511149
transform 1 0 13248 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0657_
timestamp 1644511149
transform 1 0 20608 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1644511149
transform 1 0 22724 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0660_
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19320 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 17572 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0665_
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14904 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0670_
timestamp 1644511149
transform 1 0 12880 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14720 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1644511149
transform 1 0 13156 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0674_
timestamp 1644511149
transform 1 0 12420 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 1644511149
transform 1 0 12512 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0677_
timestamp 1644511149
transform 1 0 12052 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1644511149
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0680_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0682_
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0683_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0684_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1644511149
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1644511149
transform 1 0 13616 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0687_
timestamp 1644511149
transform 1 0 16100 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0688_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0690_
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0692_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14536 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0694_
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0695_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1644511149
transform 1 0 19504 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1644511149
transform 1 0 21528 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0698_
timestamp 1644511149
transform 1 0 20240 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0701_
timestamp 1644511149
transform 1 0 20332 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0702_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0704_
timestamp 1644511149
transform 1 0 19504 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0705_
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1644511149
transform 1 0 21712 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0707_
timestamp 1644511149
transform 1 0 20516 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1644511149
transform 1 0 21712 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0709_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0710_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0711_
timestamp 1644511149
transform 1 0 23092 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0712_
timestamp 1644511149
transform 1 0 22908 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0713_
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0714_
timestamp 1644511149
transform 1 0 26128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0716_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0717_
timestamp 1644511149
transform 1 0 25024 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0719_
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0721_
timestamp 1644511149
transform 1 0 24656 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0722_
timestamp 1644511149
transform 1 0 23552 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 1644511149
transform 1 0 23460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_
timestamp 1644511149
transform 1 0 24840 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0728_
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1644511149
transform 1 0 25392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1644511149
transform 1 0 27324 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 27784 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 1644511149
transform 1 0 24840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0733_
timestamp 1644511149
transform 1 0 25576 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1644511149
transform 1 0 28428 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0735_
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1644511149
transform 1 0 26312 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0738_
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0739_
timestamp 1644511149
transform 1 0 28520 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0740_
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0743_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0744_
timestamp 1644511149
transform 1 0 24196 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1644511149
transform 1 0 25668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0746_
timestamp 1644511149
transform 1 0 24840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0748_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0749_
timestamp 1644511149
transform 1 0 24840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0750_
timestamp 1644511149
transform 1 0 20976 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0751_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0752_
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0755_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0756_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0757_
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0758_
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0759_
timestamp 1644511149
transform 1 0 19228 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0761_
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0762_
timestamp 1644511149
transform 1 0 19412 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0763_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19320 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _0764_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0765_
timestamp 1644511149
transform 1 0 25760 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0766_
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0767_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1644511149
transform 1 0 17020 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1644511149
transform 1 0 17112 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0771_
timestamp 1644511149
transform 1 0 24196 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1644511149
transform 1 0 20700 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0773_
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0774_
timestamp 1644511149
transform 1 0 21068 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0775_
timestamp 1644511149
transform 1 0 22080 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0776_
timestamp 1644511149
transform 1 0 27784 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0777_
timestamp 1644511149
transform 1 0 24564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0778_
timestamp 1644511149
transform 1 0 20424 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0779_
timestamp 1644511149
transform 1 0 20332 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0780_
timestamp 1644511149
transform 1 0 20516 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1644511149
transform 1 0 19320 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0783_
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0784_
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0786_
timestamp 1644511149
transform 1 0 22172 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0787_
timestamp 1644511149
transform 1 0 21988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0788_
timestamp 1644511149
transform 1 0 20332 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0789_
timestamp 1644511149
transform 1 0 19872 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0790_
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _0791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0792_
timestamp 1644511149
transform 1 0 22540 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1644511149
transform 1 0 22080 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0795_
timestamp 1644511149
transform 1 0 24656 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1644511149
transform 1 0 27140 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0797_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0798_
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0799_
timestamp 1644511149
transform 1 0 19596 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1644511149
transform 1 0 23736 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0801_
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0803_
timestamp 1644511149
transform 1 0 23736 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0805_
timestamp 1644511149
transform 1 0 24472 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0806_
timestamp 1644511149
transform 1 0 24748 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0807_
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0808_
timestamp 1644511149
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0809_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0810_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0811_
timestamp 1644511149
transform 1 0 22632 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0812_
timestamp 1644511149
transform 1 0 20424 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0813_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0814_
timestamp 1644511149
transform 1 0 27324 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0815_
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0816_
timestamp 1644511149
transform 1 0 28520 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1644511149
transform 1 0 26496 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0818_
timestamp 1644511149
transform 1 0 27048 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0819_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0820_
timestamp 1644511149
transform 1 0 26680 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1644511149
transform 1 0 27416 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0822_
timestamp 1644511149
transform 1 0 25852 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0823_
timestamp 1644511149
transform 1 0 25760 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0824_
timestamp 1644511149
transform 1 0 25576 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0825_
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0826_
timestamp 1644511149
transform 1 0 25668 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0827_
timestamp 1644511149
transform 1 0 15548 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0829_
timestamp 1644511149
transform 1 0 29624 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1644511149
transform 1 0 15272 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0832_
timestamp 1644511149
transform 1 0 17020 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0833_
timestamp 1644511149
transform 1 0 23092 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0834_
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1644511149
transform 1 0 23644 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1644511149
transform 1 0 23000 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0837_
timestamp 1644511149
transform 1 0 16836 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0838_
timestamp 1644511149
transform 1 0 16928 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0839_
timestamp 1644511149
transform 1 0 16008 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0840_
timestamp 1644511149
transform 1 0 14444 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0841_
timestamp 1644511149
transform 1 0 15640 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0842_
timestamp 1644511149
transform 1 0 16836 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0843_
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1644511149
transform 1 0 14628 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0845_
timestamp 1644511149
transform 1 0 15456 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1644511149
transform 1 0 15640 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0847_
timestamp 1644511149
transform 1 0 13616 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0848_
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0849_
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0850_
timestamp 1644511149
transform 1 0 14352 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0851_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0852_
timestamp 1644511149
transform 1 0 14536 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0853_
timestamp 1644511149
transform 1 0 14444 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0854_
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0855_
timestamp 1644511149
transform 1 0 17296 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0856_
timestamp 1644511149
transform 1 0 17204 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0857_
timestamp 1644511149
transform 1 0 17572 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0858_
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0859_
timestamp 1644511149
transform 1 0 17204 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0861_
timestamp 1644511149
transform 1 0 29992 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30544 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0864_
timestamp 1644511149
transform 1 0 31464 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1644511149
transform 1 0 28520 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0866_
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0867_
timestamp 1644511149
transform 1 0 26772 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0868_
timestamp 1644511149
transform 1 0 29624 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0869_
timestamp 1644511149
transform 1 0 30360 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0870_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform 1 0 29440 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0872_
timestamp 1644511149
transform 1 0 29716 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1644511149
transform 1 0 29808 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0874_
timestamp 1644511149
transform 1 0 30728 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0875_
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0876_
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0877_
timestamp 1644511149
transform 1 0 29992 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0878_
timestamp 1644511149
transform 1 0 31464 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0879_
timestamp 1644511149
transform 1 0 29992 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0880_
timestamp 1644511149
transform 1 0 29256 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0881_
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1644511149
transform 1 0 28336 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0883_
timestamp 1644511149
transform 1 0 27876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1644511149
transform 1 0 28336 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0887_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1644511149
transform 1 0 25576 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0889_
timestamp 1644511149
transform 1 0 29624 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0890_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 20976 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 27140 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 43056 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0902_
timestamp 1644511149
transform 1 0 30360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 44068 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 29072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1644511149
transform 1 0 27508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0915_
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 41400 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0921_
timestamp 1644511149
transform 1 0 25116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 37536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 39376 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 46644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 23184 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 41492 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 30452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17940 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 14996 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 15640 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 15088 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0939_
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 17112 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1644511149
transform 1 0 44068 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  _0946_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43516 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 42780 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 31188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 22356 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0958_
timestamp 1644511149
transform 1 0 44068 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 11960 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 42964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 44896 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 38732 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0964_
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 47288 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 4968 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0970_
timestamp 1644511149
transform 1 0 43608 0 -1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 43608 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 23276 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0976_
timestamp 1644511149
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0977_
timestamp 1644511149
transform 1 0 22172 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 11776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0983_
timestamp 1644511149
transform 1 0 28336 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 28520 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 32384 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 46828 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0989_
timestamp 1644511149
transform 1 0 30636 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 33028 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 47932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 42688 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0995_
timestamp 1644511149
transform 1 0 20240 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 19964 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1001_
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 29716 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform 1 0 33028 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41124 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45816 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1015_
timestamp 1644511149
transform 1 0 46092 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1016_
timestamp 1644511149
transform 1 0 46552 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1644511149
transform 1 0 45632 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1644511149
transform 1 0 45908 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1644511149
transform 1 0 43700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1021_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1644511149
transform 1 0 44528 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1023_
timestamp 1644511149
transform 1 0 47472 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1024_
timestamp 1644511149
transform 1 0 40204 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1026_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40204 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1644511149
transform 1 0 39560 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1029_
timestamp 1644511149
transform 1 0 40388 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1644511149
transform 1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _1032_
timestamp 1644511149
transform 1 0 42780 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1644511149
transform 1 0 43608 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1644511149
transform 1 0 42964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1035_
timestamp 1644511149
transform 1 0 42320 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1036_
timestamp 1644511149
transform 1 0 43792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1644511149
transform 1 0 46736 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1644511149
transform 1 0 27048 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 1644511149
transform 1 0 27784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1040_
timestamp 1644511149
transform 1 0 27600 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 1644511149
transform 1 0 27048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1042_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1043_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1044_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1045_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1644511149
transform 1 0 43056 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1047_
timestamp 1644511149
transform 1 0 43056 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43056 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1049_
timestamp 1644511149
transform 1 0 43332 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1644511149
transform 1 0 42780 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42964 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1644511149
transform 1 0 44160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44344 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1056_
timestamp 1644511149
transform 1 0 45172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1057_
timestamp 1644511149
transform 1 0 43608 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1058_
timestamp 1644511149
transform 1 0 28520 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1061_
timestamp 1644511149
transform 1 0 28704 0 -1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1644511149
transform 1 0 27048 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1064_
timestamp 1644511149
transform 1 0 28336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1065_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 1644511149
transform 1 0 29256 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 1644511149
transform 1 0 43240 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1644511149
transform 1 0 42504 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1071_
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1072_
timestamp 1644511149
transform 1 0 41124 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1073_
timestamp 1644511149
transform 1 0 32936 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1075_
timestamp 1644511149
transform 1 0 25668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1644511149
transform 1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1077_
timestamp 1644511149
transform 1 0 1840 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1079_
timestamp 1644511149
transform 1 0 46276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1081_
timestamp 1644511149
transform 1 0 34776 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform 1 0 34408 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1083_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1085_
timestamp 1644511149
transform 1 0 40204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1644511149
transform 1 0 40664 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1087_
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1089_
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 27232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 29716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1093_
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 32752 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1099_
timestamp 1644511149
transform 1 0 17848 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1644511149
transform 1 0 17112 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1644511149
transform 1 0 15548 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1644511149
transform 1 0 14168 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1644511149
transform 1 0 18308 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1644511149
transform 1 0 17664 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1111_
timestamp 1644511149
transform 1 0 20056 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1644511149
transform 1 0 27784 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 23552 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 20516 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1117_
timestamp 1644511149
transform 1 0 19872 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1644511149
transform 1 0 21896 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1644511149
transform 1 0 20516 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1644511149
transform 1 0 20056 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1123_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1644511149
transform 1 0 22448 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1644511149
transform 1 0 25208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1128_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1129_
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1130_
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1644511149
transform 1 0 26036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1132_
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1133_
timestamp 1644511149
transform 1 0 22724 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1134_
timestamp 1644511149
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1135_
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1136_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1137_
timestamp 1644511149
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1138_
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1644511149
transform 1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1140_
timestamp 1644511149
transform 1 0 17296 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1141_
timestamp 1644511149
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1644511149
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1143_
timestamp 1644511149
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1144_
timestamp 1644511149
transform 1 0 12972 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1145_
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1146_
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1147_
timestamp 1644511149
transform 1 0 11776 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1644511149
transform 1 0 11868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1149_
timestamp 1644511149
transform 1 0 11684 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1150_
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1644511149
transform 1 0 15088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1152_
timestamp 1644511149
transform 1 0 15732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1153_
timestamp 1644511149
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1154_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1155_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1156_
timestamp 1644511149
transform 1 0 27876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1157_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1158_
timestamp 1644511149
transform 1 0 30544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1159_
timestamp 1644511149
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1160_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1162_
timestamp 1644511149
transform 1 0 33304 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1163_
timestamp 1644511149
transform 1 0 31280 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1644511149
transform 1 0 32936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1644511149
transform 1 0 24472 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1644511149
transform 1 0 27968 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1644511149
transform 1 0 30820 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1644511149
transform 1 0 16744 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1644511149
transform 1 0 13800 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1644511149
transform 1 0 13892 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1644511149
transform 1 0 17480 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1644511149
transform 1 0 22172 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1644511149
transform 1 0 21896 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 1644511149
transform 1 0 19504 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1644511149
transform 1 0 21344 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1644511149
transform 1 0 19504 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1644511149
transform 1 0 19964 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1644511149
transform 1 0 21988 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1644511149
transform 1 0 17020 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1644511149
transform 1 0 18952 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1644511149
transform 1 0 21620 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1200_
timestamp 1644511149
transform 1 0 25392 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1644511149
transform 1 0 25392 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1203_
timestamp 1644511149
transform 1 0 25300 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1206_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1644511149
transform 1 0 17664 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1644511149
transform 1 0 16928 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1210_
timestamp 1644511149
transform 1 0 13340 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1644511149
transform 1 0 11500 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1214_
timestamp 1644511149
transform 1 0 11500 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1215_
timestamp 1644511149
transform 1 0 12420 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 1644511149
transform 1 0 11684 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 1644511149
transform 1 0 14628 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 1644511149
transform 1 0 21252 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1222_
timestamp 1644511149
transform 1 0 28704 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1223_
timestamp 1644511149
transform 1 0 31004 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 1644511149
transform 1 0 31280 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1226_
timestamp 1644511149
transform 1 0 34868 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1644511149
transform 1 0 33856 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1230_
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__conb_1  _1231__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1232__82
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1233__83
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1234__84
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1235__85
timestamp 1644511149
transform 1 0 47472 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1236__86
timestamp 1644511149
transform 1 0 20884 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1237__87
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1238__88
timestamp 1644511149
transform 1 0 24564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1239__89
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1240__90
timestamp 1644511149
transform 1 0 25300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1241__91
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1242__92
timestamp 1644511149
transform 1 0 1840 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1243__93
timestamp 1644511149
transform 1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1244__94
timestamp 1644511149
transform 1 0 4140 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1245__95
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1246__96
timestamp 1644511149
transform 1 0 43608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1247__97
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1248__98
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1249__99
timestamp 1644511149
transform 1 0 45632 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1250__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1251__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1252__102
timestamp 1644511149
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1253__103
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1254__104
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1255__105
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1256__106
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1257__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1258__108
timestamp 1644511149
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1259__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1260__110
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1261__111
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1262__112
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1263__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1264__114
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1265__115
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1266__116
timestamp 1644511149
transform 1 0 43332 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1267__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1268__118
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1269__119
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1270__120
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1271__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1272__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1273__123
timestamp 1644511149
transform 1 0 46368 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1274__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1275__125
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1276__126
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1277__127
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1278__128
timestamp 1644511149
transform 1 0 47748 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1279__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1280__130
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1281__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1282__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1283__133
timestamp 1644511149
transform 1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1284__134
timestamp 1644511149
transform 1 0 47472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1285__135
timestamp 1644511149
transform 1 0 42504 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 29716 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 43884 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 44068 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 45448 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 42596 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 44988 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 38824 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 27048 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 46276 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 20792 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 32200 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 42596 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1315_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1316_
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1317_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1318_
timestamp 1644511149
transform 1 0 29716 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1319_
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1320_
timestamp 1644511149
transform 1 0 21988 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1321_
timestamp 1644511149
transform 1 0 23368 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1322_
timestamp 1644511149
transform 1 0 15640 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1323_
timestamp 1644511149
transform 1 0 30360 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1324_
timestamp 1644511149
transform 1 0 22724 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1325_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1326_
timestamp 1644511149
transform 1 0 42596 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1327_
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1328_
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1329_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1330_
timestamp 1644511149
transform 1 0 11684 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1331_
timestamp 1644511149
transform 1 0 17204 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1332_
timestamp 1644511149
transform 1 0 14260 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1333_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1334_
timestamp 1644511149
transform 1 0 14260 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1335_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1336_
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1337_
timestamp 1644511149
transform 1 0 15824 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1338_
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1339_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1340_
timestamp 1644511149
transform 1 0 23828 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1341_
timestamp 1644511149
transform 1 0 14904 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1342_
timestamp 1644511149
transform 1 0 28244 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1343_
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1344_
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1345_
timestamp 1644511149
transform 1 0 36984 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1346_
timestamp 1644511149
transform 1 0 37444 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 42136 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 32292 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 32936 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 22816 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 1840 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 24472 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 42596 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 46276 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1372_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1373_
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1374_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1375_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1376_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1377_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1378_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1379_
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1380_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1381_
timestamp 1644511149
transform 1 0 44896 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 20976 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 19688 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 22632 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 27416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 47288 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 47932 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 47932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1644511149
transform 1 0 47840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 12328 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 22448 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 46460 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 47656 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1644511149
transform 1 0 31004 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 43148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 11684 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46184 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 45448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 40020 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39376 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 40572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 15824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 19872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33028 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2024 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35052 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 40664 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 36800 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2852 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45448 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35420 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46736 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 41768 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37444 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 41400 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 45172 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 40480 0 1 22848
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
